module fake_ariane_3192_n_16275 (n_2752, n_3527, n_913, n_1681, n_2163, n_3432, n_4030, n_1486, n_1507, n_1938, n_3619, n_589, n_2484, n_2866, n_3153, n_1174, n_4013, n_3152, n_2346, n_3434, n_1469, n_691, n_1353, n_3056, n_3500, n_3480, n_2679, n_1355, n_2131, n_3268, n_3853, n_2559, n_2500, n_2509, n_423, n_4085, n_1383, n_2182, n_603, n_373, n_2135, n_2334, n_2680, n_3264, n_1250, n_2030, n_1169, n_789, n_3181, n_850, n_2993, n_1916, n_2879, n_610, n_245, n_1713, n_96, n_319, n_49, n_1436, n_2407, n_690, n_2818, n_416, n_3578, n_1109, n_1430, n_2537, n_525, n_187, n_3745, n_2002, n_1463, n_2243, n_3487, n_1238, n_2694, n_3668, n_2011, n_3742, n_2729, n_1515, n_817, n_1837, n_924, n_781, n_2013, n_2786, n_1566, n_2837, n_189, n_717, n_3765, n_72, n_2006, n_4058, n_952, n_864, n_4090, n_2446, n_1096, n_4116, n_1379, n_2436, n_57, n_3352, n_3517, n_2376, n_2367, n_2671, n_2790, n_1706, n_2207, n_2461, n_2702, n_3719, n_117, n_524, n_2731, n_3703, n_1214, n_634, n_3561, n_1839, n_1246, n_1138, n_214, n_3526, n_3888, n_3954, n_2042, n_2123, n_3198, n_1853, n_764, n_1503, n_2238, n_2529, n_2374, n_4103, n_462, n_1196, n_1181, n_32, n_1999, n_3435, n_410, n_2380, n_1187, n_1131, n_1225, n_3154, n_2646, n_737, n_137, n_1298, n_2653, n_1745, n_2873, n_1366, n_232, n_52, n_2084, n_3115, n_3938, n_568, n_2278, n_4028, n_3330, n_3514, n_1088, n_77, n_1424, n_766, n_2976, n_1835, n_3383, n_3965, n_1457, n_377, n_2482, n_3905, n_1682, n_2750, n_3797, n_1836, n_3416, n_520, n_870, n_2547, n_3382, n_1453, n_279, n_945, n_958, n_3943, n_3930, n_2554, n_3145, n_3808, n_2248, n_3665, n_3063, n_813, n_3281, n_3535, n_419, n_1985, n_2288, n_2621, n_2908, n_3081, n_146, n_3858, n_270, n_4106, n_338, n_995, n_2579, n_285, n_1909, n_2156, n_1184, n_1961, n_202, n_1535, n_3220, n_2960, n_500, n_665, n_754, n_903, n_3270, n_871, n_2323, n_1073, n_2844, n_3348, n_239, n_402, n_1979, n_1277, n_2107, n_1746, n_3261, n_54, n_829, n_1761, n_1062, n_339, n_738, n_3679, n_1690, n_2221, n_2807, n_672, n_740, n_1283, n_167, n_2317, n_2838, n_1974, n_2906, n_1736, n_1018, n_2342, n_2200, n_2781, n_3283, n_3856, n_4038, n_69, n_259, n_2442, n_2735, n_953, n_1364, n_2390, n_143, n_1888, n_1224, n_3657, n_2109, n_1425, n_2634, n_2709, n_3451, n_625, n_557, n_2322, n_2746, n_3419, n_1107, n_2832, n_1688, n_989, n_242, n_645, n_1944, n_331, n_559, n_2233, n_2370, n_2663, n_267, n_495, n_2914, n_1988, n_350, n_381, n_795, n_721, n_1084, n_3545, n_1718, n_1276, n_1936, n_2149, n_2277, n_200, n_1428, n_1284, n_2878, n_1241, n_3890, n_3830, n_821, n_561, n_770, n_3252, n_1514, n_2539, n_1528, n_507, n_486, n_901, n_2782, n_3879, n_569, n_2078, n_3315, n_3929, n_1145, n_3523, n_971, n_3144, n_2359, n_3999, n_2201, n_787, n_4012, n_1650, n_31, n_1519, n_1195, n_2049, n_1522, n_518, n_1207, n_222, n_3606, n_786, n_1404, n_3347, n_3420, n_3859, n_868, n_3474, n_2232, n_1847, n_2458, n_2779, n_3627, n_3596, n_3150, n_2950, n_1542, n_3552, n_1314, n_3756, n_3639, n_3254, n_1512, n_2227, n_2301, n_1539, n_2859, n_3121, n_2847, n_884, n_3412, n_4077, n_1851, n_2162, n_3209, n_3324, n_3015, n_1415, n_3870, n_1034, n_1652, n_2192, n_1676, n_3749, n_1085, n_277, n_2988, n_1636, n_3482, n_432, n_293, n_823, n_1900, n_620, n_3948, n_93, n_1074, n_3230, n_859, n_3793, n_1765, n_4031, n_108, n_1889, n_587, n_1977, n_693, n_863, n_2650, n_303, n_1254, n_3960, n_929, n_3207, n_3641, n_2433, n_206, n_352, n_899, n_1703, n_2332, n_2391, n_3828, n_3975, n_3073, n_611, n_1295, n_2060, n_1850, n_238, n_365, n_2004, n_3183, n_3571, n_1013, n_3883, n_4032, n_4018, n_1495, n_3607, n_1637, n_3297, n_2571, n_136, n_334, n_2427, n_192, n_3325, n_3613, n_2885, n_661, n_2098, n_2616, n_1751, n_2874, n_3003, n_4117, n_300, n_533, n_3049, n_3136, n_2867, n_3634, n_1917, n_2456, n_2769, n_104, n_1924, n_438, n_1560, n_1654, n_2341, n_2899, n_1548, n_3066, n_16, n_1811, n_2045, n_3274, n_3877, n_440, n_3913, n_3817, n_3013, n_3612, n_273, n_2575, n_2722, n_1396, n_3728, n_1230, n_612, n_333, n_1840, n_2739, n_3739, n_376, n_3962, n_512, n_1597, n_4082, n_2942, n_1771, n_2902, n_1544, n_579, n_3271, n_844, n_1012, n_1267, n_2061, n_2685, n_3164, n_2094, n_3854, n_3861, n_2512, n_1354, n_1790, n_149, n_1213, n_2382, n_2956, n_237, n_2043, n_780, n_2349, n_1918, n_3652, n_3449, n_2788, n_4119, n_1021, n_1443, n_4000, n_3089, n_491, n_2595, n_1465, n_2686, n_3084, n_1949, n_1595, n_1142, n_1140, n_705, n_3458, n_570, n_260, n_2727, n_942, n_3580, n_1437, n_3860, n_3511, n_7, n_2077, n_1378, n_461, n_1121, n_1416, n_2909, n_209, n_490, n_3554, n_1461, n_17, n_2717, n_3012, n_1391, n_2981, n_1947, n_225, n_1599, n_1876, n_1006, n_1830, n_3850, n_575, n_546, n_3472, n_503, n_2527, n_1112, n_700, n_1159, n_772, n_1216, n_3126, n_3754, n_2759, n_1245, n_2743, n_1669, n_2969, n_3429, n_1675, n_2466, n_676, n_3758, n_42, n_2038, n_2263, n_3518, n_3958, n_2800, n_2568, n_2116, n_2271, n_2145, n_2326, n_1838, n_3485, n_1594, n_680, n_1935, n_2806, n_287, n_3191, n_1716, n_4108, n_302, n_3777, n_4109, n_1872, n_380, n_3562, n_1585, n_2281, n_1432, n_94, n_2245, n_4, n_3359, n_3767, n_3841, n_3119, n_249, n_1108, n_3588, n_355, n_212, n_65, n_123, n_444, n_851, n_1590, n_1351, n_3234, n_3280, n_3413, n_3692, n_3900, n_2216, n_4115, n_1274, n_3539, n_257, n_2426, n_652, n_1819, n_475, n_135, n_3095, n_947, n_2134, n_3862, n_930, n_1260, n_3698, n_3716, n_1179, n_468, n_3284, n_3909, n_102, n_2703, n_182, n_696, n_1442, n_2926, n_482, n_2620, n_798, n_577, n_1833, n_407, n_1691, n_27, n_916, n_1386, n_2810, n_3391, n_3506, n_912, n_1884, n_460, n_1555, n_1842, n_2499, n_2549, n_3678, n_366, n_762, n_1253, n_1468, n_1661, n_2791, n_555, n_2683, n_3212, n_804, n_1656, n_1382, n_3093, n_3529, n_2970, n_3159, n_966, n_992, n_955, n_3549, n_3885, n_3914, n_3624, n_1182, n_794, n_2855, n_78, n_2166, n_2848, n_1692, n_3192, n_2611, n_1562, n_514, n_2748, n_418, n_2185, n_3306, n_3250, n_3029, n_2398, n_3538, n_3915, n_1376, n_3839, n_513, n_288, n_179, n_1292, n_1178, n_1972, n_2015, n_2925, n_1435, n_3407, n_3717, n_1750, n_1026, n_1506, n_3460, n_3544, n_1610, n_3875, n_4029, n_2202, n_2072, n_3852, n_306, n_2952, n_3530, n_2415, n_2693, n_2877, n_92, n_4099, n_3120, n_203, n_2922, n_436, n_3000, n_150, n_2871, n_2930, n_3193, n_3240, n_324, n_2745, n_2087, n_669, n_931, n_1491, n_2628, n_3219, n_3362, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_3937, n_2161, n_1418, n_746, n_1357, n_292, n_1079, n_1787, n_2462, n_3510, n_1389, n_3393, n_3172, n_2155, n_2659, n_4033, n_615, n_3747, n_1139, n_2836, n_3688, n_76, n_2439, n_2864, n_517, n_1312, n_1717, n_3604, n_4045, n_0, n_1812, n_3651, n_824, n_428, n_159, n_2172, n_2601, n_3614, n_3871, n_892, n_1880, n_959, n_30, n_2365, n_2257, n_3757, n_1399, n_1101, n_1567, n_1343, n_563, n_2219, n_3116, n_1855, n_3784, n_2100, n_2333, n_3176, n_144, n_3629, n_3666, n_3372, n_3891, n_990, n_1623, n_3559, n_1903, n_3792, n_867, n_2147, n_3479, n_4020, n_2435, n_1226, n_2224, n_944, n_749, n_1932, n_1780, n_2825, n_2888, n_1970, n_3998, n_3724, n_1920, n_2083, n_815, n_542, n_3287, n_2167, n_2293, n_2753, n_1340, n_470, n_2668, n_1240, n_2921, n_3046, n_1087, n_4055, n_3980, n_2701, n_2400, n_3021, n_632, n_3257, n_477, n_650, n_3741, n_2388, n_425, n_3730, n_2273, n_2712, n_1433, n_3805, n_1911, n_3979, n_3912, n_2567, n_3950, n_3496, n_3493, n_2557, n_2695, n_2898, n_1825, n_1908, n_1155, n_2598, n_1071, n_2755, n_3700, n_3727, n_712, n_976, n_3567, n_909, n_4003, n_1392, n_767, n_1832, n_2795, n_2682, n_1841, n_1680, n_2066, n_2302, n_2762, n_964, n_1627, n_2220, n_2954, n_382, n_3014, n_489, n_2294, n_80, n_2274, n_3342, n_2895, n_2903, n_251, n_974, n_506, n_3814, n_3812, n_3127, n_3796, n_1731, n_799, n_3884, n_1147, n_2829, n_2378, n_3625, n_397, n_2467, n_3375, n_2768, n_471, n_351, n_965, n_1914, n_155, n_3760, n_2253, n_934, n_2213, n_3515, n_1447, n_2363, n_1220, n_356, n_2019, n_698, n_4056, n_2728, n_2130, n_1674, n_2021, n_2025, n_3010, n_2160, n_1992, n_124, n_3744, n_4015, n_2924, n_307, n_1209, n_4022, n_1020, n_1563, n_3673, n_3052, n_646, n_2507, n_3438, n_2142, n_1633, n_34, n_404, n_2625, n_2896, n_172, n_1913, n_2069, n_2495, n_3187, n_1058, n_2328, n_4043, n_347, n_2434, n_1042, n_3170, n_183, n_1234, n_2311, n_479, n_3936, n_1578, n_2261, n_1455, n_3147, n_2287, n_299, n_836, n_2223, n_3082, n_1279, n_3415, n_3661, n_2473, n_3320, n_2144, n_2511, n_3464, n_564, n_3414, n_133, n_66, n_205, n_1029, n_2649, n_3981, n_1247, n_760, n_522, n_2438, n_1568, n_2919, n_20, n_3210, n_1483, n_3108, n_1363, n_2681, n_3867, n_3397, n_367, n_1111, n_970, n_1689, n_2535, n_3467, n_713, n_1255, n_2632, n_1646, n_598, n_3031, n_345, n_2262, n_3179, n_2565, n_3889, n_1237, n_3262, n_927, n_261, n_1095, n_2980, n_1728, n_2335, n_3078, n_3699, n_3971, n_370, n_706, n_2120, n_286, n_3239, n_2631, n_3215, n_3311, n_3869, n_3516, n_1401, n_1419, n_3138, n_1531, n_776, n_424, n_2860, n_3816, n_2041, n_2113, n_1933, n_3528, n_1651, n_3087, n_85, n_130, n_2697, n_1387, n_466, n_1263, n_346, n_1817, n_3711, n_2404, n_2168, n_2757, n_3704, n_348, n_552, n_2312, n_670, n_2677, n_1826, n_3171, n_379, n_138, n_162, n_264, n_3577, n_2834, n_4051, n_2483, n_4074, n_3994, n_441, n_1951, n_3185, n_2490, n_1032, n_1217, n_2558, n_1496, n_2996, n_637, n_1592, n_2812, n_3660, n_73, n_327, n_2662, n_1259, n_3300, n_2801, n_1177, n_3104, n_3074, n_2655, n_1231, n_3917, n_4122, n_3246, n_2132, n_3299, n_980, n_1618, n_3774, n_1869, n_3589, n_3623, n_1743, n_905, n_2718, n_207, n_720, n_926, n_41, n_1943, n_2687, n_2296, n_3876, n_3615, n_3267, n_194, n_1802, n_2178, n_3946, n_2112, n_2765, n_1163, n_2640, n_3054, n_2811, n_3019, n_186, n_1795, n_3200, n_1384, n_3642, n_2237, n_145, n_2146, n_2983, n_1868, n_3276, n_59, n_3601, n_4089, n_1501, n_2241, n_2373, n_1173, n_3498, n_3513, n_3682, n_2350, n_3881, n_1068, n_1198, n_4096, n_2531, n_1570, n_2099, n_3759, n_3377, n_487, n_1518, n_3323, n_1456, n_4007, n_90, n_1879, n_1886, n_1648, n_2187, n_3961, n_1413, n_2617, n_2481, n_3863, n_2129, n_855, n_2327, n_158, n_3882, n_3916, n_808, n_1365, n_2476, n_553, n_2814, n_2059, n_3675, n_3968, n_2437, n_2636, n_1439, n_814, n_578, n_3466, n_2074, n_1665, n_1287, n_2841, n_405, n_1611, n_2122, n_120, n_3572, n_2975, n_3332, n_2399, n_320, n_1414, n_1134, n_2067, n_3374, n_3471, n_4075, n_1484, n_1901, n_647, n_2055, n_2998, n_3465, n_2027, n_2932, n_1423, n_2117, n_481, n_600, n_1053, n_1609, n_3118, n_4072, n_2822, n_1939, n_2308, n_2242, n_1906, n_529, n_1899, n_3039, n_2195, n_3922, n_502, n_2194, n_2937, n_218, n_3508, n_1467, n_4039, n_247, n_1828, n_2159, n_1798, n_3057, n_1304, n_1608, n_3831, n_1744, n_3335, n_3007, n_2267, n_1105, n_547, n_3599, n_3618, n_439, n_604, n_677, n_3705, n_3022, n_478, n_703, n_3983, n_1349, n_1709, n_3318, n_1061, n_3385, n_2102, n_326, n_681, n_3477, n_227, n_3286, n_3734, n_3370, n_874, n_3773, n_3949, n_2286, n_3494, n_2023, n_1278, n_707, n_3974, n_3443, n_11, n_3401, n_129, n_126, n_983, n_3036, n_2783, n_2599, n_3988, n_3788, n_3939, n_590, n_699, n_727, n_301, n_1726, n_2075, n_3263, n_3542, n_2523, n_1945, n_3569, n_3835, n_3837, n_545, n_1015, n_2418, n_1377, n_1162, n_536, n_1614, n_2031, n_2496, n_3260, n_3349, n_3761, n_3819, n_3996, n_2118, n_325, n_1740, n_3222, n_1602, n_688, n_3139, n_636, n_2853, n_427, n_3350, n_3801, n_1098, n_3009, n_1490, n_2338, n_442, n_777, n_3764, n_1553, n_1080, n_920, n_1760, n_1086, n_1092, n_3025, n_3636, n_3051, n_3205, n_2225, n_986, n_1104, n_1963, n_2802, n_3653, n_3951, n_3868, n_3035, n_3823, n_729, n_887, n_3403, n_2057, n_2218, n_1122, n_1205, n_1408, n_2593, n_163, n_1693, n_2125, n_2716, n_1132, n_390, n_1156, n_2741, n_501, n_2184, n_2714, n_314, n_1823, n_2944, n_2861, n_2780, n_3023, n_1120, n_3439, n_3942, n_1202, n_4084, n_627, n_2254, n_3130, n_3290, n_1188, n_1498, n_1371, n_2033, n_2618, n_4121, n_3602, n_233, n_957, n_388, n_1402, n_1242, n_3957, n_2754, n_2707, n_2774, n_3418, n_2849, n_1607, n_1489, n_2799, n_1218, n_2756, n_3611, n_3781, n_2217, n_221, n_321, n_86, n_2226, n_3959, n_3984, n_1586, n_861, n_3338, n_2962, n_1543, n_1431, n_877, n_3995, n_1119, n_3713, n_1863, n_1763, n_1666, n_3908, n_1500, n_616, n_2214, n_1055, n_1395, n_3892, n_1346, n_2763, n_3156, n_2256, n_1189, n_3337, n_1089, n_3750, n_3424, n_281, n_3326, n_3356, n_1859, n_2660, n_3426, n_262, n_1502, n_3044, n_1523, n_2190, n_3492, n_3501, n_1478, n_2732, n_1883, n_3737, n_2516, n_3931, n_4094, n_2776, n_2555, n_3216, n_3224, n_3568, n_1969, n_2708, n_735, n_297, n_3070, n_1005, n_3275, n_527, n_2379, n_46, n_3579, n_3245, n_84, n_1294, n_2661, n_1667, n_845, n_888, n_2894, n_2300, n_2949, n_3896, n_4049, n_4067, n_1649, n_2452, n_1677, n_2470, n_1927, n_1297, n_2827, n_178, n_3214, n_551, n_3551, n_417, n_1708, n_70, n_343, n_3085, n_3373, n_1222, n_2284, n_3005, n_3710, n_1844, n_2283, n_582, n_2526, n_1957, n_3364, n_1953, n_2643, n_755, n_1097, n_3803, n_3766, n_3985, n_1219, n_1711, n_710, n_1919, n_2994, n_534, n_1791, n_2508, n_3186, n_2124, n_1894, n_1460, n_1239, n_2594, n_3826, n_278, n_2266, n_3944, n_3417, n_2449, n_560, n_890, n_842, n_148, n_3626, n_1898, n_451, n_745, n_1741, n_1572, n_1907, n_1793, n_3180, n_3648, n_3423, n_61, n_742, n_1081, n_1373, n_1975, n_1388, n_1266, n_1540, n_1719, n_2119, n_2742, n_769, n_3671, n_1797, n_2366, n_2493, n_13, n_1753, n_1990, n_1372, n_476, n_832, n_55, n_535, n_744, n_1895, n_2821, n_3491, n_2690, n_3090, n_3696, n_2474, n_4104, n_2623, n_3392, n_982, n_1800, n_915, n_215, n_3791, n_1075, n_2008, n_454, n_298, n_1331, n_1890, n_2904, n_3064, n_3199, n_4034, n_1529, n_3353, n_1227, n_3531, n_2127, n_655, n_2946, n_3166, n_3151, n_3649, n_3684, n_3333, n_3512, n_1734, n_1860, n_3065, n_403, n_3016, n_2785, n_2460, n_4114, n_2840, n_1007, n_1580, n_1319, n_3135, n_657, n_3367, n_3669, n_3956, n_3924, n_4081, n_837, n_812, n_2448, n_3997, n_2211, n_4040, n_2292, n_2480, n_606, n_951, n_3024, n_2772, n_3564, n_862, n_1700, n_2637, n_659, n_1332, n_3795, n_2306, n_509, n_1854, n_666, n_1747, n_2071, n_2424, n_3990, n_430, n_1206, n_1729, n_722, n_1508, n_3953, n_2414, n_2082, n_2893, n_2959, n_1532, n_3277, n_1171, n_1030, n_785, n_3161, n_3208, n_2389, n_4069, n_1309, n_3582, n_999, n_2280, n_1766, n_1338, n_2978, n_1342, n_2737, n_3282, n_456, n_1867, n_3993, n_852, n_1394, n_2916, n_2576, n_3459, n_3617, n_704, n_2958, n_3365, n_1060, n_1044, n_1714, n_4113, n_2696, n_3340, n_521, n_2140, n_873, n_1301, n_1748, n_2157, n_1966, n_1243, n_2171, n_2468, n_3977, n_1400, n_4112, n_342, n_3400, n_2035, n_2614, n_1466, n_3735, n_3486, n_1513, n_1527, n_2581, n_358, n_1783, n_3656, n_608, n_2494, n_1538, n_2831, n_2457, n_2128, n_3069, n_2992, n_1037, n_3650, n_4071, n_1329, n_317, n_3197, n_1993, n_1545, n_3586, n_134, n_2629, n_3369, n_4035, n_3256, n_1257, n_1480, n_1954, n_3670, n_1668, n_1878, n_3964, n_2540, n_3836, n_3302, n_1605, n_1078, n_3060, n_266, n_2486, n_1897, n_2984, n_4009, n_157, n_3646, n_2520, n_2137, n_1161, n_2489, n_3685, n_811, n_3097, n_624, n_3507, n_791, n_876, n_618, n_1191, n_2492, n_3864, n_2939, n_3425, n_736, n_1025, n_1215, n_241, n_1449, n_3450, n_3748, n_2337, n_2265, n_687, n_2900, n_797, n_2026, n_2912, n_3524, n_1786, n_2627, n_4050, n_3173, n_480, n_1327, n_3732, n_1475, n_211, n_642, n_1804, n_2106, n_97, n_408, n_1406, n_595, n_1405, n_2684, n_3174, n_3314, n_2726, n_602, n_3813, n_2622, n_3447, n_4006, n_2272, n_3266, n_1757, n_592, n_3102, n_1499, n_854, n_1318, n_3452, n_2091, n_393, n_1632, n_1769, n_474, n_1929, n_4098, n_1950, n_2264, n_2691, n_3789, n_805, n_2032, n_2090, n_2929, n_3124, n_3811, n_3422, n_295, n_1658, n_190, n_2249, n_1072, n_3411, n_695, n_1526, n_2991, n_3463, n_1305, n_64, n_180, n_730, n_386, n_1596, n_2348, n_2656, n_1281, n_516, n_2364, n_1997, n_2574, n_1137, n_1873, n_1258, n_197, n_640, n_463, n_1476, n_1524, n_1733, n_1856, n_2016, n_2667, n_2723, n_2725, n_3925, n_2928, n_943, n_1118, n_678, n_2905, n_2884, n_3408, n_651, n_2850, n_1874, n_1293, n_3167, n_3746, n_961, n_469, n_1046, n_1807, n_726, n_1123, n_3780, n_1657, n_878, n_2857, n_3694, n_4118, n_1784, n_3110, n_3857, n_771, n_3787, n_4025, n_1321, n_3050, n_3919, n_3157, n_3753, n_3893, n_752, n_2307, n_71, n_1488, n_985, n_421, n_1330, n_906, n_3702, n_1180, n_1697, n_2295, n_2730, n_283, n_4076, n_806, n_3142, n_1984, n_1350, n_3453, n_3129, n_1556, n_649, n_1561, n_2412, n_2720, n_374, n_3298, n_3107, n_3495, n_1352, n_3843, n_2405, n_2815, n_1824, n_643, n_2606, n_2700, n_1492, n_226, n_4065, n_2383, n_2764, n_1441, n_1822, n_682, n_36, n_1616, n_2633, n_2416, n_3708, n_819, n_2386, n_2907, n_1971, n_2945, n_586, n_1324, n_1429, n_2064, n_2353, n_2528, n_1778, n_3543, n_3640, n_1776, n_3448, n_686, n_605, n_2936, n_1154, n_584, n_3609, n_1557, n_1759, n_1829, n_2325, n_1130, n_1450, n_3718, n_349, n_756, n_2022, n_3390, n_1016, n_2298, n_1149, n_1505, n_2408, n_2698, n_3740, n_2986, n_2320, n_3017, n_979, n_2329, n_2570, n_3140, n_1642, n_2417, n_2789, n_2, n_3976, n_2525, n_1815, n_2813, n_897, n_2546, n_949, n_2454, n_1493, n_2890, n_2911, n_515, n_3381, n_807, n_3455, n_3736, n_891, n_3313, n_885, n_1659, n_3955, n_2354, n_3591, n_198, n_1864, n_2760, n_3907, n_3086, n_1887, n_3165, n_1208, n_3317, n_3945, n_3726, n_3336, n_1987, n_4052, n_3357, n_3388, n_396, n_2368, n_802, n_23, n_1151, n_554, n_960, n_3635, n_2352, n_3541, n_2502, n_1256, n_87, n_714, n_3560, n_3345, n_2170, n_3605, n_790, n_2244, n_2143, n_2393, n_354, n_140, n_725, n_2377, n_1577, n_3566, n_151, n_3840, n_3421, n_1448, n_2198, n_28, n_1009, n_230, n_3548, n_2652, n_1133, n_3067, n_154, n_883, n_142, n_4097, n_4054, n_3809, n_473, n_1852, n_801, n_1286, n_2612, n_818, n_1685, n_779, n_2410, n_2314, n_2477, n_2279, n_3169, n_594, n_3236, n_2222, n_3468, n_1995, n_1877, n_1397, n_35, n_1052, n_272, n_1333, n_1306, n_1849, n_3573, n_2076, n_2133, n_2203, n_833, n_2943, n_1426, n_2250, n_3319, n_2497, n_2247, n_2230, n_879, n_1117, n_3321, n_38, n_422, n_1269, n_1303, n_1547, n_1438, n_1541, n_597, n_3291, n_3654, n_75, n_2001, n_1047, n_3783, n_95, n_2506, n_1472, n_2413, n_4008, n_1593, n_2610, n_3715, n_1050, n_2626, n_566, n_2158, n_2578, n_2607, n_3643, n_2285, n_3343, n_3184, n_152, n_3309, n_2892, n_169, n_106, n_1201, n_1288, n_173, n_2605, n_858, n_2796, n_1185, n_2475, n_2804, n_2173, n_3982, n_2715, n_3206, n_335, n_3647, n_1035, n_3475, n_1143, n_2665, n_344, n_2070, n_2136, n_426, n_433, n_3973, n_3134, n_398, n_2771, n_62, n_210, n_1090, n_2403, n_3755, n_2947, n_1367, n_3842, n_2044, n_166, n_253, n_928, n_3886, n_1153, n_271, n_465, n_3769, n_4078, n_825, n_1103, n_732, n_2619, n_1565, n_1192, n_128, n_224, n_3738, n_82, n_894, n_3098, n_1380, n_1624, n_1801, n_2854, n_3055, n_420, n_1291, n_562, n_4070, n_2020, n_748, n_3987, n_2310, n_510, n_1045, n_256, n_3341, n_3600, n_3160, n_1160, n_2968, n_1882, n_1976, n_1023, n_2711, n_3223, n_1881, n_2635, n_2999, n_988, n_3386, n_330, n_914, n_400, n_689, n_1116, n_3921, n_282, n_328, n_368, n_3043, n_3190, n_1958, n_2747, n_3667, n_3027, n_4011, n_467, n_1511, n_2177, n_3695, n_2713, n_1422, n_3800, n_2766, n_1965, n_644, n_3462, n_1197, n_3906, n_3011, n_3395, n_276, n_2820, n_2613, n_3226, n_497, n_3733, n_1165, n_3378, n_2934, n_1641, n_3967, n_3731, n_168, n_81, n_538, n_2845, n_1517, n_2036, n_576, n_843, n_511, n_2647, n_455, n_429, n_588, n_3358, n_638, n_2003, n_2533, n_2210, n_3920, n_1307, n_3444, n_1128, n_3141, n_2053, n_3851, n_4091, n_1671, n_1417, n_3476, n_1048, n_2343, n_775, n_3096, n_667, n_2419, n_1049, n_3380, n_2330, n_2826, n_14, n_869, n_141, n_846, n_1398, n_1921, n_2777, n_3238, n_2450, n_2411, n_1356, n_1341, n_2234, n_2309, n_3189, n_3233, n_1504, n_1955, n_2110, n_2431, n_1773, n_3175, n_1440, n_3289, n_2666, n_3322, n_1370, n_1603, n_305, n_312, n_56, n_60, n_728, n_413, n_2401, n_2935, n_715, n_889, n_3822, n_3255, n_3818, n_1066, n_1549, n_2588, n_2863, n_2331, n_935, n_2886, n_3827, n_2478, n_685, n_911, n_4061, n_361, n_89, n_2658, n_623, n_3509, n_3587, n_2608, n_3620, n_2920, n_1712, n_3344, n_1403, n_1065, n_453, n_1534, n_1948, n_3006, n_74, n_2767, n_810, n_3376, n_19, n_40, n_1290, n_181, n_1959, n_3497, n_617, n_3770, n_2396, n_3243, n_543, n_3368, n_1362, n_1559, n_2121, n_3456, n_3865, n_3123, n_2692, n_236, n_601, n_683, n_565, n_3927, n_628, n_1300, n_1960, n_4102, n_2068, n_3117, n_3595, n_743, n_1194, n_2862, n_4060, n_1647, n_1546, n_3384, n_1420, n_2553, n_2645, n_3790, n_907, n_2749, n_1454, n_2592, n_660, n_464, n_3490, n_2459, n_962, n_941, n_3396, n_1210, n_847, n_747, n_1622, n_1135, n_2566, n_2751, n_3113, n_3101, n_918, n_1968, n_3307, n_107, n_3662, n_1885, n_639, n_452, n_673, n_3251, n_3288, n_4093, n_2842, n_2833, n_2196, n_1038, n_3603, n_3723, n_2371, n_1978, n_414, n_571, n_3880, n_3720, n_1521, n_1694, n_1940, n_3683, n_6, n_284, n_3904, n_3887, n_593, n_3195, n_3008, n_1695, n_3242, n_4027, n_2560, n_1164, n_3405, n_37, n_58, n_2313, n_609, n_3077, n_1193, n_3048, n_3339, n_1345, n_613, n_3037, n_1022, n_1336, n_1033, n_3478, n_3062, n_1774, n_409, n_171, n_2963, n_3532, n_519, n_384, n_2609, n_2561, n_1166, n_1056, n_2007, n_526, n_1994, n_3363, n_3533, n_3978, n_1767, n_1040, n_674, n_3131, n_1158, n_316, n_3168, n_125, n_1973, n_1444, n_1803, n_820, n_1749, n_43, n_872, n_1653, n_3409, n_4079, n_3522, n_3583, n_4088, n_254, n_2882, n_2303, n_2669, n_3540, n_3911, n_3241, n_3802, n_3899, n_1157, n_1584, n_234, n_848, n_1664, n_3481, n_280, n_629, n_3563, n_1739, n_161, n_2642, n_3310, n_1814, n_532, n_3689, n_2154, n_2441, n_2236, n_1789, n_763, n_1986, n_4041, n_2174, n_2688, n_99, n_540, n_216, n_692, n_2624, n_5, n_3442, n_3972, n_2054, n_1857, n_2315, n_3926, n_984, n_1687, n_2073, n_223, n_2150, n_4004, n_1552, n_750, n_2938, n_834, n_3630, n_1612, n_2498, n_800, n_2638, n_3992, n_2046, n_1816, n_1910, n_2803, n_1756, n_2887, n_1606, n_2189, n_395, n_621, n_2648, n_3305, n_1587, n_213, n_3810, n_4062, n_2093, n_2340, n_2018, n_2672, n_1772, n_67, n_2444, n_2602, n_3354, n_1014, n_724, n_2204, n_2931, n_3433, n_1427, n_1481, n_2040, n_493, n_1311, n_2977, n_3106, n_3597, n_3991, n_2199, n_2881, n_1956, n_1589, n_114, n_4111, n_2151, n_1100, n_585, n_875, n_1617, n_2455, n_827, n_2600, n_3092, n_3437, n_2231, n_3786, n_697, n_2828, n_622, n_1626, n_3436, n_1962, n_1335, n_1715, n_3806, n_296, n_3553, n_4044, n_2305, n_3645, n_880, n_793, n_2114, n_3329, n_2927, n_3304, n_3833, n_3574, n_1175, n_2289, n_132, n_2530, n_2299, n_3751, n_3402, n_751, n_1027, n_1070, n_2406, n_3247, n_1621, n_4110, n_739, n_1485, n_1028, n_2883, n_1221, n_530, n_1785, n_792, n_1262, n_1942, n_2180, n_3406, n_2951, n_3807, n_4048, n_580, n_3664, n_1579, n_494, n_2809, n_2181, n_3550, n_434, n_2014, n_975, n_2974, n_229, n_394, n_923, n_1645, n_1124, n_1381, n_2870, n_1494, n_932, n_1893, n_1183, n_3686, n_3722, n_1326, n_2889, n_2276, n_3969, n_1805, n_2282, n_3301, n_981, n_4068, n_2910, n_2141, n_1110, n_1758, n_2503, n_3873, n_2270, n_3470, n_243, n_3785, n_3294, n_2443, n_1407, n_185, n_2465, n_3610, n_1204, n_2865, n_1554, n_3279, n_994, n_2428, n_2972, n_2586, n_2989, n_1360, n_973, n_3178, n_2858, n_268, n_972, n_3844, n_3259, n_2251, n_2923, n_3076, n_164, n_2843, n_3714, n_184, n_3410, n_856, n_3100, n_2572, n_1248, n_1176, n_3721, n_3676, n_1564, n_2010, n_3677, n_1054, n_508, n_118, n_121, n_1679, n_3292, n_3389, n_2872, n_2126, n_3701, n_3109, n_3706, n_1952, n_2425, n_2394, n_3989, n_1858, n_353, n_3125, n_1678, n_2589, n_4086, n_1482, n_1361, n_2356, n_1601, n_3537, n_1057, n_191, n_2487, n_1834, n_978, n_1011, n_1520, n_2534, n_2488, n_1509, n_828, n_2941, n_322, n_1411, n_1359, n_3079, n_3638, n_3269, n_558, n_3536, n_1721, n_2564, n_116, n_3558, n_3576, n_3782, n_39, n_2591, n_653, n_1445, n_1317, n_3034, n_2050, n_2197, n_3502, n_3248, n_783, n_4053, n_2550, n_556, n_1127, n_170, n_1536, n_3177, n_3594, n_1471, n_2385, n_160, n_3440, n_119, n_2387, n_1008, n_3963, n_332, n_3658, n_581, n_294, n_3091, n_1024, n_830, n_176, n_3404, n_2291, n_3346, n_2816, n_1980, n_2518, n_987, n_936, n_2510, n_1620, n_2501, n_2542, n_3227, n_3570, n_3105, n_1385, n_1525, n_2793, n_1998, n_2165, n_2675, n_541, n_499, n_2604, n_1775, n_788, n_12, n_908, n_2639, n_3521, n_3855, n_1036, n_2169, n_2985, n_2603, n_341, n_4083, n_1270, n_109, n_1167, n_1272, n_549, n_2630, n_591, n_4105, n_2794, n_969, n_3663, n_2028, n_919, n_1663, n_50, n_3114, n_2901, n_2092, n_3940, n_2175, n_1625, n_2086, n_3225, n_3622, n_2773, n_2817, n_1926, n_2402, n_3621, n_318, n_1458, n_103, n_244, n_679, n_1630, n_3473, n_220, n_3644, n_3047, n_663, n_1720, n_2409, n_2966, n_3163, n_3680, n_443, n_3431, n_2176, n_3565, n_1412, n_3355, n_3059, n_1738, n_1550, n_528, n_1358, n_1200, n_387, n_406, n_826, n_3897, n_139, n_2808, n_2453, n_2344, n_1922, n_3331, n_1735, n_1788, n_391, n_940, n_3520, n_2392, n_1537, n_2138, n_4005, n_3272, n_3122, n_3040, n_2065, n_2543, n_2321, n_1077, n_2597, n_607, n_956, n_445, n_3360, n_1930, n_3687, n_765, n_1809, n_2787, n_4092, n_3585, n_1843, n_1904, n_122, n_2000, n_3799, n_3133, n_2805, n_4037, n_1268, n_3804, n_2676, n_2758, n_385, n_3211, n_2395, n_917, n_2868, n_1271, n_372, n_2096, n_2440, n_2556, n_2186, n_15, n_1530, n_2215, n_4057, n_2770, n_631, n_399, n_3847, n_1170, n_2724, n_4073, n_3575, n_2258, n_1261, n_2471, n_702, n_3633, n_857, n_898, n_3042, n_363, n_968, n_1067, n_1235, n_1323, n_2584, n_2375, n_3278, n_1462, n_3328, n_4001, n_1937, n_2012, n_3182, n_2967, n_3608, n_1064, n_633, n_900, n_1446, n_1282, n_3004, n_1701, n_1093, n_1551, n_2039, n_1755, n_4021, n_1285, n_3379, n_3111, n_193, n_733, n_761, n_2212, n_3838, n_731, n_336, n_1813, n_315, n_2268, n_2997, n_3469, n_4059, n_311, n_1452, n_2835, n_1573, n_3258, n_2734, n_8, n_668, n_2569, n_758, n_4019, n_3691, n_2252, n_3598, n_2111, n_3743, n_2420, n_2948, n_3099, n_1996, n_1106, n_2009, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_2897, n_1322, n_3273, n_3829, n_2583, n_2918, n_2987, n_1473, n_835, n_3155, n_446, n_1076, n_2024, n_1348, n_2651, n_753, n_2445, n_2733, n_1770, n_701, n_1003, n_2469, n_1125, n_2103, n_4024, n_2358, n_3316, n_4023, n_1710, n_1865, n_2522, n_2641, n_3632, n_2463, n_3546, n_309, n_1344, n_115, n_2355, n_1390, n_2580, n_2699, n_401, n_485, n_1792, n_4064, n_504, n_3351, n_2062, n_483, n_435, n_3068, n_1141, n_3457, n_1629, n_3901, n_291, n_1640, n_822, n_1094, n_2973, n_840, n_1459, n_2153, n_2324, n_1510, n_3454, n_3002, n_2710, n_2505, n_2139, n_1099, n_839, n_79, n_1754, n_3, n_3146, n_3394, n_3038, n_759, n_567, n_2397, n_91, n_2521, n_240, n_369, n_1727, n_2740, n_2235, n_44, n_1991, n_1575, n_3693, n_3878, n_2721, n_1848, n_1892, n_1172, n_3132, n_2615, n_614, n_3776, n_4066, n_2775, n_3903, n_1212, n_3581, n_3778, n_831, n_3681, n_3933, n_3970, n_778, n_48, n_1619, n_2351, n_3303, n_188, n_2260, n_323, n_550, n_1315, n_1660, n_4080, n_1902, n_997, n_635, n_2206, n_2784, n_3898, n_2541, n_694, n_1643, n_1320, n_3188, n_3001, n_3232, n_1113, n_3218, n_2347, n_248, n_3768, n_1152, n_2657, n_2990, n_2447, n_2034, n_1845, n_2538, n_3932, n_1934, n_2101, n_2577, n_921, n_2362, n_1615, n_1236, n_4100, n_228, n_2104, n_1265, n_1576, n_2105, n_1470, n_671, n_1533, n_1806, n_2372, n_2552, n_3445, n_4087, n_1, n_1409, n_1148, n_1588, n_1684, n_1673, n_2422, n_2704, n_1334, n_654, n_2290, n_2933, n_3729, n_3253, n_2856, n_3235, n_3387, n_2088, n_3265, n_3952, n_1275, n_3103, n_488, n_3018, n_904, n_505, n_88, n_2005, n_3584, n_2048, n_1696, n_3446, n_498, n_3028, n_1875, n_1059, n_3148, n_3775, n_684, n_2429, n_2108, n_2736, n_3966, n_3285, n_3824, n_3825, n_1039, n_2246, n_3616, n_539, n_1150, n_977, n_449, n_2339, n_3846, n_392, n_1628, n_1289, n_1831, n_2532, n_2191, n_2971, n_3874, n_1497, n_1866, n_2472, n_2664, n_2705, n_2056, n_2852, n_459, n_1136, n_2515, n_3845, n_1782, n_458, n_1190, n_1600, n_1144, n_3203, n_383, n_838, n_1558, n_4107, n_1941, n_3628, n_1316, n_175, n_2519, n_3637, n_950, n_1017, n_711, n_3941, n_734, n_1915, n_2360, n_723, n_1393, n_2240, n_658, n_630, n_1369, n_53, n_362, n_2846, n_310, n_3371, n_1781, n_709, n_2917, n_3137, n_2544, n_24, n_809, n_3143, n_3194, n_3690, n_2085, n_2432, n_3229, n_3032, n_3872, n_1686, n_1964, n_3659, n_3928, n_235, n_881, n_1019, n_1477, n_1777, n_2188, n_1982, n_2097, n_662, n_641, n_3366, n_3461, n_2430, n_2504, n_910, n_290, n_741, n_939, n_1410, n_2297, n_3094, n_3441, n_371, n_199, n_3020, n_4002, n_217, n_2964, n_1114, n_1325, n_1742, n_708, n_308, n_1223, n_3815, n_2545, n_201, n_1768, n_2513, n_2193, n_2369, n_572, n_1199, n_2957, n_865, n_10, n_1273, n_1983, n_2982, n_1041, n_2451, n_3312, n_2115, n_2913, n_993, n_1862, n_948, n_2017, n_3752, n_3672, n_922, n_1004, n_1810, n_3061, n_448, n_2587, n_3504, n_1347, n_2839, n_3237, n_860, n_3555, n_3820, n_3072, n_1043, n_2961, n_255, n_2869, n_3534, n_450, n_4036, n_1923, n_3848, n_3655, n_2955, n_2670, n_3631, n_1764, n_2674, n_3556, n_896, n_1737, n_1479, n_1613, n_3026, n_2644, n_902, n_1031, n_2979, n_1723, n_3674, n_1638, n_853, n_3071, n_3918, n_716, n_4010, n_1571, n_1698, n_3902, n_4101, n_196, n_3866, n_1337, n_3763, n_774, n_1946, n_2148, n_933, n_3244, n_3499, n_1779, n_2562, n_596, n_954, n_2051, n_3112, n_1168, n_1821, n_4095, n_219, n_1310, n_3296, n_3196, n_3762, n_3794, n_231, n_3910, n_3947, n_656, n_492, n_574, n_3593, n_2673, n_252, n_664, n_1591, n_2585, n_2995, n_3293, n_3361, n_1229, n_1683, n_2582, n_3228, n_3327, n_2548, n_68, n_3488, n_1896, n_2164, n_1732, n_415, n_2381, n_2744, n_1967, n_2384, n_2678, n_2179, n_63, n_1280, n_544, n_1516, n_1186, n_1705, n_599, n_768, n_3707, n_1091, n_2052, n_2485, n_3779, n_3895, n_3149, n_537, n_1063, n_3934, n_25, n_991, n_2183, n_2205, n_83, n_2275, n_389, n_2563, n_1724, n_3088, n_1670, n_1707, n_1799, n_2080, n_3590, n_2058, n_3231, n_1126, n_3834, n_2761, n_2357, n_2029, n_195, n_1846, n_1912, n_3923, n_938, n_1891, n_1328, n_895, n_110, n_304, n_2875, n_1639, n_583, n_3519, n_2209, n_2421, n_1302, n_3295, n_1000, n_313, n_626, n_4042, n_378, n_1581, n_3849, n_1928, n_98, n_946, n_757, n_2047, n_3058, n_375, n_113, n_1655, n_1818, n_33, n_1146, n_2792, n_3398, n_3709, n_1634, n_2596, n_1203, n_998, n_1699, n_1598, n_3557, n_3592, n_3725, n_3986, n_2269, n_472, n_937, n_1474, n_2081, n_4026, n_2536, n_2524, n_265, n_1583, n_1604, n_208, n_1631, n_1702, n_3399, n_3894, n_156, n_174, n_275, n_100, n_3202, n_1794, n_1375, n_3053, n_147, n_204, n_1232, n_996, n_1211, n_1368, n_963, n_3772, n_1264, n_51, n_1082, n_1725, n_496, n_2891, n_2318, n_1827, n_3128, n_4120, n_866, n_26, n_246, n_925, n_1752, n_1313, n_1001, n_1722, n_2361, n_1115, n_2229, n_2819, n_2880, n_3030, n_3075, n_3505, n_1339, n_1002, n_1644, n_105, n_1051, n_3547, n_4014, n_3771, n_2551, n_719, n_131, n_263, n_1102, n_360, n_2255, n_1129, n_1252, n_2239, n_3045, n_250, n_1464, n_1296, n_3158, n_773, n_2798, n_3221, n_2316, n_165, n_3217, n_2464, n_3697, n_1010, n_2830, n_882, n_2706, n_2304, n_1249, n_101, n_803, n_1871, n_2514, n_329, n_718, n_3821, n_1434, n_340, n_1905, n_1569, n_3201, n_3334, n_4016, n_2573, n_2940, n_3503, n_289, n_9, n_112, n_45, n_548, n_3427, n_2336, n_523, n_1662, n_3162, n_457, n_1299, n_1870, n_3249, n_3430, n_3483, n_4046, n_177, n_2063, n_1925, n_782, n_364, n_258, n_2915, n_3489, n_3083, n_431, n_2654, n_3935, n_2491, n_1861, n_2079, n_1228, n_2319, n_2152, n_3213, n_2517, n_1931, n_4047, n_1244, n_3484, n_1796, n_411, n_484, n_2259, n_849, n_2095, n_2719, n_22, n_2965, n_2738, n_1820, n_2590, n_2876, n_2797, n_29, n_357, n_412, n_1251, n_1989, n_3041, n_447, n_1421, n_2208, n_2423, n_2689, n_4063, n_2778, n_1762, n_1233, n_3798, n_3080, n_1808, n_1574, n_1672, n_2228, n_1635, n_3033, n_1704, n_3832, n_893, n_3525, n_3308, n_3712, n_1582, n_841, n_2479, n_3204, n_886, n_1069, n_1981, n_2824, n_2037, n_2953, n_359, n_3428, n_1308, n_573, n_796, n_2851, n_2823, n_4017, n_127, n_531, n_2345, n_1730, n_1374, n_1451, n_2089, n_1487, n_675, n_16275);

input n_2752;
input n_3527;
input n_913;
input n_1681;
input n_2163;
input n_3432;
input n_4030;
input n_1486;
input n_1507;
input n_1938;
input n_3619;
input n_589;
input n_2484;
input n_2866;
input n_3153;
input n_1174;
input n_4013;
input n_3152;
input n_2346;
input n_3434;
input n_1469;
input n_691;
input n_1353;
input n_3056;
input n_3500;
input n_3480;
input n_2679;
input n_1355;
input n_2131;
input n_3268;
input n_3853;
input n_2559;
input n_2500;
input n_2509;
input n_423;
input n_4085;
input n_1383;
input n_2182;
input n_603;
input n_373;
input n_2135;
input n_2334;
input n_2680;
input n_3264;
input n_1250;
input n_2030;
input n_1169;
input n_789;
input n_3181;
input n_850;
input n_2993;
input n_1916;
input n_2879;
input n_610;
input n_245;
input n_1713;
input n_96;
input n_319;
input n_49;
input n_1436;
input n_2407;
input n_690;
input n_2818;
input n_416;
input n_3578;
input n_1109;
input n_1430;
input n_2537;
input n_525;
input n_187;
input n_3745;
input n_2002;
input n_1463;
input n_2243;
input n_3487;
input n_1238;
input n_2694;
input n_3668;
input n_2011;
input n_3742;
input n_2729;
input n_1515;
input n_817;
input n_1837;
input n_924;
input n_781;
input n_2013;
input n_2786;
input n_1566;
input n_2837;
input n_189;
input n_717;
input n_3765;
input n_72;
input n_2006;
input n_4058;
input n_952;
input n_864;
input n_4090;
input n_2446;
input n_1096;
input n_4116;
input n_1379;
input n_2436;
input n_57;
input n_3352;
input n_3517;
input n_2376;
input n_2367;
input n_2671;
input n_2790;
input n_1706;
input n_2207;
input n_2461;
input n_2702;
input n_3719;
input n_117;
input n_524;
input n_2731;
input n_3703;
input n_1214;
input n_634;
input n_3561;
input n_1839;
input n_1246;
input n_1138;
input n_214;
input n_3526;
input n_3888;
input n_3954;
input n_2042;
input n_2123;
input n_3198;
input n_1853;
input n_764;
input n_1503;
input n_2238;
input n_2529;
input n_2374;
input n_4103;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_1999;
input n_3435;
input n_410;
input n_2380;
input n_1187;
input n_1131;
input n_1225;
input n_3154;
input n_2646;
input n_737;
input n_137;
input n_1298;
input n_2653;
input n_1745;
input n_2873;
input n_1366;
input n_232;
input n_52;
input n_2084;
input n_3115;
input n_3938;
input n_568;
input n_2278;
input n_4028;
input n_3330;
input n_3514;
input n_1088;
input n_77;
input n_1424;
input n_766;
input n_2976;
input n_1835;
input n_3383;
input n_3965;
input n_1457;
input n_377;
input n_2482;
input n_3905;
input n_1682;
input n_2750;
input n_3797;
input n_1836;
input n_3416;
input n_520;
input n_870;
input n_2547;
input n_3382;
input n_1453;
input n_279;
input n_945;
input n_958;
input n_3943;
input n_3930;
input n_2554;
input n_3145;
input n_3808;
input n_2248;
input n_3665;
input n_3063;
input n_813;
input n_3281;
input n_3535;
input n_419;
input n_1985;
input n_2288;
input n_2621;
input n_2908;
input n_3081;
input n_146;
input n_3858;
input n_270;
input n_4106;
input n_338;
input n_995;
input n_2579;
input n_285;
input n_1909;
input n_2156;
input n_1184;
input n_1961;
input n_202;
input n_1535;
input n_3220;
input n_2960;
input n_500;
input n_665;
input n_754;
input n_903;
input n_3270;
input n_871;
input n_2323;
input n_1073;
input n_2844;
input n_3348;
input n_239;
input n_402;
input n_1979;
input n_1277;
input n_2107;
input n_1746;
input n_3261;
input n_54;
input n_829;
input n_1761;
input n_1062;
input n_339;
input n_738;
input n_3679;
input n_1690;
input n_2221;
input n_2807;
input n_672;
input n_740;
input n_1283;
input n_167;
input n_2317;
input n_2838;
input n_1974;
input n_2906;
input n_1736;
input n_1018;
input n_2342;
input n_2200;
input n_2781;
input n_3283;
input n_3856;
input n_4038;
input n_69;
input n_259;
input n_2442;
input n_2735;
input n_953;
input n_1364;
input n_2390;
input n_143;
input n_1888;
input n_1224;
input n_3657;
input n_2109;
input n_1425;
input n_2634;
input n_2709;
input n_3451;
input n_625;
input n_557;
input n_2322;
input n_2746;
input n_3419;
input n_1107;
input n_2832;
input n_1688;
input n_989;
input n_242;
input n_645;
input n_1944;
input n_331;
input n_559;
input n_2233;
input n_2370;
input n_2663;
input n_267;
input n_495;
input n_2914;
input n_1988;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_3545;
input n_1718;
input n_1276;
input n_1936;
input n_2149;
input n_2277;
input n_200;
input n_1428;
input n_1284;
input n_2878;
input n_1241;
input n_3890;
input n_3830;
input n_821;
input n_561;
input n_770;
input n_3252;
input n_1514;
input n_2539;
input n_1528;
input n_507;
input n_486;
input n_901;
input n_2782;
input n_3879;
input n_569;
input n_2078;
input n_3315;
input n_3929;
input n_1145;
input n_3523;
input n_971;
input n_3144;
input n_2359;
input n_3999;
input n_2201;
input n_787;
input n_4012;
input n_1650;
input n_31;
input n_1519;
input n_1195;
input n_2049;
input n_1522;
input n_518;
input n_1207;
input n_222;
input n_3606;
input n_786;
input n_1404;
input n_3347;
input n_3420;
input n_3859;
input n_868;
input n_3474;
input n_2232;
input n_1847;
input n_2458;
input n_2779;
input n_3627;
input n_3596;
input n_3150;
input n_2950;
input n_1542;
input n_3552;
input n_1314;
input n_3756;
input n_3639;
input n_3254;
input n_1512;
input n_2227;
input n_2301;
input n_1539;
input n_2859;
input n_3121;
input n_2847;
input n_884;
input n_3412;
input n_4077;
input n_1851;
input n_2162;
input n_3209;
input n_3324;
input n_3015;
input n_1415;
input n_3870;
input n_1034;
input n_1652;
input n_2192;
input n_1676;
input n_3749;
input n_1085;
input n_277;
input n_2988;
input n_1636;
input n_3482;
input n_432;
input n_293;
input n_823;
input n_1900;
input n_620;
input n_3948;
input n_93;
input n_1074;
input n_3230;
input n_859;
input n_3793;
input n_1765;
input n_4031;
input n_108;
input n_1889;
input n_587;
input n_1977;
input n_693;
input n_863;
input n_2650;
input n_303;
input n_1254;
input n_3960;
input n_929;
input n_3207;
input n_3641;
input n_2433;
input n_206;
input n_352;
input n_899;
input n_1703;
input n_2332;
input n_2391;
input n_3828;
input n_3975;
input n_3073;
input n_611;
input n_1295;
input n_2060;
input n_1850;
input n_238;
input n_365;
input n_2004;
input n_3183;
input n_3571;
input n_1013;
input n_3883;
input n_4032;
input n_4018;
input n_1495;
input n_3607;
input n_1637;
input n_3297;
input n_2571;
input n_136;
input n_334;
input n_2427;
input n_192;
input n_3325;
input n_3613;
input n_2885;
input n_661;
input n_2098;
input n_2616;
input n_1751;
input n_2874;
input n_3003;
input n_4117;
input n_300;
input n_533;
input n_3049;
input n_3136;
input n_2867;
input n_3634;
input n_1917;
input n_2456;
input n_2769;
input n_104;
input n_1924;
input n_438;
input n_1560;
input n_1654;
input n_2341;
input n_2899;
input n_1548;
input n_3066;
input n_16;
input n_1811;
input n_2045;
input n_3274;
input n_3877;
input n_440;
input n_3913;
input n_3817;
input n_3013;
input n_3612;
input n_273;
input n_2575;
input n_2722;
input n_1396;
input n_3728;
input n_1230;
input n_612;
input n_333;
input n_1840;
input n_2739;
input n_3739;
input n_376;
input n_3962;
input n_512;
input n_1597;
input n_4082;
input n_2942;
input n_1771;
input n_2902;
input n_1544;
input n_579;
input n_3271;
input n_844;
input n_1012;
input n_1267;
input n_2061;
input n_2685;
input n_3164;
input n_2094;
input n_3854;
input n_3861;
input n_2512;
input n_1354;
input n_1790;
input n_149;
input n_1213;
input n_2382;
input n_2956;
input n_237;
input n_2043;
input n_780;
input n_2349;
input n_1918;
input n_3652;
input n_3449;
input n_2788;
input n_4119;
input n_1021;
input n_1443;
input n_4000;
input n_3089;
input n_491;
input n_2595;
input n_1465;
input n_2686;
input n_3084;
input n_1949;
input n_1595;
input n_1142;
input n_1140;
input n_705;
input n_3458;
input n_570;
input n_260;
input n_2727;
input n_942;
input n_3580;
input n_1437;
input n_3860;
input n_3511;
input n_7;
input n_2077;
input n_1378;
input n_461;
input n_1121;
input n_1416;
input n_2909;
input n_209;
input n_490;
input n_3554;
input n_1461;
input n_17;
input n_2717;
input n_3012;
input n_1391;
input n_2981;
input n_1947;
input n_225;
input n_1599;
input n_1876;
input n_1006;
input n_1830;
input n_3850;
input n_575;
input n_546;
input n_3472;
input n_503;
input n_2527;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_3126;
input n_3754;
input n_2759;
input n_1245;
input n_2743;
input n_1669;
input n_2969;
input n_3429;
input n_1675;
input n_2466;
input n_676;
input n_3758;
input n_42;
input n_2038;
input n_2263;
input n_3518;
input n_3958;
input n_2800;
input n_2568;
input n_2116;
input n_2271;
input n_2145;
input n_2326;
input n_1838;
input n_3485;
input n_1594;
input n_680;
input n_1935;
input n_2806;
input n_287;
input n_3191;
input n_1716;
input n_4108;
input n_302;
input n_3777;
input n_4109;
input n_1872;
input n_380;
input n_3562;
input n_1585;
input n_2281;
input n_1432;
input n_94;
input n_2245;
input n_4;
input n_3359;
input n_3767;
input n_3841;
input n_3119;
input n_249;
input n_1108;
input n_3588;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_1590;
input n_1351;
input n_3234;
input n_3280;
input n_3413;
input n_3692;
input n_3900;
input n_2216;
input n_4115;
input n_1274;
input n_3539;
input n_257;
input n_2426;
input n_652;
input n_1819;
input n_475;
input n_135;
input n_3095;
input n_947;
input n_2134;
input n_3862;
input n_930;
input n_1260;
input n_3698;
input n_3716;
input n_1179;
input n_468;
input n_3284;
input n_3909;
input n_102;
input n_2703;
input n_182;
input n_696;
input n_1442;
input n_2926;
input n_482;
input n_2620;
input n_798;
input n_577;
input n_1833;
input n_407;
input n_1691;
input n_27;
input n_916;
input n_1386;
input n_2810;
input n_3391;
input n_3506;
input n_912;
input n_1884;
input n_460;
input n_1555;
input n_1842;
input n_2499;
input n_2549;
input n_3678;
input n_366;
input n_762;
input n_1253;
input n_1468;
input n_1661;
input n_2791;
input n_555;
input n_2683;
input n_3212;
input n_804;
input n_1656;
input n_1382;
input n_3093;
input n_3529;
input n_2970;
input n_3159;
input n_966;
input n_992;
input n_955;
input n_3549;
input n_3885;
input n_3914;
input n_3624;
input n_1182;
input n_794;
input n_2855;
input n_78;
input n_2166;
input n_2848;
input n_1692;
input n_3192;
input n_2611;
input n_1562;
input n_514;
input n_2748;
input n_418;
input n_2185;
input n_3306;
input n_3250;
input n_3029;
input n_2398;
input n_3538;
input n_3915;
input n_1376;
input n_3839;
input n_513;
input n_288;
input n_179;
input n_1292;
input n_1178;
input n_1972;
input n_2015;
input n_2925;
input n_1435;
input n_3407;
input n_3717;
input n_1750;
input n_1026;
input n_1506;
input n_3460;
input n_3544;
input n_1610;
input n_3875;
input n_4029;
input n_2202;
input n_2072;
input n_3852;
input n_306;
input n_2952;
input n_3530;
input n_2415;
input n_2693;
input n_2877;
input n_92;
input n_4099;
input n_3120;
input n_203;
input n_2922;
input n_436;
input n_3000;
input n_150;
input n_2871;
input n_2930;
input n_3193;
input n_3240;
input n_324;
input n_2745;
input n_2087;
input n_669;
input n_931;
input n_1491;
input n_2628;
input n_3219;
input n_3362;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_3937;
input n_2161;
input n_1418;
input n_746;
input n_1357;
input n_292;
input n_1079;
input n_1787;
input n_2462;
input n_3510;
input n_1389;
input n_3393;
input n_3172;
input n_2155;
input n_2659;
input n_4033;
input n_615;
input n_3747;
input n_1139;
input n_2836;
input n_3688;
input n_76;
input n_2439;
input n_2864;
input n_517;
input n_1312;
input n_1717;
input n_3604;
input n_4045;
input n_0;
input n_1812;
input n_3651;
input n_824;
input n_428;
input n_159;
input n_2172;
input n_2601;
input n_3614;
input n_3871;
input n_892;
input n_1880;
input n_959;
input n_30;
input n_2365;
input n_2257;
input n_3757;
input n_1399;
input n_1101;
input n_1567;
input n_1343;
input n_563;
input n_2219;
input n_3116;
input n_1855;
input n_3784;
input n_2100;
input n_2333;
input n_3176;
input n_144;
input n_3629;
input n_3666;
input n_3372;
input n_3891;
input n_990;
input n_1623;
input n_3559;
input n_1903;
input n_3792;
input n_867;
input n_2147;
input n_3479;
input n_4020;
input n_2435;
input n_1226;
input n_2224;
input n_944;
input n_749;
input n_1932;
input n_1780;
input n_2825;
input n_2888;
input n_1970;
input n_3998;
input n_3724;
input n_1920;
input n_2083;
input n_815;
input n_542;
input n_3287;
input n_2167;
input n_2293;
input n_2753;
input n_1340;
input n_470;
input n_2668;
input n_1240;
input n_2921;
input n_3046;
input n_1087;
input n_4055;
input n_3980;
input n_2701;
input n_2400;
input n_3021;
input n_632;
input n_3257;
input n_477;
input n_650;
input n_3741;
input n_2388;
input n_425;
input n_3730;
input n_2273;
input n_2712;
input n_1433;
input n_3805;
input n_1911;
input n_3979;
input n_3912;
input n_2567;
input n_3950;
input n_3496;
input n_3493;
input n_2557;
input n_2695;
input n_2898;
input n_1825;
input n_1908;
input n_1155;
input n_2598;
input n_1071;
input n_2755;
input n_3700;
input n_3727;
input n_712;
input n_976;
input n_3567;
input n_909;
input n_4003;
input n_1392;
input n_767;
input n_1832;
input n_2795;
input n_2682;
input n_1841;
input n_1680;
input n_2066;
input n_2302;
input n_2762;
input n_964;
input n_1627;
input n_2220;
input n_2954;
input n_382;
input n_3014;
input n_489;
input n_2294;
input n_80;
input n_2274;
input n_3342;
input n_2895;
input n_2903;
input n_251;
input n_974;
input n_506;
input n_3814;
input n_3812;
input n_3127;
input n_3796;
input n_1731;
input n_799;
input n_3884;
input n_1147;
input n_2829;
input n_2378;
input n_3625;
input n_397;
input n_2467;
input n_3375;
input n_2768;
input n_471;
input n_351;
input n_965;
input n_1914;
input n_155;
input n_3760;
input n_2253;
input n_934;
input n_2213;
input n_3515;
input n_1447;
input n_2363;
input n_1220;
input n_356;
input n_2019;
input n_698;
input n_4056;
input n_2728;
input n_2130;
input n_1674;
input n_2021;
input n_2025;
input n_3010;
input n_2160;
input n_1992;
input n_124;
input n_3744;
input n_4015;
input n_2924;
input n_307;
input n_1209;
input n_4022;
input n_1020;
input n_1563;
input n_3673;
input n_3052;
input n_646;
input n_2507;
input n_3438;
input n_2142;
input n_1633;
input n_34;
input n_404;
input n_2625;
input n_2896;
input n_172;
input n_1913;
input n_2069;
input n_2495;
input n_3187;
input n_1058;
input n_2328;
input n_4043;
input n_347;
input n_2434;
input n_1042;
input n_3170;
input n_183;
input n_1234;
input n_2311;
input n_479;
input n_3936;
input n_1578;
input n_2261;
input n_1455;
input n_3147;
input n_2287;
input n_299;
input n_836;
input n_2223;
input n_3082;
input n_1279;
input n_3415;
input n_3661;
input n_2473;
input n_3320;
input n_2144;
input n_2511;
input n_3464;
input n_564;
input n_3414;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_2649;
input n_3981;
input n_1247;
input n_760;
input n_522;
input n_2438;
input n_1568;
input n_2919;
input n_20;
input n_3210;
input n_1483;
input n_3108;
input n_1363;
input n_2681;
input n_3867;
input n_3397;
input n_367;
input n_1111;
input n_970;
input n_1689;
input n_2535;
input n_3467;
input n_713;
input n_1255;
input n_2632;
input n_1646;
input n_598;
input n_3031;
input n_345;
input n_2262;
input n_3179;
input n_2565;
input n_3889;
input n_1237;
input n_3262;
input n_927;
input n_261;
input n_1095;
input n_2980;
input n_1728;
input n_2335;
input n_3078;
input n_3699;
input n_3971;
input n_370;
input n_706;
input n_2120;
input n_286;
input n_3239;
input n_2631;
input n_3215;
input n_3311;
input n_3869;
input n_3516;
input n_1401;
input n_1419;
input n_3138;
input n_1531;
input n_776;
input n_424;
input n_2860;
input n_3816;
input n_2041;
input n_2113;
input n_1933;
input n_3528;
input n_1651;
input n_3087;
input n_85;
input n_130;
input n_2697;
input n_1387;
input n_466;
input n_1263;
input n_346;
input n_1817;
input n_3711;
input n_2404;
input n_2168;
input n_2757;
input n_3704;
input n_348;
input n_552;
input n_2312;
input n_670;
input n_2677;
input n_1826;
input n_3171;
input n_379;
input n_138;
input n_162;
input n_264;
input n_3577;
input n_2834;
input n_4051;
input n_2483;
input n_4074;
input n_3994;
input n_441;
input n_1951;
input n_3185;
input n_2490;
input n_1032;
input n_1217;
input n_2558;
input n_1496;
input n_2996;
input n_637;
input n_1592;
input n_2812;
input n_3660;
input n_73;
input n_327;
input n_2662;
input n_1259;
input n_3300;
input n_2801;
input n_1177;
input n_3104;
input n_3074;
input n_2655;
input n_1231;
input n_3917;
input n_4122;
input n_3246;
input n_2132;
input n_3299;
input n_980;
input n_1618;
input n_3774;
input n_1869;
input n_3589;
input n_3623;
input n_1743;
input n_905;
input n_2718;
input n_207;
input n_720;
input n_926;
input n_41;
input n_1943;
input n_2687;
input n_2296;
input n_3876;
input n_3615;
input n_3267;
input n_194;
input n_1802;
input n_2178;
input n_3946;
input n_2112;
input n_2765;
input n_1163;
input n_2640;
input n_3054;
input n_2811;
input n_3019;
input n_186;
input n_1795;
input n_3200;
input n_1384;
input n_3642;
input n_2237;
input n_145;
input n_2146;
input n_2983;
input n_1868;
input n_3276;
input n_59;
input n_3601;
input n_4089;
input n_1501;
input n_2241;
input n_2373;
input n_1173;
input n_3498;
input n_3513;
input n_3682;
input n_2350;
input n_3881;
input n_1068;
input n_1198;
input n_4096;
input n_2531;
input n_1570;
input n_2099;
input n_3759;
input n_3377;
input n_487;
input n_1518;
input n_3323;
input n_1456;
input n_4007;
input n_90;
input n_1879;
input n_1886;
input n_1648;
input n_2187;
input n_3961;
input n_1413;
input n_2617;
input n_2481;
input n_3863;
input n_2129;
input n_855;
input n_2327;
input n_158;
input n_3882;
input n_3916;
input n_808;
input n_1365;
input n_2476;
input n_553;
input n_2814;
input n_2059;
input n_3675;
input n_3968;
input n_2437;
input n_2636;
input n_1439;
input n_814;
input n_578;
input n_3466;
input n_2074;
input n_1665;
input n_1287;
input n_2841;
input n_405;
input n_1611;
input n_2122;
input n_120;
input n_3572;
input n_2975;
input n_3332;
input n_2399;
input n_320;
input n_1414;
input n_1134;
input n_2067;
input n_3374;
input n_3471;
input n_4075;
input n_1484;
input n_1901;
input n_647;
input n_2055;
input n_2998;
input n_3465;
input n_2027;
input n_2932;
input n_1423;
input n_2117;
input n_481;
input n_600;
input n_1053;
input n_1609;
input n_3118;
input n_4072;
input n_2822;
input n_1939;
input n_2308;
input n_2242;
input n_1906;
input n_529;
input n_1899;
input n_3039;
input n_2195;
input n_3922;
input n_502;
input n_2194;
input n_2937;
input n_218;
input n_3508;
input n_1467;
input n_4039;
input n_247;
input n_1828;
input n_2159;
input n_1798;
input n_3057;
input n_1304;
input n_1608;
input n_3831;
input n_1744;
input n_3335;
input n_3007;
input n_2267;
input n_1105;
input n_547;
input n_3599;
input n_3618;
input n_439;
input n_604;
input n_677;
input n_3705;
input n_3022;
input n_478;
input n_703;
input n_3983;
input n_1349;
input n_1709;
input n_3318;
input n_1061;
input n_3385;
input n_2102;
input n_326;
input n_681;
input n_3477;
input n_227;
input n_3286;
input n_3734;
input n_3370;
input n_874;
input n_3773;
input n_3949;
input n_2286;
input n_3494;
input n_2023;
input n_1278;
input n_707;
input n_3974;
input n_3443;
input n_11;
input n_3401;
input n_129;
input n_126;
input n_983;
input n_3036;
input n_2783;
input n_2599;
input n_3988;
input n_3788;
input n_3939;
input n_590;
input n_699;
input n_727;
input n_301;
input n_1726;
input n_2075;
input n_3263;
input n_3542;
input n_2523;
input n_1945;
input n_3569;
input n_3835;
input n_3837;
input n_545;
input n_1015;
input n_2418;
input n_1377;
input n_1162;
input n_536;
input n_1614;
input n_2031;
input n_2496;
input n_3260;
input n_3349;
input n_3761;
input n_3819;
input n_3996;
input n_2118;
input n_325;
input n_1740;
input n_3222;
input n_1602;
input n_688;
input n_3139;
input n_636;
input n_2853;
input n_427;
input n_3350;
input n_3801;
input n_1098;
input n_3009;
input n_1490;
input n_2338;
input n_442;
input n_777;
input n_3764;
input n_1553;
input n_1080;
input n_920;
input n_1760;
input n_1086;
input n_1092;
input n_3025;
input n_3636;
input n_3051;
input n_3205;
input n_2225;
input n_986;
input n_1104;
input n_1963;
input n_2802;
input n_3653;
input n_3951;
input n_3868;
input n_3035;
input n_3823;
input n_729;
input n_887;
input n_3403;
input n_2057;
input n_2218;
input n_1122;
input n_1205;
input n_1408;
input n_2593;
input n_163;
input n_1693;
input n_2125;
input n_2716;
input n_1132;
input n_390;
input n_1156;
input n_2741;
input n_501;
input n_2184;
input n_2714;
input n_314;
input n_1823;
input n_2944;
input n_2861;
input n_2780;
input n_3023;
input n_1120;
input n_3439;
input n_3942;
input n_1202;
input n_4084;
input n_627;
input n_2254;
input n_3130;
input n_3290;
input n_1188;
input n_1498;
input n_1371;
input n_2033;
input n_2618;
input n_4121;
input n_3602;
input n_233;
input n_957;
input n_388;
input n_1402;
input n_1242;
input n_3957;
input n_2754;
input n_2707;
input n_2774;
input n_3418;
input n_2849;
input n_1607;
input n_1489;
input n_2799;
input n_1218;
input n_2756;
input n_3611;
input n_3781;
input n_2217;
input n_221;
input n_321;
input n_86;
input n_2226;
input n_3959;
input n_3984;
input n_1586;
input n_861;
input n_3338;
input n_2962;
input n_1543;
input n_1431;
input n_877;
input n_3995;
input n_1119;
input n_3713;
input n_1863;
input n_1763;
input n_1666;
input n_3908;
input n_1500;
input n_616;
input n_2214;
input n_1055;
input n_1395;
input n_3892;
input n_1346;
input n_2763;
input n_3156;
input n_2256;
input n_1189;
input n_3337;
input n_1089;
input n_3750;
input n_3424;
input n_281;
input n_3326;
input n_3356;
input n_1859;
input n_2660;
input n_3426;
input n_262;
input n_1502;
input n_3044;
input n_1523;
input n_2190;
input n_3492;
input n_3501;
input n_1478;
input n_2732;
input n_1883;
input n_3737;
input n_2516;
input n_3931;
input n_4094;
input n_2776;
input n_2555;
input n_3216;
input n_3224;
input n_3568;
input n_1969;
input n_2708;
input n_735;
input n_297;
input n_3070;
input n_1005;
input n_3275;
input n_527;
input n_2379;
input n_46;
input n_3579;
input n_3245;
input n_84;
input n_1294;
input n_2661;
input n_1667;
input n_845;
input n_888;
input n_2894;
input n_2300;
input n_2949;
input n_3896;
input n_4049;
input n_4067;
input n_1649;
input n_2452;
input n_1677;
input n_2470;
input n_1927;
input n_1297;
input n_2827;
input n_178;
input n_3214;
input n_551;
input n_3551;
input n_417;
input n_1708;
input n_70;
input n_343;
input n_3085;
input n_3373;
input n_1222;
input n_2284;
input n_3005;
input n_3710;
input n_1844;
input n_2283;
input n_582;
input n_2526;
input n_1957;
input n_3364;
input n_1953;
input n_2643;
input n_755;
input n_1097;
input n_3803;
input n_3766;
input n_3985;
input n_1219;
input n_1711;
input n_710;
input n_1919;
input n_2994;
input n_534;
input n_1791;
input n_2508;
input n_3186;
input n_2124;
input n_1894;
input n_1460;
input n_1239;
input n_2594;
input n_3826;
input n_278;
input n_2266;
input n_3944;
input n_3417;
input n_2449;
input n_560;
input n_890;
input n_842;
input n_148;
input n_3626;
input n_1898;
input n_451;
input n_745;
input n_1741;
input n_1572;
input n_1907;
input n_1793;
input n_3180;
input n_3648;
input n_3423;
input n_61;
input n_742;
input n_1081;
input n_1373;
input n_1975;
input n_1388;
input n_1266;
input n_1540;
input n_1719;
input n_2119;
input n_2742;
input n_769;
input n_3671;
input n_1797;
input n_2366;
input n_2493;
input n_13;
input n_1753;
input n_1990;
input n_1372;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_1895;
input n_2821;
input n_3491;
input n_2690;
input n_3090;
input n_3696;
input n_2474;
input n_4104;
input n_2623;
input n_3392;
input n_982;
input n_1800;
input n_915;
input n_215;
input n_3791;
input n_1075;
input n_2008;
input n_454;
input n_298;
input n_1331;
input n_1890;
input n_2904;
input n_3064;
input n_3199;
input n_4034;
input n_1529;
input n_3353;
input n_1227;
input n_3531;
input n_2127;
input n_655;
input n_2946;
input n_3166;
input n_3151;
input n_3649;
input n_3684;
input n_3333;
input n_3512;
input n_1734;
input n_1860;
input n_3065;
input n_403;
input n_3016;
input n_2785;
input n_2460;
input n_4114;
input n_2840;
input n_1007;
input n_1580;
input n_1319;
input n_3135;
input n_657;
input n_3367;
input n_3669;
input n_3956;
input n_3924;
input n_4081;
input n_837;
input n_812;
input n_2448;
input n_3997;
input n_2211;
input n_4040;
input n_2292;
input n_2480;
input n_606;
input n_951;
input n_3024;
input n_2772;
input n_3564;
input n_862;
input n_1700;
input n_2637;
input n_659;
input n_1332;
input n_3795;
input n_2306;
input n_509;
input n_1854;
input n_666;
input n_1747;
input n_2071;
input n_2424;
input n_3990;
input n_430;
input n_1206;
input n_1729;
input n_722;
input n_1508;
input n_3953;
input n_2414;
input n_2082;
input n_2893;
input n_2959;
input n_1532;
input n_3277;
input n_1171;
input n_1030;
input n_785;
input n_3161;
input n_3208;
input n_2389;
input n_4069;
input n_1309;
input n_3582;
input n_999;
input n_2280;
input n_1766;
input n_1338;
input n_2978;
input n_1342;
input n_2737;
input n_3282;
input n_456;
input n_1867;
input n_3993;
input n_852;
input n_1394;
input n_2916;
input n_2576;
input n_3459;
input n_3617;
input n_704;
input n_2958;
input n_3365;
input n_1060;
input n_1044;
input n_1714;
input n_4113;
input n_2696;
input n_3340;
input n_521;
input n_2140;
input n_873;
input n_1301;
input n_1748;
input n_2157;
input n_1966;
input n_1243;
input n_2171;
input n_2468;
input n_3977;
input n_1400;
input n_4112;
input n_342;
input n_3400;
input n_2035;
input n_2614;
input n_1466;
input n_3735;
input n_3486;
input n_1513;
input n_1527;
input n_2581;
input n_358;
input n_1783;
input n_3656;
input n_608;
input n_2494;
input n_1538;
input n_2831;
input n_2457;
input n_2128;
input n_3069;
input n_2992;
input n_1037;
input n_3650;
input n_4071;
input n_1329;
input n_317;
input n_3197;
input n_1993;
input n_1545;
input n_3586;
input n_134;
input n_2629;
input n_3369;
input n_4035;
input n_3256;
input n_1257;
input n_1480;
input n_1954;
input n_3670;
input n_1668;
input n_1878;
input n_3964;
input n_2540;
input n_3836;
input n_3302;
input n_1605;
input n_1078;
input n_3060;
input n_266;
input n_2486;
input n_1897;
input n_2984;
input n_4009;
input n_157;
input n_3646;
input n_2520;
input n_2137;
input n_1161;
input n_2489;
input n_3685;
input n_811;
input n_3097;
input n_624;
input n_3507;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_2492;
input n_3864;
input n_2939;
input n_3425;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_1449;
input n_3450;
input n_3748;
input n_2337;
input n_2265;
input n_687;
input n_2900;
input n_797;
input n_2026;
input n_2912;
input n_3524;
input n_1786;
input n_2627;
input n_4050;
input n_3173;
input n_480;
input n_1327;
input n_3732;
input n_1475;
input n_211;
input n_642;
input n_1804;
input n_2106;
input n_97;
input n_408;
input n_1406;
input n_595;
input n_1405;
input n_2684;
input n_3174;
input n_3314;
input n_2726;
input n_602;
input n_3813;
input n_2622;
input n_3447;
input n_4006;
input n_2272;
input n_3266;
input n_1757;
input n_592;
input n_3102;
input n_1499;
input n_854;
input n_1318;
input n_3452;
input n_2091;
input n_393;
input n_1632;
input n_1769;
input n_474;
input n_1929;
input n_4098;
input n_1950;
input n_2264;
input n_2691;
input n_3789;
input n_805;
input n_2032;
input n_2090;
input n_2929;
input n_3124;
input n_3811;
input n_3422;
input n_295;
input n_1658;
input n_190;
input n_2249;
input n_1072;
input n_3411;
input n_695;
input n_1526;
input n_2991;
input n_3463;
input n_1305;
input n_64;
input n_180;
input n_730;
input n_386;
input n_1596;
input n_2348;
input n_2656;
input n_1281;
input n_516;
input n_2364;
input n_1997;
input n_2574;
input n_1137;
input n_1873;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_1476;
input n_1524;
input n_1733;
input n_1856;
input n_2016;
input n_2667;
input n_2723;
input n_2725;
input n_3925;
input n_2928;
input n_943;
input n_1118;
input n_678;
input n_2905;
input n_2884;
input n_3408;
input n_651;
input n_2850;
input n_1874;
input n_1293;
input n_3167;
input n_3746;
input n_961;
input n_469;
input n_1046;
input n_1807;
input n_726;
input n_1123;
input n_3780;
input n_1657;
input n_878;
input n_2857;
input n_3694;
input n_4118;
input n_1784;
input n_3110;
input n_3857;
input n_771;
input n_3787;
input n_4025;
input n_1321;
input n_3050;
input n_3919;
input n_3157;
input n_3753;
input n_3893;
input n_752;
input n_2307;
input n_71;
input n_1488;
input n_985;
input n_421;
input n_1330;
input n_906;
input n_3702;
input n_1180;
input n_1697;
input n_2295;
input n_2730;
input n_283;
input n_4076;
input n_806;
input n_3142;
input n_1984;
input n_1350;
input n_3453;
input n_3129;
input n_1556;
input n_649;
input n_1561;
input n_2412;
input n_2720;
input n_374;
input n_3298;
input n_3107;
input n_3495;
input n_1352;
input n_3843;
input n_2405;
input n_2815;
input n_1824;
input n_643;
input n_2606;
input n_2700;
input n_1492;
input n_226;
input n_4065;
input n_2383;
input n_2764;
input n_1441;
input n_1822;
input n_682;
input n_36;
input n_1616;
input n_2633;
input n_2416;
input n_3708;
input n_819;
input n_2386;
input n_2907;
input n_1971;
input n_2945;
input n_586;
input n_1324;
input n_1429;
input n_2064;
input n_2353;
input n_2528;
input n_1778;
input n_3543;
input n_3640;
input n_1776;
input n_3448;
input n_686;
input n_605;
input n_2936;
input n_1154;
input n_584;
input n_3609;
input n_1557;
input n_1759;
input n_1829;
input n_2325;
input n_1130;
input n_1450;
input n_3718;
input n_349;
input n_756;
input n_2022;
input n_3390;
input n_1016;
input n_2298;
input n_1149;
input n_1505;
input n_2408;
input n_2698;
input n_3740;
input n_2986;
input n_2320;
input n_3017;
input n_979;
input n_2329;
input n_2570;
input n_3140;
input n_1642;
input n_2417;
input n_2789;
input n_2;
input n_3976;
input n_2525;
input n_1815;
input n_2813;
input n_897;
input n_2546;
input n_949;
input n_2454;
input n_1493;
input n_2890;
input n_2911;
input n_515;
input n_3381;
input n_807;
input n_3455;
input n_3736;
input n_891;
input n_3313;
input n_885;
input n_1659;
input n_3955;
input n_2354;
input n_3591;
input n_198;
input n_1864;
input n_2760;
input n_3907;
input n_3086;
input n_1887;
input n_3165;
input n_1208;
input n_3317;
input n_3945;
input n_3726;
input n_3336;
input n_1987;
input n_4052;
input n_3357;
input n_3388;
input n_396;
input n_2368;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_3635;
input n_2352;
input n_3541;
input n_2502;
input n_1256;
input n_87;
input n_714;
input n_3560;
input n_3345;
input n_2170;
input n_3605;
input n_790;
input n_2244;
input n_2143;
input n_2393;
input n_354;
input n_140;
input n_725;
input n_2377;
input n_1577;
input n_3566;
input n_151;
input n_3840;
input n_3421;
input n_1448;
input n_2198;
input n_28;
input n_1009;
input n_230;
input n_3548;
input n_2652;
input n_1133;
input n_3067;
input n_154;
input n_883;
input n_142;
input n_4097;
input n_4054;
input n_3809;
input n_473;
input n_1852;
input n_801;
input n_1286;
input n_2612;
input n_818;
input n_1685;
input n_779;
input n_2410;
input n_2314;
input n_2477;
input n_2279;
input n_3169;
input n_594;
input n_3236;
input n_2222;
input n_3468;
input n_1995;
input n_1877;
input n_1397;
input n_35;
input n_1052;
input n_272;
input n_1333;
input n_1306;
input n_1849;
input n_3573;
input n_2076;
input n_2133;
input n_2203;
input n_833;
input n_2943;
input n_1426;
input n_2250;
input n_3319;
input n_2497;
input n_2247;
input n_2230;
input n_879;
input n_1117;
input n_3321;
input n_38;
input n_422;
input n_1269;
input n_1303;
input n_1547;
input n_1438;
input n_1541;
input n_597;
input n_3291;
input n_3654;
input n_75;
input n_2001;
input n_1047;
input n_3783;
input n_95;
input n_2506;
input n_1472;
input n_2413;
input n_4008;
input n_1593;
input n_2610;
input n_3715;
input n_1050;
input n_2626;
input n_566;
input n_2158;
input n_2578;
input n_2607;
input n_3643;
input n_2285;
input n_3343;
input n_3184;
input n_152;
input n_3309;
input n_2892;
input n_169;
input n_106;
input n_1201;
input n_1288;
input n_173;
input n_2605;
input n_858;
input n_2796;
input n_1185;
input n_2475;
input n_2804;
input n_2173;
input n_3982;
input n_2715;
input n_3206;
input n_335;
input n_3647;
input n_1035;
input n_3475;
input n_1143;
input n_2665;
input n_344;
input n_2070;
input n_2136;
input n_426;
input n_433;
input n_3973;
input n_3134;
input n_398;
input n_2771;
input n_62;
input n_210;
input n_1090;
input n_2403;
input n_3755;
input n_2947;
input n_1367;
input n_3842;
input n_2044;
input n_166;
input n_253;
input n_928;
input n_3886;
input n_1153;
input n_271;
input n_465;
input n_3769;
input n_4078;
input n_825;
input n_1103;
input n_732;
input n_2619;
input n_1565;
input n_1192;
input n_128;
input n_224;
input n_3738;
input n_82;
input n_894;
input n_3098;
input n_1380;
input n_1624;
input n_1801;
input n_2854;
input n_3055;
input n_420;
input n_1291;
input n_562;
input n_4070;
input n_2020;
input n_748;
input n_3987;
input n_2310;
input n_510;
input n_1045;
input n_256;
input n_3341;
input n_3600;
input n_3160;
input n_1160;
input n_2968;
input n_1882;
input n_1976;
input n_1023;
input n_2711;
input n_3223;
input n_1881;
input n_2635;
input n_2999;
input n_988;
input n_3386;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_3921;
input n_282;
input n_328;
input n_368;
input n_3043;
input n_3190;
input n_1958;
input n_2747;
input n_3667;
input n_3027;
input n_4011;
input n_467;
input n_1511;
input n_2177;
input n_3695;
input n_2713;
input n_1422;
input n_3800;
input n_2766;
input n_1965;
input n_644;
input n_3462;
input n_1197;
input n_3906;
input n_3011;
input n_3395;
input n_276;
input n_2820;
input n_2613;
input n_3226;
input n_497;
input n_3733;
input n_1165;
input n_3378;
input n_2934;
input n_1641;
input n_3967;
input n_3731;
input n_168;
input n_81;
input n_538;
input n_2845;
input n_1517;
input n_2036;
input n_576;
input n_843;
input n_511;
input n_2647;
input n_455;
input n_429;
input n_588;
input n_3358;
input n_638;
input n_2003;
input n_2533;
input n_2210;
input n_3920;
input n_1307;
input n_3444;
input n_1128;
input n_3141;
input n_2053;
input n_3851;
input n_4091;
input n_1671;
input n_1417;
input n_3476;
input n_1048;
input n_2343;
input n_775;
input n_3096;
input n_667;
input n_2419;
input n_1049;
input n_3380;
input n_2330;
input n_2826;
input n_14;
input n_869;
input n_141;
input n_846;
input n_1398;
input n_1921;
input n_2777;
input n_3238;
input n_2450;
input n_2411;
input n_1356;
input n_1341;
input n_2234;
input n_2309;
input n_3189;
input n_3233;
input n_1504;
input n_1955;
input n_2110;
input n_2431;
input n_1773;
input n_3175;
input n_1440;
input n_3289;
input n_2666;
input n_3322;
input n_1370;
input n_1603;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_2401;
input n_2935;
input n_715;
input n_889;
input n_3822;
input n_3255;
input n_3818;
input n_1066;
input n_1549;
input n_2588;
input n_2863;
input n_2331;
input n_935;
input n_2886;
input n_3827;
input n_2478;
input n_685;
input n_911;
input n_4061;
input n_361;
input n_89;
input n_2658;
input n_623;
input n_3509;
input n_3587;
input n_2608;
input n_3620;
input n_2920;
input n_1712;
input n_3344;
input n_1403;
input n_1065;
input n_453;
input n_1534;
input n_1948;
input n_3006;
input n_74;
input n_2767;
input n_810;
input n_3376;
input n_19;
input n_40;
input n_1290;
input n_181;
input n_1959;
input n_3497;
input n_617;
input n_3770;
input n_2396;
input n_3243;
input n_543;
input n_3368;
input n_1362;
input n_1559;
input n_2121;
input n_3456;
input n_3865;
input n_3123;
input n_2692;
input n_236;
input n_601;
input n_683;
input n_565;
input n_3927;
input n_628;
input n_1300;
input n_1960;
input n_4102;
input n_2068;
input n_3117;
input n_3595;
input n_743;
input n_1194;
input n_2862;
input n_4060;
input n_1647;
input n_1546;
input n_3384;
input n_1420;
input n_2553;
input n_2645;
input n_3790;
input n_907;
input n_2749;
input n_1454;
input n_2592;
input n_660;
input n_464;
input n_3490;
input n_2459;
input n_962;
input n_941;
input n_3396;
input n_1210;
input n_847;
input n_747;
input n_1622;
input n_1135;
input n_2566;
input n_2751;
input n_3113;
input n_3101;
input n_918;
input n_1968;
input n_3307;
input n_107;
input n_3662;
input n_1885;
input n_639;
input n_452;
input n_673;
input n_3251;
input n_3288;
input n_4093;
input n_2842;
input n_2833;
input n_2196;
input n_1038;
input n_3603;
input n_3723;
input n_2371;
input n_1978;
input n_414;
input n_571;
input n_3880;
input n_3720;
input n_1521;
input n_1694;
input n_1940;
input n_3683;
input n_6;
input n_284;
input n_3904;
input n_3887;
input n_593;
input n_3195;
input n_3008;
input n_1695;
input n_3242;
input n_4027;
input n_2560;
input n_1164;
input n_3405;
input n_37;
input n_58;
input n_2313;
input n_609;
input n_3077;
input n_1193;
input n_3048;
input n_3339;
input n_1345;
input n_613;
input n_3037;
input n_1022;
input n_1336;
input n_1033;
input n_3478;
input n_3062;
input n_1774;
input n_409;
input n_171;
input n_2963;
input n_3532;
input n_519;
input n_384;
input n_2609;
input n_2561;
input n_1166;
input n_1056;
input n_2007;
input n_526;
input n_1994;
input n_3363;
input n_3533;
input n_3978;
input n_1767;
input n_1040;
input n_674;
input n_3131;
input n_1158;
input n_316;
input n_3168;
input n_125;
input n_1973;
input n_1444;
input n_1803;
input n_820;
input n_1749;
input n_43;
input n_872;
input n_1653;
input n_3409;
input n_4079;
input n_3522;
input n_3583;
input n_4088;
input n_254;
input n_2882;
input n_2303;
input n_2669;
input n_3540;
input n_3911;
input n_3241;
input n_3802;
input n_3899;
input n_1157;
input n_1584;
input n_234;
input n_848;
input n_1664;
input n_3481;
input n_280;
input n_629;
input n_3563;
input n_1739;
input n_161;
input n_2642;
input n_3310;
input n_1814;
input n_532;
input n_3689;
input n_2154;
input n_2441;
input n_2236;
input n_1789;
input n_763;
input n_1986;
input n_4041;
input n_2174;
input n_2688;
input n_99;
input n_540;
input n_216;
input n_692;
input n_2624;
input n_5;
input n_3442;
input n_3972;
input n_2054;
input n_1857;
input n_2315;
input n_3926;
input n_984;
input n_1687;
input n_2073;
input n_223;
input n_2150;
input n_4004;
input n_1552;
input n_750;
input n_2938;
input n_834;
input n_3630;
input n_1612;
input n_2498;
input n_800;
input n_2638;
input n_3992;
input n_2046;
input n_1816;
input n_1910;
input n_2803;
input n_1756;
input n_2887;
input n_1606;
input n_2189;
input n_395;
input n_621;
input n_2648;
input n_3305;
input n_1587;
input n_213;
input n_3810;
input n_4062;
input n_2093;
input n_2340;
input n_2018;
input n_2672;
input n_1772;
input n_67;
input n_2444;
input n_2602;
input n_3354;
input n_1014;
input n_724;
input n_2204;
input n_2931;
input n_3433;
input n_1427;
input n_1481;
input n_2040;
input n_493;
input n_1311;
input n_2977;
input n_3106;
input n_3597;
input n_3991;
input n_2199;
input n_2881;
input n_1956;
input n_1589;
input n_114;
input n_4111;
input n_2151;
input n_1100;
input n_585;
input n_875;
input n_1617;
input n_2455;
input n_827;
input n_2600;
input n_3092;
input n_3437;
input n_2231;
input n_3786;
input n_697;
input n_2828;
input n_622;
input n_1626;
input n_3436;
input n_1962;
input n_1335;
input n_1715;
input n_3806;
input n_296;
input n_3553;
input n_4044;
input n_2305;
input n_3645;
input n_880;
input n_793;
input n_2114;
input n_3329;
input n_2927;
input n_3304;
input n_3833;
input n_3574;
input n_1175;
input n_2289;
input n_132;
input n_2530;
input n_2299;
input n_3751;
input n_3402;
input n_751;
input n_1027;
input n_1070;
input n_2406;
input n_3247;
input n_1621;
input n_4110;
input n_739;
input n_1485;
input n_1028;
input n_2883;
input n_1221;
input n_530;
input n_1785;
input n_792;
input n_1262;
input n_1942;
input n_2180;
input n_3406;
input n_2951;
input n_3807;
input n_4048;
input n_580;
input n_3664;
input n_1579;
input n_494;
input n_2809;
input n_2181;
input n_3550;
input n_434;
input n_2014;
input n_975;
input n_2974;
input n_229;
input n_394;
input n_923;
input n_1645;
input n_1124;
input n_1381;
input n_2870;
input n_1494;
input n_932;
input n_1893;
input n_1183;
input n_3686;
input n_3722;
input n_1326;
input n_2889;
input n_2276;
input n_3969;
input n_1805;
input n_2282;
input n_3301;
input n_981;
input n_4068;
input n_2910;
input n_2141;
input n_1110;
input n_1758;
input n_2503;
input n_3873;
input n_2270;
input n_3470;
input n_243;
input n_3785;
input n_3294;
input n_2443;
input n_1407;
input n_185;
input n_2465;
input n_3610;
input n_1204;
input n_2865;
input n_1554;
input n_3279;
input n_994;
input n_2428;
input n_2972;
input n_2586;
input n_2989;
input n_1360;
input n_973;
input n_3178;
input n_2858;
input n_268;
input n_972;
input n_3844;
input n_3259;
input n_2251;
input n_2923;
input n_3076;
input n_164;
input n_2843;
input n_3714;
input n_184;
input n_3410;
input n_856;
input n_3100;
input n_2572;
input n_1248;
input n_1176;
input n_3721;
input n_3676;
input n_1564;
input n_2010;
input n_3677;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_1679;
input n_3292;
input n_3389;
input n_2872;
input n_2126;
input n_3701;
input n_3109;
input n_3706;
input n_1952;
input n_2425;
input n_2394;
input n_3989;
input n_1858;
input n_353;
input n_3125;
input n_1678;
input n_2589;
input n_4086;
input n_1482;
input n_1361;
input n_2356;
input n_1601;
input n_3537;
input n_1057;
input n_191;
input n_2487;
input n_1834;
input n_978;
input n_1011;
input n_1520;
input n_2534;
input n_2488;
input n_1509;
input n_828;
input n_2941;
input n_322;
input n_1411;
input n_1359;
input n_3079;
input n_3638;
input n_3269;
input n_558;
input n_3536;
input n_1721;
input n_2564;
input n_116;
input n_3558;
input n_3576;
input n_3782;
input n_39;
input n_2591;
input n_653;
input n_1445;
input n_1317;
input n_3034;
input n_2050;
input n_2197;
input n_3502;
input n_3248;
input n_783;
input n_4053;
input n_2550;
input n_556;
input n_1127;
input n_170;
input n_1536;
input n_3177;
input n_3594;
input n_1471;
input n_2385;
input n_160;
input n_3440;
input n_119;
input n_2387;
input n_1008;
input n_3963;
input n_332;
input n_3658;
input n_581;
input n_294;
input n_3091;
input n_1024;
input n_830;
input n_176;
input n_3404;
input n_2291;
input n_3346;
input n_2816;
input n_1980;
input n_2518;
input n_987;
input n_936;
input n_2510;
input n_1620;
input n_2501;
input n_2542;
input n_3227;
input n_3570;
input n_3105;
input n_1385;
input n_1525;
input n_2793;
input n_1998;
input n_2165;
input n_2675;
input n_541;
input n_499;
input n_2604;
input n_1775;
input n_788;
input n_12;
input n_908;
input n_2639;
input n_3521;
input n_3855;
input n_1036;
input n_2169;
input n_2985;
input n_2603;
input n_341;
input n_4083;
input n_1270;
input n_109;
input n_1167;
input n_1272;
input n_549;
input n_2630;
input n_591;
input n_4105;
input n_2794;
input n_969;
input n_3663;
input n_2028;
input n_919;
input n_1663;
input n_50;
input n_3114;
input n_2901;
input n_2092;
input n_3940;
input n_2175;
input n_1625;
input n_2086;
input n_3225;
input n_3622;
input n_2773;
input n_2817;
input n_1926;
input n_2402;
input n_3621;
input n_318;
input n_1458;
input n_103;
input n_244;
input n_679;
input n_1630;
input n_3473;
input n_220;
input n_3644;
input n_3047;
input n_663;
input n_1720;
input n_2409;
input n_2966;
input n_3163;
input n_3680;
input n_443;
input n_3431;
input n_2176;
input n_3565;
input n_1412;
input n_3355;
input n_3059;
input n_1738;
input n_1550;
input n_528;
input n_1358;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_3897;
input n_139;
input n_2808;
input n_2453;
input n_2344;
input n_1922;
input n_3331;
input n_1735;
input n_1788;
input n_391;
input n_940;
input n_3520;
input n_2392;
input n_1537;
input n_2138;
input n_4005;
input n_3272;
input n_3122;
input n_3040;
input n_2065;
input n_2543;
input n_2321;
input n_1077;
input n_2597;
input n_607;
input n_956;
input n_445;
input n_3360;
input n_1930;
input n_3687;
input n_765;
input n_1809;
input n_2787;
input n_4092;
input n_3585;
input n_1843;
input n_1904;
input n_122;
input n_2000;
input n_3799;
input n_3133;
input n_2805;
input n_4037;
input n_1268;
input n_3804;
input n_2676;
input n_2758;
input n_385;
input n_3211;
input n_2395;
input n_917;
input n_2868;
input n_1271;
input n_372;
input n_2096;
input n_2440;
input n_2556;
input n_2186;
input n_15;
input n_1530;
input n_2215;
input n_4057;
input n_2770;
input n_631;
input n_399;
input n_3847;
input n_1170;
input n_2724;
input n_4073;
input n_3575;
input n_2258;
input n_1261;
input n_2471;
input n_702;
input n_3633;
input n_857;
input n_898;
input n_3042;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1323;
input n_2584;
input n_2375;
input n_3278;
input n_1462;
input n_3328;
input n_4001;
input n_1937;
input n_2012;
input n_3182;
input n_2967;
input n_3608;
input n_1064;
input n_633;
input n_900;
input n_1446;
input n_1282;
input n_3004;
input n_1701;
input n_1093;
input n_1551;
input n_2039;
input n_1755;
input n_4021;
input n_1285;
input n_3379;
input n_3111;
input n_193;
input n_733;
input n_761;
input n_2212;
input n_3838;
input n_731;
input n_336;
input n_1813;
input n_315;
input n_2268;
input n_2997;
input n_3469;
input n_4059;
input n_311;
input n_1452;
input n_2835;
input n_1573;
input n_3258;
input n_2734;
input n_8;
input n_668;
input n_2569;
input n_758;
input n_4019;
input n_3691;
input n_2252;
input n_3598;
input n_2111;
input n_3743;
input n_2420;
input n_2948;
input n_3099;
input n_1996;
input n_1106;
input n_2009;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_2897;
input n_1322;
input n_3273;
input n_3829;
input n_2583;
input n_2918;
input n_2987;
input n_1473;
input n_835;
input n_3155;
input n_446;
input n_1076;
input n_2024;
input n_1348;
input n_2651;
input n_753;
input n_2445;
input n_2733;
input n_1770;
input n_701;
input n_1003;
input n_2469;
input n_1125;
input n_2103;
input n_4024;
input n_2358;
input n_3316;
input n_4023;
input n_1710;
input n_1865;
input n_2522;
input n_2641;
input n_3632;
input n_2463;
input n_3546;
input n_309;
input n_1344;
input n_115;
input n_2355;
input n_1390;
input n_2580;
input n_2699;
input n_401;
input n_485;
input n_1792;
input n_4064;
input n_504;
input n_3351;
input n_2062;
input n_483;
input n_435;
input n_3068;
input n_1141;
input n_3457;
input n_1629;
input n_3901;
input n_291;
input n_1640;
input n_822;
input n_1094;
input n_2973;
input n_840;
input n_1459;
input n_2153;
input n_2324;
input n_1510;
input n_3454;
input n_3002;
input n_2710;
input n_2505;
input n_2139;
input n_1099;
input n_839;
input n_79;
input n_1754;
input n_3;
input n_3146;
input n_3394;
input n_3038;
input n_759;
input n_567;
input n_2397;
input n_91;
input n_2521;
input n_240;
input n_369;
input n_1727;
input n_2740;
input n_2235;
input n_44;
input n_1991;
input n_1575;
input n_3693;
input n_3878;
input n_2721;
input n_1848;
input n_1892;
input n_1172;
input n_3132;
input n_2615;
input n_614;
input n_3776;
input n_4066;
input n_2775;
input n_3903;
input n_1212;
input n_3581;
input n_3778;
input n_831;
input n_3681;
input n_3933;
input n_3970;
input n_778;
input n_48;
input n_1619;
input n_2351;
input n_3303;
input n_188;
input n_2260;
input n_323;
input n_550;
input n_1315;
input n_1660;
input n_4080;
input n_1902;
input n_997;
input n_635;
input n_2206;
input n_2784;
input n_3898;
input n_2541;
input n_694;
input n_1643;
input n_1320;
input n_3188;
input n_3001;
input n_3232;
input n_1113;
input n_3218;
input n_2347;
input n_248;
input n_3768;
input n_1152;
input n_2657;
input n_2990;
input n_2447;
input n_2034;
input n_1845;
input n_2538;
input n_3932;
input n_1934;
input n_2101;
input n_2577;
input n_921;
input n_2362;
input n_1615;
input n_1236;
input n_4100;
input n_228;
input n_2104;
input n_1265;
input n_1576;
input n_2105;
input n_1470;
input n_671;
input n_1533;
input n_1806;
input n_2372;
input n_2552;
input n_3445;
input n_4087;
input n_1;
input n_1409;
input n_1148;
input n_1588;
input n_1684;
input n_1673;
input n_2422;
input n_2704;
input n_1334;
input n_654;
input n_2290;
input n_2933;
input n_3729;
input n_3253;
input n_2856;
input n_3235;
input n_3387;
input n_2088;
input n_3265;
input n_3952;
input n_1275;
input n_3103;
input n_488;
input n_3018;
input n_904;
input n_505;
input n_88;
input n_2005;
input n_3584;
input n_2048;
input n_1696;
input n_3446;
input n_498;
input n_3028;
input n_1875;
input n_1059;
input n_3148;
input n_3775;
input n_684;
input n_2429;
input n_2108;
input n_2736;
input n_3966;
input n_3285;
input n_3824;
input n_3825;
input n_1039;
input n_2246;
input n_3616;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_2339;
input n_3846;
input n_392;
input n_1628;
input n_1289;
input n_1831;
input n_2532;
input n_2191;
input n_2971;
input n_3874;
input n_1497;
input n_1866;
input n_2472;
input n_2664;
input n_2705;
input n_2056;
input n_2852;
input n_459;
input n_1136;
input n_2515;
input n_3845;
input n_1782;
input n_458;
input n_1190;
input n_1600;
input n_1144;
input n_3203;
input n_383;
input n_838;
input n_1558;
input n_4107;
input n_1941;
input n_3628;
input n_1316;
input n_175;
input n_2519;
input n_3637;
input n_950;
input n_1017;
input n_711;
input n_3941;
input n_734;
input n_1915;
input n_2360;
input n_723;
input n_1393;
input n_2240;
input n_658;
input n_630;
input n_1369;
input n_53;
input n_362;
input n_2846;
input n_310;
input n_3371;
input n_1781;
input n_709;
input n_2917;
input n_3137;
input n_2544;
input n_24;
input n_809;
input n_3143;
input n_3194;
input n_3690;
input n_2085;
input n_2432;
input n_3229;
input n_3032;
input n_3872;
input n_1686;
input n_1964;
input n_3659;
input n_3928;
input n_235;
input n_881;
input n_1019;
input n_1477;
input n_1777;
input n_2188;
input n_1982;
input n_2097;
input n_662;
input n_641;
input n_3366;
input n_3461;
input n_2430;
input n_2504;
input n_910;
input n_290;
input n_741;
input n_939;
input n_1410;
input n_2297;
input n_3094;
input n_3441;
input n_371;
input n_199;
input n_3020;
input n_4002;
input n_217;
input n_2964;
input n_1114;
input n_1325;
input n_1742;
input n_708;
input n_308;
input n_1223;
input n_3815;
input n_2545;
input n_201;
input n_1768;
input n_2513;
input n_2193;
input n_2369;
input n_572;
input n_1199;
input n_2957;
input n_865;
input n_10;
input n_1273;
input n_1983;
input n_2982;
input n_1041;
input n_2451;
input n_3312;
input n_2115;
input n_2913;
input n_993;
input n_1862;
input n_948;
input n_2017;
input n_3752;
input n_3672;
input n_922;
input n_1004;
input n_1810;
input n_3061;
input n_448;
input n_2587;
input n_3504;
input n_1347;
input n_2839;
input n_3237;
input n_860;
input n_3555;
input n_3820;
input n_3072;
input n_1043;
input n_2961;
input n_255;
input n_2869;
input n_3534;
input n_450;
input n_4036;
input n_1923;
input n_3848;
input n_3655;
input n_2955;
input n_2670;
input n_3631;
input n_1764;
input n_2674;
input n_3556;
input n_896;
input n_1737;
input n_1479;
input n_1613;
input n_3026;
input n_2644;
input n_902;
input n_1031;
input n_2979;
input n_1723;
input n_3674;
input n_1638;
input n_853;
input n_3071;
input n_3918;
input n_716;
input n_4010;
input n_1571;
input n_1698;
input n_3902;
input n_4101;
input n_196;
input n_3866;
input n_1337;
input n_3763;
input n_774;
input n_1946;
input n_2148;
input n_933;
input n_3244;
input n_3499;
input n_1779;
input n_2562;
input n_596;
input n_954;
input n_2051;
input n_3112;
input n_1168;
input n_1821;
input n_4095;
input n_219;
input n_1310;
input n_3296;
input n_3196;
input n_3762;
input n_3794;
input n_231;
input n_3910;
input n_3947;
input n_656;
input n_492;
input n_574;
input n_3593;
input n_2673;
input n_252;
input n_664;
input n_1591;
input n_2585;
input n_2995;
input n_3293;
input n_3361;
input n_1229;
input n_1683;
input n_2582;
input n_3228;
input n_3327;
input n_2548;
input n_68;
input n_3488;
input n_1896;
input n_2164;
input n_1732;
input n_415;
input n_2381;
input n_2744;
input n_1967;
input n_2384;
input n_2678;
input n_2179;
input n_63;
input n_1280;
input n_544;
input n_1516;
input n_1186;
input n_1705;
input n_599;
input n_768;
input n_3707;
input n_1091;
input n_2052;
input n_2485;
input n_3779;
input n_3895;
input n_3149;
input n_537;
input n_1063;
input n_3934;
input n_25;
input n_991;
input n_2183;
input n_2205;
input n_83;
input n_2275;
input n_389;
input n_2563;
input n_1724;
input n_3088;
input n_1670;
input n_1707;
input n_1799;
input n_2080;
input n_3590;
input n_2058;
input n_3231;
input n_1126;
input n_3834;
input n_2761;
input n_2357;
input n_2029;
input n_195;
input n_1846;
input n_1912;
input n_3923;
input n_938;
input n_1891;
input n_1328;
input n_895;
input n_110;
input n_304;
input n_2875;
input n_1639;
input n_583;
input n_3519;
input n_2209;
input n_2421;
input n_1302;
input n_3295;
input n_1000;
input n_313;
input n_626;
input n_4042;
input n_378;
input n_1581;
input n_3849;
input n_1928;
input n_98;
input n_946;
input n_757;
input n_2047;
input n_3058;
input n_375;
input n_113;
input n_1655;
input n_1818;
input n_33;
input n_1146;
input n_2792;
input n_3398;
input n_3709;
input n_1634;
input n_2596;
input n_1203;
input n_998;
input n_1699;
input n_1598;
input n_3557;
input n_3592;
input n_3725;
input n_3986;
input n_2269;
input n_472;
input n_937;
input n_1474;
input n_2081;
input n_4026;
input n_2536;
input n_2524;
input n_265;
input n_1583;
input n_1604;
input n_208;
input n_1631;
input n_1702;
input n_3399;
input n_3894;
input n_156;
input n_174;
input n_275;
input n_100;
input n_3202;
input n_1794;
input n_1375;
input n_3053;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_1368;
input n_963;
input n_3772;
input n_1264;
input n_51;
input n_1082;
input n_1725;
input n_496;
input n_2891;
input n_2318;
input n_1827;
input n_3128;
input n_4120;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1752;
input n_1313;
input n_1001;
input n_1722;
input n_2361;
input n_1115;
input n_2229;
input n_2819;
input n_2880;
input n_3030;
input n_3075;
input n_3505;
input n_1339;
input n_1002;
input n_1644;
input n_105;
input n_1051;
input n_3547;
input n_4014;
input n_3771;
input n_2551;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_2255;
input n_1129;
input n_1252;
input n_2239;
input n_3045;
input n_250;
input n_1464;
input n_1296;
input n_3158;
input n_773;
input n_2798;
input n_3221;
input n_2316;
input n_165;
input n_3217;
input n_2464;
input n_3697;
input n_1010;
input n_2830;
input n_882;
input n_2706;
input n_2304;
input n_1249;
input n_101;
input n_803;
input n_1871;
input n_2514;
input n_329;
input n_718;
input n_3821;
input n_1434;
input n_340;
input n_1905;
input n_1569;
input n_3201;
input n_3334;
input n_4016;
input n_2573;
input n_2940;
input n_3503;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_3427;
input n_2336;
input n_523;
input n_1662;
input n_3162;
input n_457;
input n_1299;
input n_1870;
input n_3249;
input n_3430;
input n_3483;
input n_4046;
input n_177;
input n_2063;
input n_1925;
input n_782;
input n_364;
input n_258;
input n_2915;
input n_3489;
input n_3083;
input n_431;
input n_2654;
input n_3935;
input n_2491;
input n_1861;
input n_2079;
input n_1228;
input n_2319;
input n_2152;
input n_3213;
input n_2517;
input n_1931;
input n_4047;
input n_1244;
input n_3484;
input n_1796;
input n_411;
input n_484;
input n_2259;
input n_849;
input n_2095;
input n_2719;
input n_22;
input n_2965;
input n_2738;
input n_1820;
input n_2590;
input n_2876;
input n_2797;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_1989;
input n_3041;
input n_447;
input n_1421;
input n_2208;
input n_2423;
input n_2689;
input n_4063;
input n_2778;
input n_1762;
input n_1233;
input n_3798;
input n_3080;
input n_1808;
input n_1574;
input n_1672;
input n_2228;
input n_1635;
input n_3033;
input n_1704;
input n_3832;
input n_893;
input n_3525;
input n_3308;
input n_3712;
input n_1582;
input n_841;
input n_2479;
input n_3204;
input n_886;
input n_1069;
input n_1981;
input n_2824;
input n_2037;
input n_2953;
input n_359;
input n_3428;
input n_1308;
input n_573;
input n_796;
input n_2851;
input n_2823;
input n_4017;
input n_127;
input n_531;
input n_2345;
input n_1730;
input n_1374;
input n_1451;
input n_2089;
input n_1487;
input n_675;

output n_16275;

wire n_4474;
wire n_9872;
wire n_14741;
wire n_16050;
wire n_9604;
wire n_10943;
wire n_10453;
wire n_12407;
wire n_7329;
wire n_15048;
wire n_12343;
wire n_13909;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_14469;
wire n_11913;
wire n_8165;
wire n_5093;
wire n_12760;
wire n_4586;
wire n_11172;
wire n_12018;
wire n_14470;
wire n_15304;
wire n_6603;
wire n_6557;
wire n_10678;
wire n_5402;
wire n_11190;
wire n_13957;
wire n_6581;
wire n_15154;
wire n_16227;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_11458;
wire n_11999;
wire n_5717;
wire n_10649;
wire n_13176;
wire n_10794;
wire n_12945;
wire n_4283;
wire n_9297;
wire n_11627;
wire n_4403;
wire n_10557;
wire n_13125;
wire n_8139;
wire n_15369;
wire n_11453;
wire n_4962;
wire n_14456;
wire n_7832;
wire n_16166;
wire n_8438;
wire n_12806;
wire n_12244;
wire n_11135;
wire n_11306;
wire n_15390;
wire n_15157;
wire n_4302;
wire n_14658;
wire n_12589;
wire n_5791;
wire n_7127;
wire n_13109;
wire n_4547;
wire n_14209;
wire n_13718;
wire n_5090;
wire n_8321;
wire n_5302;
wire n_15105;
wire n_10000;
wire n_12103;
wire n_7922;
wire n_7805;
wire n_9807;
wire n_7542;
wire n_12354;
wire n_11783;
wire n_7053;
wire n_16181;
wire n_11614;
wire n_9892;
wire n_5712;
wire n_14807;
wire n_11143;
wire n_6297;
wire n_4982;
wire n_10704;
wire n_14334;
wire n_11431;
wire n_11799;
wire n_8699;
wire n_9263;
wire n_9734;
wire n_8037;
wire n_5479;
wire n_8257;
wire n_4610;
wire n_6058;
wire n_11246;
wire n_10213;
wire n_11377;
wire n_13029;
wire n_9886;
wire n_15093;
wire n_5263;
wire n_10904;
wire n_15293;
wire n_5565;
wire n_9096;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_8997;
wire n_13215;
wire n_14066;
wire n_9985;
wire n_15841;
wire n_9665;
wire n_14300;
wire n_12233;
wire n_11349;
wire n_7001;
wire n_10169;
wire n_10903;
wire n_13875;
wire n_11906;
wire n_6129;
wire n_13755;
wire n_14335;
wire n_14473;
wire n_13910;
wire n_15347;
wire n_4321;
wire n_15801;
wire n_10574;
wire n_13066;
wire n_5590;
wire n_10468;
wire n_14226;
wire n_6524;
wire n_9241;
wire n_16188;
wire n_16032;
wire n_9286;
wire n_4853;
wire n_8744;
wire n_9592;
wire n_5229;
wire n_15921;
wire n_12574;
wire n_6313;
wire n_12260;
wire n_7464;
wire n_8449;
wire n_15404;
wire n_9683;
wire n_10380;
wire n_10968;
wire n_14979;
wire n_4260;
wire n_13491;
wire n_7626;
wire n_9939;
wire n_15874;
wire n_12315;
wire n_10688;
wire n_9358;
wire n_16157;
wire n_9466;
wire n_8953;
wire n_11756;
wire n_7965;
wire n_13636;
wire n_7368;
wire n_9787;
wire n_8399;
wire n_6664;
wire n_8598;
wire n_10276;
wire n_15671;
wire n_7562;
wire n_11604;
wire n_9997;
wire n_7534;
wire n_13196;
wire n_7428;
wire n_12581;
wire n_4512;
wire n_6190;
wire n_8460;
wire n_12085;
wire n_14960;
wire n_4132;
wire n_16108;
wire n_13980;
wire n_14861;
wire n_7373;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_9318;
wire n_10281;
wire n_16224;
wire n_13715;
wire n_12089;
wire n_8734;
wire n_12671;
wire n_14592;
wire n_15750;
wire n_8720;
wire n_10528;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_12993;
wire n_13120;
wire n_8114;
wire n_4824;
wire n_8422;
wire n_12728;
wire n_7467;
wire n_14572;
wire n_8126;
wire n_5340;
wire n_6797;
wire n_7392;
wire n_9714;
wire n_14405;
wire n_14598;
wire n_16147;
wire n_15441;
wire n_10399;
wire n_4741;
wire n_7526;
wire n_8664;
wire n_10131;
wire n_11721;
wire n_14378;
wire n_11736;
wire n_4143;
wire n_14430;
wire n_10634;
wire n_4273;
wire n_11444;
wire n_11891;
wire n_13058;
wire n_4136;
wire n_14094;
wire n_9809;
wire n_11492;
wire n_14636;
wire n_9613;
wire n_9354;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_12647;
wire n_9897;
wire n_9295;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_15363;
wire n_15602;
wire n_10595;
wire n_11767;
wire n_13180;
wire n_6253;
wire n_15577;
wire n_9119;
wire n_6128;
wire n_9058;
wire n_6197;
wire n_7200;
wire n_8326;
wire n_11807;
wire n_11944;
wire n_13090;
wire n_15161;
wire n_11474;
wire n_5589;
wire n_11819;
wire n_15423;
wire n_8504;
wire n_8920;
wire n_5744;
wire n_12080;
wire n_6808;
wire n_5691;
wire n_7937;
wire n_16257;
wire n_8985;
wire n_7490;
wire n_13069;
wire n_6295;
wire n_11409;
wire n_5403;
wire n_11692;
wire n_13138;
wire n_12599;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_6992;
wire n_10644;
wire n_12863;
wire n_8035;
wire n_11856;
wire n_5830;
wire n_9516;
wire n_15063;
wire n_13996;
wire n_13064;
wire n_8660;
wire n_15593;
wire n_6681;
wire n_4227;
wire n_15788;
wire n_5158;
wire n_9917;
wire n_12185;
wire n_5152;
wire n_8939;
wire n_11737;
wire n_11652;
wire n_15326;
wire n_11038;
wire n_5092;
wire n_13991;
wire n_6542;
wire n_13466;
wire n_9202;
wire n_13689;
wire n_13896;
wire n_11925;
wire n_14115;
wire n_6161;
wire n_15930;
wire n_4505;
wire n_11974;
wire n_12457;
wire n_6452;
wire n_10426;
wire n_5247;
wire n_9512;
wire n_9923;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_10070;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_12792;
wire n_7507;
wire n_13458;
wire n_8176;
wire n_9677;
wire n_7215;
wire n_7379;
wire n_7441;
wire n_5210;
wire n_15481;
wire n_5292;
wire n_8327;
wire n_12556;
wire n_8991;
wire n_7438;
wire n_11200;
wire n_8855;
wire n_4443;
wire n_9811;
wire n_13762;
wire n_9508;
wire n_13441;
wire n_13532;
wire n_5086;
wire n_6136;
wire n_14236;
wire n_11597;
wire n_5843;
wire n_7874;
wire n_11309;
wire n_14156;
wire n_15702;
wire n_8539;
wire n_13118;
wire n_8630;
wire n_9308;
wire n_14587;
wire n_15566;
wire n_8533;
wire n_13830;
wire n_11233;
wire n_7108;
wire n_11047;
wire n_9638;
wire n_15665;
wire n_11068;
wire n_13912;
wire n_15057;
wire n_15429;
wire n_13768;
wire n_4529;
wire n_11476;
wire n_8435;
wire n_7695;
wire n_10245;
wire n_6156;
wire n_11611;
wire n_13111;
wire n_8098;
wire n_4908;
wire n_11957;
wire n_8204;
wire n_5060;
wire n_13290;
wire n_12509;
wire n_12663;
wire n_9199;
wire n_12155;
wire n_15221;
wire n_13379;
wire n_15828;
wire n_7162;
wire n_4432;
wire n_11210;
wire n_9808;
wire n_7331;
wire n_10457;
wire n_5913;
wire n_8958;
wire n_13838;
wire n_4530;
wire n_11333;
wire n_11682;
wire n_9821;
wire n_5614;
wire n_13692;
wire n_16187;
wire n_5391;
wire n_5452;
wire n_10715;
wire n_11381;
wire n_7944;
wire n_11922;
wire n_5249;
wire n_13126;
wire n_14762;
wire n_12068;
wire n_10579;
wire n_7850;
wire n_5076;
wire n_10707;
wire n_5757;
wire n_15682;
wire n_9265;
wire n_6872;
wire n_15357;
wire n_15098;
wire n_12332;
wire n_12858;
wire n_6644;
wire n_11352;
wire n_9143;
wire n_5062;
wire n_12641;
wire n_4912;
wire n_12140;
wire n_9845;
wire n_4226;
wire n_10112;
wire n_14505;
wire n_10556;
wire n_14150;
wire n_4311;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_7607;
wire n_14292;
wire n_13330;
wire n_7642;
wire n_8373;
wire n_16075;
wire n_8424;
wire n_13417;
wire n_8442;
wire n_9304;
wire n_14492;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_15909;
wire n_4827;
wire n_6801;
wire n_11152;
wire n_13505;
wire n_4993;
wire n_7397;
wire n_7205;
wire n_10080;
wire n_14951;
wire n_11022;
wire n_4871;
wire n_11025;
wire n_12517;
wire n_4405;
wire n_16228;
wire n_6563;
wire n_5968;
wire n_11251;
wire n_13821;
wire n_10766;
wire n_13787;
wire n_6398;
wire n_11222;
wire n_5586;
wire n_14065;
wire n_7461;
wire n_8519;
wire n_11650;
wire n_14310;
wire n_15420;
wire n_14958;
wire n_15690;
wire n_8075;
wire n_5468;
wire n_7638;
wire n_4745;
wire n_10781;
wire n_11091;
wire n_13243;
wire n_13531;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_8642;
wire n_15565;
wire n_11713;
wire n_8648;
wire n_10217;
wire n_7224;
wire n_6966;
wire n_9791;
wire n_5056;
wire n_9449;
wire n_9934;
wire n_9149;
wire n_9686;
wire n_13063;
wire n_13186;
wire n_14639;
wire n_15101;
wire n_13463;
wire n_15748;
wire n_7259;
wire n_7838;
wire n_8556;
wire n_5984;
wire n_12961;
wire n_14039;
wire n_11398;
wire n_9844;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_12389;
wire n_7307;
wire n_6776;
wire n_15472;
wire n_11208;
wire n_9458;
wire n_4951;
wire n_4959;
wire n_8585;
wire n_7840;
wire n_15994;
wire n_9717;
wire n_11858;
wire n_12595;
wire n_11487;
wire n_14194;
wire n_8455;
wire n_8444;
wire n_13237;
wire n_9128;
wire n_14788;
wire n_10638;
wire n_14559;
wire n_14255;
wire n_11745;
wire n_10239;
wire n_12368;
wire n_13353;
wire n_6624;
wire n_7888;
wire n_8560;
wire n_15360;
wire n_12816;
wire n_14730;
wire n_11525;
wire n_6710;
wire n_6883;
wire n_9558;
wire n_8108;
wire n_8158;
wire n_14990;
wire n_16076;
wire n_10464;
wire n_13054;
wire n_15923;
wire n_10446;
wire n_15010;
wire n_15957;
wire n_6553;
wire n_9715;
wire n_14166;
wire n_4905;
wire n_10219;
wire n_9016;
wire n_4508;
wire n_5897;
wire n_6261;
wire n_4894;
wire n_6659;
wire n_9399;
wire n_15615;
wire n_15215;
wire n_7351;
wire n_7256;
wire n_12967;
wire n_14458;
wire n_12907;
wire n_14353;
wire n_12020;
wire n_4141;
wire n_13877;
wire n_15368;
wire n_16211;
wire n_6893;
wire n_12377;
wire n_13272;
wire n_4422;
wire n_12007;
wire n_11087;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_15779;
wire n_5179;
wire n_10394;
wire n_15700;
wire n_6337;
wire n_5680;
wire n_6210;
wire n_7583;
wire n_14368;
wire n_5685;
wire n_13394;
wire n_15240;
wire n_5974;
wire n_10776;
wire n_14032;
wire n_14375;
wire n_10917;
wire n_5723;
wire n_14914;
wire n_15815;
wire n_15085;
wire n_5922;
wire n_6378;
wire n_14822;
wire n_5549;
wire n_13536;
wire n_9094;
wire n_13524;
wire n_8130;
wire n_15212;
wire n_11483;
wire n_14075;
wire n_14093;
wire n_4364;
wire n_14705;
wire n_12944;
wire n_9510;
wire n_11049;
wire n_7488;
wire n_16101;
wire n_7690;
wire n_12706;
wire n_14817;
wire n_12973;
wire n_12319;
wire n_4307;
wire n_14178;
wire n_14053;
wire n_6044;
wire n_15825;
wire n_16138;
wire n_12388;
wire n_6206;
wire n_7893;
wire n_11031;
wire n_9429;
wire n_14929;
wire n_11599;
wire n_4438;
wire n_11292;
wire n_15740;
wire n_6538;
wire n_11568;
wire n_15016;
wire n_7966;
wire n_6996;
wire n_5831;
wire n_9653;
wire n_4367;
wire n_5134;
wire n_11468;
wire n_13815;
wire n_7599;
wire n_9648;
wire n_7231;
wire n_14626;
wire n_10240;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_12470;
wire n_12711;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_15483;
wire n_8675;
wire n_12216;
wire n_9095;
wire n_7900;
wire n_11203;
wire n_5708;
wire n_8123;
wire n_9003;
wire n_9048;
wire n_16080;
wire n_12879;
wire n_14228;
wire n_13801;
wire n_5454;
wire n_14472;
wire n_13659;
wire n_4254;
wire n_10578;
wire n_14946;
wire n_11206;
wire n_12649;
wire n_12093;
wire n_13473;
wire n_8913;
wire n_9932;
wire n_15247;
wire n_8220;
wire n_12165;
wire n_15170;
wire n_11779;
wire n_13497;
wire n_16262;
wire n_9309;
wire n_8355;
wire n_12724;
wire n_9661;
wire n_14557;
wire n_9799;
wire n_12447;
wire n_5373;
wire n_7403;
wire n_6665;
wire n_8883;
wire n_15480;
wire n_15910;
wire n_13822;
wire n_7168;
wire n_10427;
wire n_15514;
wire n_15527;
wire n_4179;
wire n_11609;
wire n_11927;
wire n_10626;
wire n_11676;
wire n_6461;
wire n_6033;
wire n_10138;
wire n_15556;
wire n_6860;
wire n_9063;
wire n_7322;
wire n_10364;
wire n_6060;
wire n_10532;
wire n_5788;
wire n_5983;
wire n_15734;
wire n_15719;
wire n_9895;
wire n_10288;
wire n_6709;
wire n_11602;
wire n_15601;
wire n_13843;
wire n_11865;
wire n_15263;
wire n_12566;
wire n_5557;
wire n_12383;
wire n_6914;
wire n_8816;
wire n_15873;
wire n_4314;
wire n_8418;
wire n_14943;
wire n_5951;
wire n_4315;
wire n_5647;
wire n_16145;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_12035;
wire n_15684;
wire n_12212;
wire n_9110;
wire n_11427;
wire n_11613;
wire n_15739;
wire n_4442;
wire n_10668;
wire n_4857;
wire n_8739;
wire n_9969;
wire n_11375;
wire n_8927;
wire n_10398;
wire n_15749;
wire n_6009;
wire n_7221;
wire n_11870;
wire n_4637;
wire n_5523;
wire n_12053;
wire n_13250;
wire n_15004;
wire n_8243;
wire n_8798;
wire n_13228;
wire n_7963;
wire n_13893;
wire n_6382;
wire n_8423;
wire n_13869;
wire n_15278;
wire n_14326;
wire n_9028;
wire n_15335;
wire n_4296;
wire n_14699;
wire n_13100;
wire n_9654;
wire n_10683;
wire n_14232;
wire n_10249;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_9810;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_12852;
wire n_12123;
wire n_9701;
wire n_5392;
wire n_4714;
wire n_9270;
wire n_11373;
wire n_11878;
wire n_6418;
wire n_8548;
wire n_9437;
wire n_8996;
wire n_13185;
wire n_9483;
wire n_6263;
wire n_14593;
wire n_6731;
wire n_8156;
wire n_15774;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_16151;
wire n_6048;
wire n_13738;
wire n_7185;
wire n_10229;
wire n_12268;
wire n_5149;
wire n_9256;
wire n_5280;
wire n_4970;
wire n_10889;
wire n_11070;
wire n_6234;
wire n_16046;
wire n_4153;
wire n_14966;
wire n_8992;
wire n_5052;
wire n_7141;
wire n_5137;
wire n_15459;
wire n_11107;
wire n_14116;
wire n_13195;
wire n_12298;
wire n_6224;
wire n_12930;
wire n_8510;
wire n_5089;
wire n_11394;
wire n_5775;
wire n_9854;
wire n_15190;
wire n_9737;
wire n_8961;
wire n_12890;
wire n_14551;
wire n_9964;
wire n_11154;
wire n_14940;
wire n_4643;
wire n_9719;
wire n_6142;
wire n_10826;
wire n_6119;
wire n_10358;
wire n_12301;
wire n_15086;
wire n_13886;
wire n_6619;
wire n_11973;
wire n_13200;
wire n_4133;
wire n_11073;
wire n_13876;
wire n_6759;
wire n_6903;
wire n_7416;
wire n_15466;
wire n_6768;
wire n_5031;
wire n_7092;
wire n_7233;
wire n_4543;
wire n_14442;
wire n_4337;
wire n_9679;
wire n_9669;
wire n_11186;
wire n_12382;
wire n_5082;
wire n_4788;
wire n_10835;
wire n_12996;
wire n_13095;
wire n_15947;
wire n_4555;
wire n_5230;
wire n_4486;
wire n_10416;
wire n_12661;
wire n_8402;
wire n_8978;
wire n_14097;
wire n_7191;
wire n_15125;
wire n_14279;
wire n_6189;
wire n_5796;
wire n_15339;
wire n_13907;
wire n_9105;
wire n_13085;
wire n_14411;
wire n_9699;
wire n_11360;
wire n_5296;
wire n_5398;
wire n_6761;
wire n_14304;
wire n_9673;
wire n_15313;
wire n_10860;
wire n_11823;
wire n_4780;
wire n_4640;
wire n_8685;
wire n_10997;
wire n_9240;
wire n_15162;
wire n_7202;
wire n_14033;
wire n_5960;
wire n_7445;
wire n_9212;
wire n_5858;
wire n_13889;
wire n_5985;
wire n_8595;
wire n_10602;
wire n_15327;
wire n_12088;
wire n_11181;
wire n_9040;
wire n_9478;
wire n_10261;
wire n_10817;
wire n_12062;
wire n_12277;
wire n_14045;
wire n_4157;
wire n_9742;
wire n_11806;
wire n_7868;
wire n_10124;
wire n_13386;
wire n_16238;
wire n_7654;
wire n_8779;
wire n_5192;
wire n_15844;
wire n_4247;
wire n_5051;
wire n_10132;
wire n_15034;
wire n_5336;
wire n_8520;
wire n_4583;
wire n_14305;
wire n_8555;
wire n_12421;
wire n_10730;
wire n_9456;
wire n_6366;
wire n_11321;
wire n_6304;
wire n_4292;
wire n_9146;
wire n_11702;
wire n_7176;
wire n_14233;
wire n_14835;
wire n_8565;
wire n_8334;
wire n_13605;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_12133;
wire n_11970;
wire n_15167;
wire n_15083;
wire n_13283;
wire n_4773;
wire n_5028;
wire n_13596;
wire n_15912;
wire n_9573;
wire n_14983;
wire n_15257;
wire n_11286;
wire n_8030;
wire n_8513;
wire n_14511;
wire n_13746;
wire n_13327;
wire n_14550;
wire n_9379;
wire n_10948;
wire n_9219;
wire n_13534;
wire n_16186;
wire n_14056;
wire n_10927;
wire n_11496;
wire n_15356;
wire n_14151;
wire n_13149;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_8245;
wire n_13727;
wire n_13992;
wire n_14846;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_12186;
wire n_8753;
wire n_15230;
wire n_7527;
wire n_9706;
wire n_4856;
wire n_7948;
wire n_7096;
wire n_11863;
wire n_15776;
wire n_4216;
wire n_9206;
wire n_14139;
wire n_15002;
wire n_8485;
wire n_5596;
wire n_6482;
wire n_10118;
wire n_8106;
wire n_15585;
wire n_15847;
wire n_8325;
wire n_15329;
wire n_14619;
wire n_10875;
wire n_4864;
wire n_11225;
wire n_15018;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_15239;
wire n_10731;
wire n_4313;
wire n_14071;
wire n_15169;
wire n_11355;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_9434;
wire n_6229;
wire n_13113;
wire n_5933;
wire n_13198;
wire n_5536;
wire n_13097;
wire n_15256;
wire n_15928;
wire n_4798;
wire n_10350;
wire n_10654;
wire n_7293;
wire n_9874;
wire n_11261;
wire n_11862;
wire n_13369;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_12579;
wire n_4229;
wire n_5071;
wire n_5810;
wire n_10564;
wire n_12342;
wire n_13653;
wire n_14832;
wire n_14691;
wire n_11584;
wire n_9082;
wire n_7144;
wire n_12877;
wire n_12256;
wire n_4991;
wire n_13360;
wire n_11893;
wire n_10262;
wire n_11500;
wire n_11044;
wire n_7316;
wire n_7508;
wire n_13785;
wire n_9596;
wire n_15861;
wire n_8677;
wire n_15065;
wire n_5818;
wire n_5198;
wire n_11109;
wire n_12909;
wire n_13044;
wire n_12859;
wire n_16025;
wire n_10729;
wire n_9559;
wire n_15463;
wire n_9709;
wire n_10973;
wire n_15525;
wire n_4182;
wire n_8626;
wire n_12822;
wire n_7869;
wire n_13217;
wire n_13943;
wire n_10069;
wire n_10810;
wire n_16001;
wire n_12468;
wire n_8166;
wire n_9356;
wire n_14948;
wire n_5539;
wire n_4252;
wire n_5009;
wire n_12267;
wire n_15515;
wire n_12170;
wire n_12426;
wire n_15689;
wire n_15876;
wire n_6943;
wire n_10791;
wire n_12900;
wire n_10553;
wire n_14555;
wire n_6631;
wire n_5889;
wire n_12846;
wire n_8602;
wire n_9609;
wire n_7151;
wire n_10284;
wire n_15467;
wire n_7762;
wire n_13469;
wire n_15346;
wire n_13840;
wire n_13836;
wire n_5632;
wire n_12855;
wire n_11501;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_16260;
wire n_13569;
wire n_4446;
wire n_5613;
wire n_4662;
wire n_7472;
wire n_9342;
wire n_14229;
wire n_4800;
wire n_14425;
wire n_15324;
wire n_7075;
wire n_13076;
wire n_14917;
wire n_5427;
wire n_12234;
wire n_4440;
wire n_4425;
wire n_6770;
wire n_14317;
wire n_5450;
wire n_7611;
wire n_11437;
wire n_7796;
wire n_6508;
wire n_14682;
wire n_7989;
wire n_13320;
wire n_8047;
wire n_12120;
wire n_13082;
wire n_15863;
wire n_15064;
wire n_9233;
wire n_10474;
wire n_7936;
wire n_10694;
wire n_10529;
wire n_13117;
wire n_15622;
wire n_4781;
wire n_12042;
wire n_6031;
wire n_14328;
wire n_15457;
wire n_5124;
wire n_16084;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_11722;
wire n_4828;
wire n_12568;
wire n_14444;
wire n_12149;
wire n_15138;
wire n_8800;
wire n_4652;
wire n_12278;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_10622;
wire n_9435;
wire n_13318;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_9557;
wire n_11639;
wire n_9551;
wire n_8955;
wire n_8039;
wire n_8193;
wire n_12231;
wire n_12116;
wire n_9073;
wire n_13677;
wire n_7546;
wire n_8432;
wire n_15343;
wire n_14422;
wire n_5904;
wire n_11997;
wire n_14876;
wire n_16088;
wire n_6628;
wire n_5318;
wire n_8684;
wire n_5374;
wire n_10270;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_16069;
wire n_13158;
wire n_7407;
wire n_12014;
wire n_13230;
wire n_9388;
wire n_10463;
wire n_9721;
wire n_11731;
wire n_14061;
wire n_4863;
wire n_10880;
wire n_11610;
wire n_12097;
wire n_14612;
wire n_12363;
wire n_13115;
wire n_15599;
wire n_13427;
wire n_5463;
wire n_6328;
wire n_11498;
wire n_6929;
wire n_12008;
wire n_11509;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_15097;
wire n_14401;
wire n_14034;
wire n_15518;
wire n_15820;
wire n_13559;
wire n_15400;
wire n_6012;
wire n_15723;
wire n_7481;
wire n_11447;
wire n_4429;
wire n_6484;
wire n_5435;
wire n_11706;
wire n_5053;
wire n_7182;
wire n_14498;
wire n_11055;
wire n_14517;
wire n_10689;
wire n_9507;
wire n_5476;
wire n_5483;
wire n_12534;
wire n_9539;
wire n_8617;
wire n_14297;
wire n_7605;
wire n_8591;
wire n_8090;
wire n_15513;
wire n_9268;
wire n_5511;
wire n_9718;
wire n_8661;
wire n_13512;
wire n_10068;
wire n_15330;
wire n_6639;
wire n_11258;
wire n_9672;
wire n_12748;
wire n_11168;
wire n_9890;
wire n_12272;
wire n_9187;
wire n_9572;
wire n_16272;
wire n_12148;
wire n_10363;
wire n_6124;
wire n_16130;
wire n_12615;
wire n_12142;
wire n_16164;
wire n_13201;
wire n_9527;
wire n_11234;
wire n_15375;
wire n_9949;
wire n_13388;
wire n_14484;
wire n_7423;
wire n_13674;
wire n_15115;
wire n_7375;
wire n_7076;
wire n_16269;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_8811;
wire n_13858;
wire n_9952;
wire n_11612;
wire n_7736;
wire n_6435;
wire n_13949;
wire n_10888;
wire n_12714;
wire n_13782;
wire n_14486;
wire n_14759;
wire n_5829;
wire n_14580;
wire n_7419;
wire n_13612;
wire n_6600;
wire n_14087;
wire n_13681;
wire n_7010;
wire n_13700;
wire n_14421;
wire n_16095;
wire n_14193;
wire n_10277;
wire n_15242;
wire n_5881;
wire n_9798;
wire n_4694;
wire n_11895;
wire n_8192;
wire n_9251;
wire n_4664;
wire n_6201;
wire n_10537;
wire n_14703;
wire n_14684;
wire n_14653;
wire n_8573;
wire n_4633;
wire n_13770;
wire n_10807;
wire n_14048;
wire n_13920;
wire n_7918;
wire n_9546;
wire n_10331;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_13130;
wire n_6735;
wire n_9181;
wire n_9602;
wire n_12812;
wire n_13377;
wire n_15846;
wire n_11455;
wire n_6803;
wire n_4288;
wire n_14816;
wire n_10981;
wire n_5894;
wire n_13750;
wire n_9635;
wire n_11868;
wire n_4511;
wire n_12639;
wire n_12189;
wire n_14063;
wire n_15542;
wire n_14521;
wire n_4675;
wire n_13701;
wire n_11934;
wire n_13518;
wire n_5419;
wire n_8339;
wire n_14737;
wire n_11969;
wire n_13668;
wire n_4289;
wire n_4972;
wire n_11571;
wire n_7346;
wire n_6036;
wire n_9405;
wire n_15255;
wire n_12428;
wire n_12069;
wire n_14384;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_10780;
wire n_10158;
wire n_11481;
wire n_6102;
wire n_5077;
wire n_16173;
wire n_14276;
wire n_12057;
wire n_12050;
wire n_13587;
wire n_9726;
wire n_13488;
wire n_15852;
wire n_8804;
wire n_9577;
wire n_6650;
wire n_10024;
wire n_6573;
wire n_11774;
wire n_6904;
wire n_15271;
wire n_12214;
wire n_13805;
wire n_6329;
wire n_7385;
wire n_15425;
wire n_9802;
wire n_6244;
wire n_4846;
wire n_9540;
wire n_6204;
wire n_9250;
wire n_13365;
wire n_13767;
wire n_13972;
wire n_12381;
wire n_10191;
wire n_5225;
wire n_7295;
wire n_7824;
wire n_12157;
wire n_7148;
wire n_13938;
wire n_9171;
wire n_7169;
wire n_16054;
wire n_13443;
wire n_15297;
wire n_9350;
wire n_11257;
wire n_12330;
wire n_6756;
wire n_4805;
wire n_9441;
wire n_7600;
wire n_15268;
wire n_15838;
wire n_15814;
wire n_9124;
wire n_10675;
wire n_5826;
wire n_8697;
wire n_11598;
wire n_9626;
wire n_14011;
wire n_14645;
wire n_4822;
wire n_11327;
wire n_6946;
wire n_12926;
wire n_7947;
wire n_8645;
wire n_5931;
wire n_8820;
wire n_8146;
wire n_9408;
wire n_14712;
wire n_4635;
wire n_8154;
wire n_7847;
wire n_12824;
wire n_12392;
wire n_13094;
wire n_5532;
wire n_14545;
wire n_7311;
wire n_6804;
wire n_16189;
wire n_6179;
wire n_5441;
wire n_14103;
wire n_6059;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_14976;
wire n_8063;
wire n_13798;
wire n_14677;
wire n_8406;
wire n_15580;
wire n_6427;
wire n_14474;
wire n_14459;
wire n_4281;
wire n_5994;
wire n_12070;
wire n_8480;
wire n_11265;
wire n_14037;
wire n_11788;
wire n_14112;
wire n_14811;
wire n_9754;
wire n_10477;
wire n_4419;
wire n_14296;
wire n_11904;
wire n_8849;
wire n_13071;
wire n_5405;
wire n_9750;
wire n_10296;
wire n_7660;
wire n_13676;
wire n_13735;
wire n_14127;
wire n_5365;
wire n_9529;
wire n_9566;
wire n_5772;
wire n_11901;
wire n_12848;
wire n_10339;
wire n_15528;
wire n_6442;
wire n_8241;
wire n_10307;
wire n_10606;
wire n_6188;
wire n_12161;
wire n_16249;
wire n_10066;
wire n_11755;
wire n_4906;
wire n_11754;
wire n_15610;
wire n_6846;
wire n_13825;
wire n_10054;
wire n_4630;
wire n_8261;
wire n_10343;
wire n_6840;
wire n_6645;
wire n_15020;
wire n_8535;
wire n_8348;
wire n_4829;
wire n_13985;
wire n_6749;
wire n_12238;
wire n_6915;
wire n_12956;
wire n_12320;
wire n_8138;
wire n_7831;
wire n_13342;
wire n_11413;
wire n_13953;
wire n_10652;
wire n_13040;
wire n_5259;
wire n_15735;
wire n_8702;
wire n_11601;
wire n_7455;
wire n_8273;
wire n_14250;
wire n_10944;
wire n_6247;
wire n_5921;
wire n_10367;
wire n_15365;
wire n_11129;
wire n_11710;
wire n_4966;
wire n_14602;
wire n_8235;
wire n_15510;
wire n_13685;
wire n_6104;
wire n_15476;
wire n_9940;
wire n_15444;
wire n_8294;
wire n_12476;
wire n_4188;
wire n_10016;
wire n_15273;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_9283;
wire n_6205;
wire n_11010;
wire n_8349;
wire n_15901;
wire n_4825;
wire n_9822;
wire n_10036;
wire n_15199;
wire n_9607;
wire n_9443;
wire n_7497;
wire n_16201;
wire n_10749;
wire n_7315;
wire n_10166;
wire n_8429;
wire n_13765;
wire n_6939;
wire n_16214;
wire n_7887;
wire n_10419;
wire n_15726;
wire n_9298;
wire n_5884;
wire n_15470;
wire n_5006;
wire n_14200;
wire n_4882;
wire n_10006;
wire n_5728;
wire n_13334;
wire n_14902;
wire n_4878;
wire n_8486;
wire n_11240;
wire n_9052;
wire n_6706;
wire n_13123;
wire n_12154;
wire n_16149;
wire n_7431;
wire n_8140;
wire n_11734;
wire n_14450;
wire n_15276;
wire n_14477;
wire n_4202;
wire n_6909;
wire n_13933;
wire n_5679;
wire n_6487;
wire n_8117;
wire n_12668;
wire n_15143;
wire n_15633;
wire n_10348;
wire n_13884;
wire n_7521;
wire n_10058;
wire n_5141;
wire n_6627;
wire n_4503;
wire n_15975;
wire n_8129;
wire n_10355;
wire n_11156;
wire n_7253;
wire n_5208;
wire n_9535;
wire n_13511;
wire n_5113;
wire n_10304;
wire n_12928;
wire n_11955;
wire n_5205;
wire n_4249;
wire n_15110;
wire n_9943;
wire n_7569;
wire n_12538;
wire n_13745;
wire n_12151;
wire n_16202;
wire n_10966;
wire n_14697;
wire n_13112;
wire n_13646;
wire n_12130;
wire n_14608;
wire n_15049;
wire n_7452;
wire n_12409;
wire n_13031;
wire n_6551;
wire n_12350;
wire n_15767;
wire n_7972;
wire n_8672;
wire n_13455;
wire n_15411;
wire n_7505;
wire n_13993;
wire n_14280;
wire n_13946;
wire n_6516;
wire n_14567;
wire n_10060;
wire n_7524;
wire n_15763;
wire n_13931;
wire n_4196;
wire n_11270;
wire n_8934;
wire n_14961;
wire n_11020;
wire n_7318;
wire n_9977;
wire n_10722;
wire n_7411;
wire n_13314;
wire n_7326;
wire n_13378;
wire n_5667;
wire n_9555;
wire n_15980;
wire n_13618;
wire n_10957;
wire n_14277;
wire n_8847;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_11344;
wire n_15446;
wire n_14952;
wire n_5879;
wire n_6500;
wire n_11303;
wire n_5027;
wire n_12847;
wire n_14340;
wire n_5688;
wire n_9030;
wire n_5825;
wire n_11216;
wire n_15652;
wire n_8221;
wire n_13638;
wire n_7573;
wire n_6630;
wire n_14886;
wire n_5759;
wire n_5629;
wire n_10409;
wire n_13167;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_13758;
wire n_5999;
wire n_9590;
wire n_14646;
wire n_11511;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_10322;
wire n_11339;
wire n_11346;
wire n_11829;
wire n_12680;
wire n_5377;
wire n_6180;
wire n_12530;
wire n_11581;
wire n_8225;
wire n_7453;
wire n_4355;
wire n_12163;
wire n_16184;
wire n_14131;
wire n_7932;
wire n_9651;
wire n_7890;
wire n_5599;
wire n_10825;
wire n_16199;
wire n_16129;
wire n_15575;
wire n_6004;
wire n_9583;
wire n_9763;
wire n_10349;
wire n_9944;
wire n_13709;
wire n_13035;
wire n_6652;
wire n_9888;
wire n_7183;
wire n_4155;
wire n_4278;
wire n_10040;
wire n_10636;
wire n_4710;
wire n_10844;
wire n_12738;
wire n_6275;
wire n_6395;
wire n_6403;
wire n_9862;
wire n_14622;
wire n_6578;
wire n_4542;
wire n_5451;
wire n_15267;
wire n_4326;
wire n_9966;
wire n_15455;
wire n_10242;
wire n_6350;
wire n_16023;
wire n_5460;
wire n_4685;
wire n_16115;
wire n_9936;
wire n_6141;
wire n_8559;
wire n_11165;
wire n_6875;
wire n_7189;
wire n_9617;
wire n_10727;
wire n_9341;
wire n_6194;
wire n_14984;
wire n_14864;
wire n_15000;
wire n_8689;
wire n_11231;
wire n_9749;
wire n_5517;
wire n_9629;
wire n_13654;
wire n_5807;
wire n_14985;
wire n_15944;
wire n_11448;
wire n_12227;
wire n_5426;
wire n_6475;
wire n_12525;
wire n_10679;
wire n_11132;
wire n_10524;
wire n_12282;
wire n_5693;
wire n_13426;
wire n_5695;
wire n_12932;
wire n_14849;
wire n_4123;
wire n_13799;
wire n_14207;
wire n_16064;
wire n_4294;
wire n_8330;
wire n_10011;
wire n_12037;
wire n_6502;
wire n_10030;
wire n_6944;
wire n_11410;
wire n_14365;
wire n_4452;
wire n_15147;
wire n_8304;
wire n_9349;
wire n_13480;
wire n_15658;
wire n_5587;
wire n_4722;
wire n_11267;
wire n_13780;
wire n_6318;
wire n_10119;
wire n_11348;
wire n_11940;
wire n_13613;
wire n_10845;
wire n_8163;
wire n_6805;
wire n_11947;
wire n_4164;
wire n_4126;
wire n_7240;
wire n_5030;
wire n_15630;
wire n_8907;
wire n_14227;
wire n_5674;
wire n_7499;
wire n_9423;
wire n_5584;
wire n_12424;
wire n_5320;
wire n_15227;
wire n_6075;
wire n_10063;
wire n_12942;
wire n_6559;
wire n_9038;
wire n_8777;
wire n_11149;
wire n_8698;
wire n_10709;
wire n_6068;
wire n_12236;
wire n_4366;
wire n_6248;
wire n_6541;
wire n_11436;
wire n_9034;
wire n_5125;
wire n_4922;
wire n_11909;
wire n_12547;
wire n_13554;
wire n_6066;
wire n_6080;
wire n_14372;
wire n_13421;
wire n_4733;
wire n_7927;
wire n_8928;
wire n_13967;
wire n_13150;
wire n_13014;
wire n_7219;
wire n_10526;
wire n_11439;
wire n_8081;
wire n_12192;
wire n_12747;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_11462;
wire n_14564;
wire n_16155;
wire n_7063;
wire n_7402;
wire n_9676;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_7382;
wire n_8384;
wire n_10861;
wire n_5238;
wire n_13795;
wire n_8650;
wire n_14729;
wire n_14989;
wire n_11272;
wire n_14992;
wire n_14044;
wire n_12989;
wire n_5906;
wire n_16005;
wire n_7767;
wire n_5732;
wire n_4194;
wire n_11759;
wire n_14431;
wire n_10494;
wire n_16258;
wire n_5780;
wire n_10478;
wire n_11061;
wire n_11653;
wire n_8284;
wire n_10534;
wire n_8374;
wire n_5556;
wire n_6006;
wire n_6474;
wire n_13662;
wire n_13864;
wire n_5743;
wire n_6481;
wire n_10078;
wire n_11478;
wire n_5633;
wire n_12273;
wire n_7510;
wire n_15475;
wire n_9041;
wire n_15809;
wire n_9995;
wire n_12200;
wire n_6022;
wire n_6991;
wire n_10629;
wire n_13863;
wire n_7434;
wire n_5950;
wire n_9035;
wire n_13926;
wire n_9011;
wire n_14240;
wire n_4204;
wire n_7691;
wire n_11748;
wire n_5323;
wire n_7745;
wire n_14331;
wire n_14165;
wire n_9135;
wire n_6744;
wire n_9776;
wire n_15055;
wire n_5705;
wire n_12660;
wire n_11867;
wire n_14192;
wire n_6927;
wire n_14678;
wire n_15673;
wire n_7335;
wire n_12400;
wire n_13072;
wire n_14708;
wire n_10472;
wire n_10695;
wire n_10286;
wire n_9413;
wire n_4996;
wire n_9107;
wire n_4411;
wire n_15823;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_15713;
wire n_6116;
wire n_9548;
wire n_8074;
wire n_15117;
wire n_15479;
wire n_14246;
wire n_8780;
wire n_15631;
wire n_7956;
wire n_5510;
wire n_15536;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_9775;
wire n_13857;
wire n_16143;
wire n_13033;
wire n_12922;
wire n_8580;
wire n_15736;
wire n_5440;
wire n_12193;
wire n_9288;
wire n_4163;
wire n_15594;
wire n_16036;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_15047;
wire n_12243;
wire n_5513;
wire n_10218;
wire n_5875;
wire n_14671;
wire n_8358;
wire n_7734;
wire n_4262;
wire n_10441;
wire n_9305;
wire n_9093;
wire n_11764;
wire n_7671;
wire n_13696;
wire n_15200;
wire n_15924;
wire n_16045;
wire n_12950;
wire n_10043;
wire n_4832;
wire n_8033;
wire n_5197;
wire n_6485;
wire n_13041;
wire n_15021;
wire n_5848;
wire n_5834;
wire n_14269;
wire n_7926;
wire n_11882;
wire n_5784;
wire n_13418;
wire n_14820;
wire n_12250;
wire n_5128;
wire n_10628;
wire n_13498;
wire n_14290;
wire n_15806;
wire n_8643;
wire n_15715;
wire n_14792;
wire n_11787;
wire n_12403;
wire n_5618;
wire n_11539;
wire n_15760;
wire n_15099;
wire n_10440;
wire n_15618;
wire n_10134;
wire n_12904;
wire n_6495;
wire n_7528;
wire n_14669;
wire n_12444;
wire n_11163;
wire n_6209;
wire n_16107;
wire n_4672;
wire n_8094;
wire n_11695;
wire n_9425;
wire n_13489;
wire n_14520;
wire n_15225;
wire n_13373;
wire n_13739;
wire n_10317;
wire n_11730;
wire n_13101;
wire n_11916;
wire n_13723;
wire n_13000;
wire n_13556;
wire n_15238;
wire n_14821;
wire n_11311;
wire n_14525;
wire n_7413;
wire n_14435;
wire n_7993;
wire n_11980;
wire n_7821;
wire n_11151;
wire n_14238;
wire n_7620;
wire n_15520;
wire n_13153;
wire n_12837;
wire n_12356;
wire n_15195;
wire n_13091;
wire n_13937;
wire n_13032;
wire n_6274;
wire n_5157;
wire n_12764;
wire n_14654;
wire n_4496;
wire n_9347;
wire n_12269;
wire n_14556;
wire n_12079;
wire n_14687;
wire n_13508;
wire n_10706;
wire n_4596;
wire n_5178;
wire n_9420;
wire n_13350;
wire n_13901;
wire n_12972;
wire n_6237;
wire n_13635;
wire n_4628;
wire n_6802;
wire n_13224;
wire n_7343;
wire n_16163;
wire n_5982;
wire n_8477;
wire n_13306;
wire n_9344;
wire n_14657;
wire n_7109;
wire n_12438;
wire n_8028;
wire n_15435;
wire n_16082;
wire n_14245;
wire n_14254;
wire n_12125;
wire n_14993;
wire n_12554;
wire n_10297;
wire n_15608;
wire n_6155;
wire n_7506;
wire n_9530;
wire n_6809;
wire n_10160;
wire n_6099;
wire n_10849;
wire n_10605;
wire n_11296;
wire n_13259;
wire n_14217;
wire n_8530;
wire n_14343;
wire n_15165;
wire n_10379;
wire n_9446;
wire n_15434;
wire n_5529;
wire n_15094;
wire n_16234;
wire n_7561;
wire n_6349;
wire n_13278;
wire n_11081;
wire n_8500;
wire n_6716;
wire n_8713;
wire n_12860;
wire n_14554;
wire n_7885;
wire n_8297;
wire n_14100;
wire n_15410;
wire n_6905;
wire n_15519;
wire n_15616;
wire n_8926;
wire n_9865;
wire n_14974;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_11230;
wire n_5824;
wire n_8025;
wire n_10282;
wire n_5354;
wire n_15498;
wire n_7898;
wire n_11357;
wire n_13179;
wire n_11027;
wire n_10458;
wire n_12206;
wire n_11393;
wire n_6203;
wire n_12947;
wire n_6407;
wire n_14468;
wire n_4230;
wire n_11892;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_7070;
wire n_9025;
wire n_5276;
wire n_11105;
wire n_9713;
wire n_11160;
wire n_13043;
wire n_14675;
wire n_4659;
wire n_8293;
wire n_13962;
wire n_7299;
wire n_5196;
wire n_10382;
wire n_8029;
wire n_14892;
wire n_13468;
wire n_9314;
wire n_12270;
wire n_15830;
wire n_15325;
wire n_6960;
wire n_14235;
wire n_8880;
wire n_7249;
wire n_9660;
wire n_5763;
wire n_15062;
wire n_13018;
wire n_12739;
wire n_6061;
wire n_13831;
wire n_16105;
wire n_9769;
wire n_8471;
wire n_15031;
wire n_5701;
wire n_7002;
wire n_14529;
wire n_15940;
wire n_15688;
wire n_12906;
wire n_12490;
wire n_9902;
wire n_6273;
wire n_14424;
wire n_7094;
wire n_7396;
wire n_12751;
wire n_11397;
wire n_8726;
wire n_10640;
wire n_8977;
wire n_7018;
wire n_11897;
wire n_14949;
wire n_10522;
wire n_6746;
wire n_15248;
wire n_10691;
wire n_12650;
wire n_10764;
wire n_10244;
wire n_10914;
wire n_13348;
wire n_10272;
wire n_8316;
wire n_6174;
wire n_15070;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_14690;
wire n_15116;
wire n_13415;
wire n_5907;
wire n_7297;
wire n_4339;
wire n_7730;
wire n_10980;
wire n_12279;
wire n_13265;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_14916;
wire n_6279;
wire n_5895;
wire n_9410;
wire n_9588;
wire n_12242;
wire n_4169;
wire n_10071;
wire n_8610;
wire n_4253;
wire n_7637;
wire n_12588;
wire n_16241;
wire n_6131;
wire n_5478;
wire n_13382;
wire n_10176;
wire n_6113;
wire n_9740;
wire n_14767;
wire n_6477;
wire n_5384;
wire n_7486;
wire n_6575;
wire n_11719;
wire n_5283;
wire n_9910;
wire n_5961;
wire n_7544;
wire n_7613;
wire n_9061;
wire n_15178;
wire n_15810;
wire n_7995;
wire n_9941;
wire n_14794;
wire n_8113;
wire n_9579;
wire n_5686;
wire n_6391;
wire n_10254;
wire n_14446;
wire n_8724;
wire n_14121;
wire n_10332;
wire n_7140;
wire n_14955;
wire n_15769;
wire n_15877;
wire n_16117;
wire n_12775;
wire n_12173;
wire n_10938;
wire n_10257;
wire n_9668;
wire n_6252;
wire n_6426;
wire n_14031;
wire n_4681;
wire n_11956;
wire n_8253;
wire n_12167;
wire n_15091;
wire n_9258;
wire n_15033;
wire n_9228;
wire n_13461;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_10214;
wire n_11874;
wire n_5094;
wire n_10195;
wire n_14918;
wire n_16096;
wire n_13979;
wire n_9598;
wire n_10354;
wire n_7741;
wire n_12060;
wire n_4295;
wire n_10436;
wire n_11450;
wire n_11723;
wire n_6668;
wire n_9311;
wire n_11982;
wire n_14062;
wire n_14448;
wire n_11822;
wire n_12179;
wire n_11522;
wire n_8232;
wire n_12842;
wire n_8803;
wire n_10866;
wire n_4473;
wire n_14715;
wire n_4619;
wire n_12499;
wire n_6670;
wire n_5371;
wire n_4398;
wire n_5026;
wire n_5350;
wire n_7679;
wire n_8818;
wire n_12693;
wire n_14906;
wire n_10811;
wire n_7698;
wire n_10073;
wire n_14873;
wire n_6962;
wire n_14187;
wire n_6779;
wire n_9608;
wire n_5286;
wire n_10164;
wire n_4449;
wire n_14779;
wire n_13172;
wire n_4607;
wire n_10205;
wire n_5676;
wire n_16065;
wire n_14716;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_10515;
wire n_7800;
wire n_12326;
wire n_15438;
wire n_4266;
wire n_6336;
wire n_13713;
wire n_4407;
wire n_15384;
wire n_4695;
wire n_6503;
wire n_15362;
wire n_7835;
wire n_12542;
wire n_16040;
wire n_15080;
wire n_13650;
wire n_15187;
wire n_6049;
wire n_5885;
wire n_11499;
wire n_14390;
wire n_9818;
wire n_7100;
wire n_7243;
wire n_4777;
wire n_5243;
wire n_11034;
wire n_7415;
wire n_14747;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_9433;
wire n_14004;
wire n_11746;
wire n_11698;
wire n_15462;
wire n_8795;
wire n_10430;
wire n_12934;
wire n_10338;
wire n_11560;
wire n_9599;
wire n_8674;
wire n_9186;
wire n_14054;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_13941;
wire n_15805;
wire n_5760;
wire n_12483;
wire n_7747;
wire n_9935;
wire n_14263;
wire n_12404;
wire n_12258;
wire n_4415;
wire n_5110;
wire n_8966;
wire n_11871;
wire n_14694;
wire n_7552;
wire n_14872;
wire n_14826;
wire n_10500;
wire n_9537;
wire n_10018;
wire n_9552;
wire n_9421;
wire n_15537;
wire n_6998;
wire n_7395;
wire n_13209;
wire n_15888;
wire n_5844;
wire n_10359;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_12823;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_14775;
wire n_15795;
wire n_6609;
wire n_10548;
wire n_7635;
wire n_4408;
wire n_12905;
wire n_10291;
wire n_15124;
wire n_8567;
wire n_8259;
wire n_15638;
wire n_10667;
wire n_12274;
wire n_12849;
wire n_11167;
wire n_11297;
wire n_4976;
wire n_9473;
wire n_10208;
wire n_6525;
wire n_11183;
wire n_9469;
wire n_11285;
wire n_5938;
wire n_14270;
wire n_7274;
wire n_11740;
wire n_8578;
wire n_14859;
wire n_10757;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_15428;
wire n_14679;
wire n_13975;
wire n_6494;
wire n_15680;
wire n_4574;
wire n_15624;
wire n_8160;
wire n_8980;
wire n_6132;
wire n_10631;
wire n_10864;
wire n_11136;
wire n_4557;
wire n_11434;
wire n_8336;
wire n_11133;
wire n_14710;
wire n_14781;
wire n_13711;
wire n_7788;
wire n_5548;
wire n_16261;
wire n_6974;
wire n_13477;
wire n_10748;
wire n_14783;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_15087;
wire n_9909;
wire n_15718;
wire n_4624;
wire n_16024;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_12303;
wire n_6562;
wire n_4902;
wire n_12002;
wire n_15512;
wire n_8600;
wire n_8229;
wire n_12442;
wire n_4686;
wire n_9236;
wire n_9751;
wire n_10751;
wire n_14649;
wire n_7794;
wire n_13579;
wire n_10434;
wire n_16079;
wire n_9369;
wire n_13634;
wire n_14844;
wire n_4338;
wire n_13987;
wire n_12597;
wire n_5917;
wire n_15853;
wire n_9757;
wire n_12419;
wire n_6965;
wire n_11886;
wire n_14804;
wire n_14210;
wire n_8761;
wire n_15732;
wire n_14316;
wire n_7630;
wire n_15607;
wire n_11804;
wire n_13262;
wire n_4161;
wire n_14673;
wire n_9076;
wire n_6168;
wire n_5304;
wire n_15943;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_5355;
wire n_9729;
wire n_13706;
wire n_11531;
wire n_12943;
wire n_13543;
wire n_6284;
wire n_12039;
wire n_15024;
wire n_16203;
wire n_10663;
wire n_14393;
wire n_5321;
wire n_14144;
wire n_7454;
wire n_10263;
wire n_12295;
wire n_8473;
wire n_9366;
wire n_4772;
wire n_11883;
wire n_6931;
wire n_6521;
wire n_8351;
wire n_5915;
wire n_7276;
wire n_11792;
wire n_6379;
wire n_16059;
wire n_9647;
wire n_12410;
wire n_7085;
wire n_6306;
wire n_12938;
wire n_7753;
wire n_12891;
wire n_13493;
wire n_12304;
wire n_6834;
wire n_4716;
wire n_4654;
wire n_8948;
wire n_13166;
wire n_14760;
wire n_13541;
wire n_15412;
wire n_15695;
wire n_12572;
wire n_10318;
wire n_13551;
wire n_14356;
wire n_5116;
wire n_10740;
wire n_15131;
wire n_7225;
wire n_11634;
wire n_15535;
wire n_7541;
wire n_11039;
wire n_10062;
wire n_7913;
wire n_10128;
wire n_8020;
wire n_7946;
wire n_8944;
wire n_10717;
wire n_11965;
wire n_5500;
wire n_13890;
wire n_9275;
wire n_4622;
wire n_15158;
wire n_15265;
wire n_4757;
wire n_15955;
wire n_9520;
wire n_6471;
wire n_6949;
wire n_11477;
wire n_5669;
wire n_5672;
wire n_5621;
wire n_9493;
wire n_6760;
wire n_14852;
wire n_15006;
wire n_8875;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_9102;
wire n_14128;
wire n_5515;
wire n_11588;
wire n_11818;
wire n_6589;
wire n_11592;
wire n_4570;
wire n_10721;
wire n_7014;
wire n_10945;
wire n_12290;
wire n_9801;
wire n_11742;
wire n_13902;
wire n_12718;
wire n_7920;
wire n_11312;
wire n_5559;
wire n_8649;
wire n_5337;
wire n_11235;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_14185;
wire n_7841;
wire n_9424;
wire n_10013;
wire n_7324;
wire n_7160;
wire n_9333;
wire n_16099;
wire n_8205;
wire n_11505;
wire n_12469;
wire n_15387;
wire n_15986;
wire n_6046;
wire n_11673;
wire n_7054;
wire n_4493;
wire n_8975;
wire n_6055;
wire n_7161;
wire n_9004;
wire n_6364;
wire n_8919;
wire n_6091;
wire n_6348;
wire n_9987;
wire n_8440;
wire n_11555;
wire n_13917;
wire n_15102;
wire n_15663;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_9860;
wire n_10565;
wire n_14327;
wire n_7837;
wire n_9670;
wire n_6788;
wire n_13548;
wire n_13903;
wire n_11241;
wire n_6144;
wire n_15730;
wire n_15868;
wire n_10389;
wire n_9200;
wire n_5528;
wire n_15035;
wire n_7806;
wire n_5605;
wire n_15905;
wire n_12336;
wire n_13080;
wire n_9417;
wire n_11059;
wire n_6896;
wire n_15534;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_15681;
wire n_12248;
wire n_12931;
wire n_14047;
wire n_11066;
wire n_16200;
wire n_4901;
wire n_8757;
wire n_10020;
wire n_7201;
wire n_13408;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_9386;
wire n_12713;
wire n_8897;
wire n_12810;
wire n_7676;
wire n_8177;
wire n_11683;
wire n_13733;
wire n_14311;
wire n_5467;
wire n_7241;
wire n_15612;
wire n_14147;
wire n_5493;
wire n_9207;
wire n_13592;
wire n_6285;
wire n_10356;
wire n_12717;
wire n_13915;
wire n_7644;
wire n_9276;
wire n_4602;
wire n_7816;
wire n_8829;
wire n_12119;
wire n_14186;
wire n_14149;
wire n_4900;
wire n_10110;
wire n_6748;
wire n_11275;
wire n_7430;
wire n_14540;
wire n_13589;
wire n_16267;
wire n_11329;
wire n_8638;
wire n_14272;
wire n_13189;
wire n_13260;
wire n_5901;
wire n_9980;
wire n_11923;
wire n_11718;
wire n_6582;
wire n_7724;
wire n_5360;
wire n_10501;
wire n_7269;
wire n_15160;
wire n_16058;
wire n_12003;
wire n_7047;
wire n_12292;
wire n_16113;
wire n_10908;
wire n_9176;
wire n_6937;
wire n_4363;
wire n_12405;
wire n_9728;
wire n_11809;
wire n_10777;
wire n_8101;
wire n_13712;
wire n_15549;
wire n_8687;
wire n_5439;
wire n_6115;
wire n_9866;
wire n_14685;
wire n_8721;
wire n_8749;
wire n_12780;
wire n_13349;
wire n_9465;
wire n_13277;
wire n_11975;
wire n_8937;
wire n_6272;
wire n_7067;
wire n_12087;
wire n_13233;
wire n_13808;
wire n_14478;
wire n_4736;
wire n_5250;
wire n_4842;
wire n_12662;
wire n_10965;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_11441;
wire n_12416;
wire n_14895;
wire n_15555;
wire n_9702;
wire n_10998;
wire n_13503;
wire n_6607;
wire n_12854;
wire n_4439;
wire n_4985;
wire n_12936;
wire n_9000;
wire n_13056;
wire n_13300;
wire n_7117;
wire n_11743;
wire n_12765;
wire n_13087;
wire n_9610;
wire n_5471;
wire n_4660;
wire n_8503;
wire n_10082;
wire n_10870;
wire n_12796;
wire n_11914;
wire n_15364;
wire n_6446;
wire n_10756;
wire n_5497;
wire n_9139;
wire n_13287;
wire n_5519;
wire n_6071;
wire n_12028;
wire n_8315;
wire n_11175;
wire n_15563;
wire n_10411;
wire n_6849;
wire n_6807;
wire n_15236;
wire n_11753;
wire n_8197;
wire n_13726;
wire n_11790;
wire n_9407;
wire n_12294;
wire n_6616;
wire n_6719;
wire n_14621;
wire n_15883;
wire n_10423;
wire n_4814;
wire n_8019;
wire n_8801;
wire n_12190;
wire n_14396;
wire n_15134;
wire n_6178;
wire n_11249;
wire n_8707;
wire n_6677;
wire n_11791;
wire n_12786;
wire n_7875;
wire n_15983;
wire n_5502;
wire n_8962;
wire n_13665;
wire n_8931;
wire n_8248;
wire n_14177;
wire n_7550;
wire n_14533;
wire n_8554;
wire n_13242;
wire n_11879;
wire n_13900;
wire n_15269;
wire n_10782;
wire n_13837;
wire n_7302;
wire n_6191;
wire n_12386;
wire n_13121;
wire n_13679;
wire n_13680;
wire n_9357;
wire n_9477;
wire n_11911;
wire n_16274;
wire n_13734;
wire n_14591;
wire n_15756;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_11842;
wire n_5706;
wire n_12746;
wire n_14023;
wire n_13047;
wire n_11320;
wire n_11304;
wire n_15728;
wire n_7292;
wire n_13146;
wire n_7804;
wire n_10251;
wire n_15780;
wire n_12128;
wire n_11776;
wire n_14544;
wire n_11471;
wire n_14904;
wire n_5098;
wire n_15253;
wire n_13475;
wire n_6000;
wire n_6774;
wire n_9289;
wire n_11794;
wire n_6443;
wire n_9828;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_13236;
wire n_15656;
wire n_7248;
wire n_10737;
wire n_10475;
wire n_6647;
wire n_11198;
wire n_8040;
wire n_13336;
wire n_5466;
wire n_14465;
wire n_6941;
wire n_7239;
wire n_9797;
wire n_15015;
wire n_6552;
wire n_7826;
wire n_10665;
wire n_9981;
wire n_6094;
wire n_12761;
wire n_14482;
wire n_12113;
wire n_8102;
wire n_14440;
wire n_10541;
wire n_13393;
wire n_14765;
wire n_9793;
wire n_11419;
wire n_14214;
wire n_13202;
wire n_8196;
wire n_11171;
wire n_7112;
wire n_8822;
wire n_5213;
wire n_12017;
wire n_14483;
wire n_5738;
wire n_9514;
wire n_7971;
wire n_12139;
wire n_8885;
wire n_11564;
wire n_5592;
wire n_11078;
wire n_5620;
wire n_12802;
wire n_5491;
wire n_4831;
wire n_10633;
wire n_12592;
wire n_4782;
wire n_9825;
wire n_10573;
wire n_5216;
wire n_11218;
wire n_5953;
wire n_15799;
wire n_8474;
wire n_15315;
wire n_5703;
wire n_10258;
wire n_6886;
wire n_7078;
wire n_4597;
wire n_12791;
wire n_9501;
wire n_12352;
wire n_13811;
wire n_12296;
wire n_11459;
wire n_9043;
wire n_8152;
wire n_12491;
wire n_11998;
wire n_8269;
wire n_4546;
wire n_11775;
wire n_5187;
wire n_7006;
wire n_5119;
wire n_11288;
wire n_4147;
wire n_16066;
wire n_12454;
wire n_10042;
wire n_12162;
wire n_10570;
wire n_13151;
wire n_6531;
wire n_9481;
wire n_11768;
wire n_7577;
wire n_4576;
wire n_12992;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_11456;
wire n_15109;
wire n_14706;
wire n_11708;
wire n_15407;
wire n_14330;
wire n_12960;
wire n_8144;
wire n_5148;
wire n_6726;
wire n_11662;
wire n_6983;
wire n_13617;
wire n_16013;
wire n_7513;
wire n_10098;
wire n_4340;
wire n_15320;
wire n_7812;
wire n_5330;
wire n_9766;
wire n_9351;
wire n_13935;
wire n_13930;
wire n_6935;
wire n_6984;
wire n_6778;
wire n_10106;
wire n_8058;
wire n_11877;
wire n_12046;
wire n_8909;
wire n_6897;
wire n_4284;
wire n_5526;
wire n_5202;
wire n_12074;
wire n_15819;
wire n_14380;
wire n_6345;
wire n_9242;
wire n_10754;
wire n_6386;
wire n_12749;
wire n_6596;
wire n_14630;
wire n_15303;
wire n_5107;
wire n_7165;
wire n_15598;
wire n_9777;
wire n_15302;
wire n_4680;
wire n_5067;
wire n_11932;
wire n_11821;
wire n_12485;
wire n_14464;
wire n_15188;
wire n_15183;
wire n_9522;
wire n_15904;
wire n_15113;
wire n_14560;
wire n_6830;
wire n_9748;
wire n_5987;
wire n_12488;
wire n_14028;
wire n_12252;
wire n_10851;
wire n_9005;
wire n_12090;
wire n_11395;
wire n_10387;
wire n_6642;
wire n_6291;
wire n_9666;
wire n_6510;
wire n_10615;
wire n_5264;
wire n_14081;
wire n_14281;
wire n_10790;
wire n_10028;
wire n_15842;
wire n_10555;
wire n_12896;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_11532;
wire n_8024;
wire n_7123;
wire n_14670;
wire n_4562;
wire n_10222;
wire n_12868;
wire n_15233;
wire n_6509;
wire n_10671;
wire n_8107;
wire n_6376;
wire n_9605;
wire n_10498;
wire n_13959;
wire n_15747;
wire n_9947;
wire n_16033;
wire n_9930;
wire n_14921;
wire n_14755;
wire n_13292;
wire n_4995;
wire n_15250;
wire n_5873;
wire n_6514;
wire n_10420;
wire n_4498;
wire n_6741;
wire n_10083;
wire n_10520;
wire n_14839;
wire n_6434;
wire n_9662;
wire n_5741;
wire n_9768;
wire n_12583;
wire n_6593;
wire n_7827;
wire n_7631;
wire n_15934;
wire n_8748;
wire n_14420;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_10255;
wire n_8742;
wire n_8393;
wire n_9835;
wire n_11117;
wire n_11494;
wire n_9656;
wire n_11643;
wire n_14613;
wire n_12462;
wire n_12618;
wire n_14090;
wire n_14604;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_9475;
wire n_16226;
wire n_14347;
wire n_11475;
wire n_8122;
wire n_11004;
wire n_9724;
wire n_6947;
wire n_8403;
wire n_8912;
wire n_10612;
wire n_4850;
wire n_15613;
wire n_15676;
wire n_10007;
wire n_9154;
wire n_12127;
wire n_13651;
wire n_15773;
wire n_11223;
wire n_11570;
wire n_7157;
wire n_15945;
wire n_10937;
wire n_4937;
wire n_8740;
wire n_10493;
wire n_13631;
wire n_5574;
wire n_13264;
wire n_15012;
wire n_13678;
wire n_8310;
wire n_5877;
wire n_14406;
wire n_10104;
wire n_6375;
wire n_11212;
wire n_10552;
wire n_7781;
wire n_13294;
wire n_4786;
wire n_6042;
wire n_14746;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_10295;
wire n_8296;
wire n_10954;
wire n_7091;
wire n_9833;
wire n_9788;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_9589;
wire n_6315;
wire n_16133;
wire n_7855;
wire n_15314;
wire n_15560;
wire n_14590;
wire n_8850;
wire n_9861;
wire n_15526;
wire n_7886;
wire n_14740;
wire n_7675;
wire n_11122;
wire n_6775;
wire n_8943;
wire n_4345;
wire n_8993;
wire n_11159;
wire n_12329;
wire n_9205;
wire n_15450;
wire n_11631;
wire n_9418;
wire n_9946;
wire n_10376;
wire n_7774;
wire n_8634;
wire n_12611;
wire n_11715;
wire n_13625;
wire n_8831;
wire n_6970;
wire n_13034;
wire n_9979;
wire n_12205;
wire n_13122;
wire n_6948;
wire n_14324;
wire n_14956;
wire n_13210;
wire n_5155;
wire n_8676;
wire n_14337;
wire n_15119;
wire n_11889;
wire n_14509;
wire n_6133;
wire n_6920;
wire n_10087;
wire n_7409;
wire n_10341;
wire n_5408;
wire n_11278;
wire n_12606;
wire n_14692;
wire n_8758;
wire n_11671;
wire n_5812;
wire n_15008;
wire n_9973;
wire n_5540;
wire n_11782;
wire n_7381;
wire n_5804;
wire n_9007;
wire n_8544;
wire n_7999;
wire n_5066;
wire n_14253;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_9020;
wire n_10027;
wire n_9260;
wire n_5130;
wire n_14212;
wire n_4175;
wire n_10154;
wire n_6241;
wire n_13597;
wire n_9619;
wire n_14392;
wire n_13510;
wire n_5200;
wire n_9235;
wire n_14973;
wire n_15822;
wire n_10161;
wire n_13003;
wire n_8652;
wire n_15203;
wire n_9112;
wire n_12365;
wire n_12423;
wire n_7873;
wire n_12843;
wire n_4456;
wire n_11372;
wire n_15219;
wire n_9691;
wire n_5992;
wire n_8646;
wire n_15782;
wire n_13573;
wire n_12518;
wire n_12861;
wire n_9133;
wire n_5684;
wire n_13708;
wire n_7228;
wire n_5981;
wire n_14987;
wire n_7784;
wire n_9752;
wire n_6632;
wire n_8999;
wire n_4948;
wire n_15041;
wire n_10902;
wire n_5413;
wire n_15477;
wire n_7713;
wire n_6623;
wire n_9395;
wire n_5111;
wire n_5150;
wire n_6933;
wire n_15770;
wire n_10294;
wire n_9353;
wire n_11155;
wire n_11714;
wire n_12293;
wire n_13947;
wire n_15908;
wire n_4984;
wire n_5444;
wire n_4410;
wire n_8031;
wire n_11590;
wire n_9804;
wire n_12450;
wire n_5737;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_8439;
wire n_8575;
wire n_5615;
wire n_6908;
wire n_13648;
wire n_5097;
wire n_10323;
wire n_7084;
wire n_11976;
wire n_13274;
wire n_6083;
wire n_6537;
wire n_8499;
wire n_9397;
wire n_10969;
wire n_13015;
wire n_13472;
wire n_13322;
wire n_13870;
wire n_6390;
wire n_7640;
wire n_12000;
wire n_6799;
wire n_8772;
wire n_10806;
wire n_9767;
wire n_12903;
wire n_7912;
wire n_6278;
wire n_11430;
wire n_7195;
wire n_12309;
wire n_15072;
wire n_5640;
wire n_13401;
wire n_13891;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_16007;
wire n_9384;
wire n_4492;
wire n_15284;
wire n_13850;
wire n_15894;
wire n_13835;
wire n_5550;
wire n_15224;
wire n_10666;
wire n_12895;
wire n_5661;
wire n_7641;
wire n_15029;
wire n_4975;
wire n_11638;
wire n_12687;
wire n_12023;
wire n_14460;
wire n_5306;
wire n_5905;
wire n_13908;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_11659;
wire n_9906;
wire n_15942;
wire n_8679;
wire n_5457;
wire n_5159;
wire n_11948;
wire n_15640;
wire n_7115;
wire n_16216;
wire n_9310;
wire n_11843;
wire n_15382;
wire n_16196;
wire n_10659;
wire n_11689;
wire n_7764;
wire n_8446;
wire n_9163;
wire n_11535;
wire n_12022;
wire n_12624;
wire n_4336;
wire n_11808;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_9322;
wire n_12719;
wire n_7616;
wire n_14493;
wire n_10793;
wire n_14868;
wire n_14491;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_6412;
wire n_15495;
wire n_6271;
wire n_11108;
wire n_9377;
wire n_7235;
wire n_6572;
wire n_9224;
wire n_10211;
wire n_10837;
wire n_14381;
wire n_12664;
wire n_13020;
wire n_11577;
wire n_15045;
wire n_7271;
wire n_9055;
wire n_15686;
wire n_13749;
wire n_13311;
wire n_7222;
wire n_8678;
wire n_9971;
wire n_8605;
wire n_12981;
wire n_13945;
wire n_10976;
wire n_9624;
wire n_14766;
wire n_6930;
wire n_10045;
wire n_15026;
wire n_14172;
wire n_10289;
wire n_5482;
wire n_9145;
wire n_12716;
wire n_10232;
wire n_13079;
wire n_11098;
wire n_15177;
wire n_15130;
wire n_8443;
wire n_8525;
wire n_12166;
wire n_12507;
wire n_8312;
wire n_10819;
wire n_16035;
wire n_15968;
wire n_8901;
wire n_13786;
wire n_13645;
wire n_6584;
wire n_4494;
wire n_9887;
wire n_12044;
wire n_6387;
wire n_9373;
wire n_4201;
wire n_15359;
wire n_14374;
wire n_6470;
wire n_7206;
wire n_16019;
wire n_8869;
wire n_11279;
wire n_11729;
wire n_14012;
wire n_9770;
wire n_11514;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_15440;
wire n_5651;
wire n_15587;
wire n_15401;
wire n_6625;
wire n_14569;
wire n_7383;
wire n_12430;
wire n_4636;
wire n_11606;
wire n_4983;
wire n_6826;
wire n_10306;
wire n_12902;
wire n_14664;
wire n_12257;
wire n_11727;
wire n_13299;
wire n_10103;
wire n_11337;
wire n_6341;
wire n_4386;
wire n_6374;
wire n_10183;
wire n_12839;
wire n_13693;
wire n_5623;
wire n_16255;
wire n_11778;
wire n_12925;
wire n_11658;
wire n_10710;
wire n_8870;
wire n_9753;
wire n_5041;
wire n_4275;
wire n_5023;
wire n_10931;
wire n_9468;
wire n_11433;
wire n_8178;
wire n_7854;
wire n_5524;
wire n_9517;
wire n_15821;
wire n_16179;
wire n_9544;
wire n_7959;
wire n_5735;
wire n_14338;
wire n_14728;
wire n_15009;
wire n_8234;
wire n_6363;
wire n_13434;
wire n_6588;
wire n_11369;
wire n_14865;
wire n_15642;
wire n_4243;
wire n_12759;
wire n_7897;
wire n_11720;
wire n_14418;
wire n_15197;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_13500;
wire n_14815;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_8488;
wire n_11840;
wire n_6865;
wire n_11284;
wire n_12553;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_9774;
wire n_16194;
wire n_7132;
wire n_11987;
wire n_12016;
wire n_12496;
wire n_11052;
wire n_7533;
wire n_9586;
wire n_10670;
wire n_13655;
wire n_10150;
wire n_16042;
wire n_6722;
wire n_9780;
wire n_13476;
wire n_11177;
wire n_6420;
wire n_14900;
wire n_14803;
wire n_10004;
wire n_4907;
wire n_11169;
wire n_5153;
wire n_7766;
wire n_8862;
wire n_13229;
wire n_14092;
wire n_8184;
wire n_13950;
wire n_5787;
wire n_4713;
wire n_6911;
wire n_11221;
wire n_14219;
wire n_13344;
wire n_10353;
wire n_10151;
wire n_16111;
wire n_11095;
wire n_10187;
wire n_10171;
wire n_11211;
wire n_7129;
wire n_12138;
wire n_7080;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_10406;
wire n_8695;
wire n_12230;
wire n_12521;
wire n_11236;
wire n_11931;
wire n_7436;
wire n_8767;
wire n_11036;
wire n_12562;
wire n_8571;
wire n_7020;
wire n_11600;
wire n_15517;
wire n_5935;
wire n_8064;
wire n_14117;
wire n_15925;
wire n_14588;
wire n_6696;
wire n_13721;
wire n_4916;
wire n_8472;
wire n_10796;
wire n_13302;
wire n_5967;
wire n_15334;
wire n_15295;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_6045;
wire n_5376;
wire n_12217;
wire n_13535;
wire n_14261;
wire n_15581;
wire n_6300;
wire n_13704;
wire n_6653;
wire n_6372;
wire n_13969;
wire n_4129;
wire n_14016;
wire n_7120;
wire n_11114;
wire n_10479;
wire n_7978;
wire n_10033;
wire n_5488;
wire n_9099;
wire n_6900;
wire n_10034;
wire n_5727;
wire n_11336;
wire n_15344;
wire n_15137;
wire n_6660;
wire n_8787;
wire n_11009;
wire n_9543;
wire n_8131;
wire n_5988;
wire n_16248;
wire n_6424;
wire n_10696;
wire n_14633;
wire n_16264;
wire n_11480;
wire n_5646;
wire n_14538;
wire n_7448;
wire n_16209;
wire n_4480;
wire n_5711;
wire n_7694;
wire n_6787;
wire n_8771;
wire n_9245;
wire n_15142;
wire n_5832;
wire n_15418;
wire n_13269;
wire n_6254;
wire n_7460;
wire n_7142;
wire n_10360;
wire n_6423;
wire n_16230;
wire n_6526;
wire n_8150;
wire n_5891;
wire n_14891;
wire n_9168;
wire n_11423;
wire n_16136;
wire n_12691;
wire n_5328;
wire n_9074;
wire n_12159;
wire n_5016;
wire n_6011;
wire n_4616;
wire n_11665;
wire n_12259;
wire n_12975;
wire n_9367;
wire n_9330;
wire n_7465;
wire n_11556;
wire n_11685;
wire n_13402;
wire n_14231;
wire n_15662;
wire n_5470;
wire n_10230;
wire n_11801;
wire n_12117;
wire n_8917;
wire n_12587;
wire n_15995;
wire n_11573;
wire n_4374;
wire n_6176;
wire n_9300;
wire n_16011;
wire n_14489;
wire n_13619;
wire n_14663;
wire n_11589;
wire n_14395;
wire n_11667;
wire n_8230;
wire n_10414;
wire n_6222;
wire n_13110;
wire n_12422;
wire n_8352;
wire n_7760;
wire n_15042;
wire n_9918;
wire n_12977;
wire n_6969;
wire n_13060;
wire n_15651;
wire n_9496;
wire n_13177;
wire n_15214;
wire n_8914;
wire n_10953;
wire n_14082;
wire n_8821;
wire n_11446;
wire n_13853;
wire n_8465;
wire n_15285;
wire n_6587;
wire n_6688;
wire n_8360;
wire n_6505;
wire n_13586;
wire n_15163;
wire n_9837;
wire n_12772;
wire n_15979;
wire n_5362;
wire n_8209;
wire n_15421;
wire n_8986;
wire n_14701;
wire n_4580;
wire n_15867;
wire n_6762;
wire n_15191;
wire n_11633;
wire n_5147;
wire n_15697;
wire n_4826;
wire n_11011;
wire n_4514;
wire n_7629;
wire n_12145;
wire n_10787;
wire n_6987;
wire n_7567;
wire n_8743;
wire n_11342;
wire n_8963;
wire n_9191;
wire n_11812;
wire n_6453;
wire n_9114;
wire n_6308;
wire n_11142;
wire n_13074;
wire n_10896;
wire n_8396;
wire n_13773;
wire n_15582;
wire n_8514;
wire n_12196;
wire n_16177;
wire n_13482;
wire n_8550;
wire n_7449;
wire n_11959;
wire n_8151;
wire n_13927;
wire n_14688;
wire n_16242;
wire n_15579;
wire n_12889;
wire n_15793;
wire n_13096;
wire n_12493;
wire n_9913;
wire n_6187;
wire n_15436;
wire n_11626;
wire n_6597;
wire n_13810;
wire n_11178;
wire n_12440;
wire n_4844;
wire n_9329;
wire n_6220;
wire n_13684;
wire n_14452;
wire n_12608;
wire n_15439;
wire n_13800;
wire n_10598;
wire n_13008;
wire n_7479;
wire n_7882;
wire n_13607;
wire n_11750;
wire n_13742;
wire n_7517;
wire n_16002;
wire n_9627;
wire n_13412;
wire n_11283;
wire n_10271;
wire n_11338;
wire n_5037;
wire n_11295;
wire n_15668;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_5189;
wire n_4677;
wire n_8070;
wire n_15342;
wire n_14896;
wire n_4525;
wire n_8866;
wire n_10402;
wire n_6149;
wire n_11191;
wire n_15595;
wire n_10064;
wire n_11661;
wire n_13329;
wire n_10137;
wire n_9585;
wire n_14863;
wire n_5055;
wire n_7878;
wire n_9376;
wire n_4369;
wire n_12515;
wire n_15232;
wire n_16135;
wire n_5648;
wire n_12249;
wire n_11644;
wire n_15742;
wire n_6439;
wire n_4324;
wire n_11354;
wire n_15298;
wire n_13537;
wire n_8797;
wire n_14247;
wire n_14462;
wire n_6547;
wire n_13075;
wire n_11126;
wire n_9524;
wire n_7177;
wire n_7902;
wire n_11408;
wire n_12623;
wire n_5160;
wire n_12971;
wire n_13051;
wire n_15206;
wire n_12674;
wire n_15193;
wire n_5762;
wire n_9606;
wire n_15768;
wire n_14419;
wire n_10800;
wire n_5484;
wire n_12026;
wire n_13038;
wire n_14514;
wire n_13812;
wire n_14733;
wire n_10019;
wire n_10762;
wire n_14135;
wire n_7353;
wire n_11935;
wire n_8054;
wire n_10047;
wire n_6478;
wire n_16221;
wire n_11037;
wire n_4989;
wire n_5874;
wire n_13977;
wire n_8841;
wire n_11396;
wire n_9084;
wire n_14681;
wire n_7050;
wire n_7590;
wire n_14453;
wire n_6906;
wire n_6739;
wire n_15657;
wire n_15720;
wire n_10995;
wire n_4898;
wire n_14869;
wire n_4528;
wire n_14036;
wire n_15490;
wire n_10597;
wire n_10561;
wire n_14994;
wire n_7818;
wire n_12345;
wire n_7645;
wire n_15655;
wire n_7482;
wire n_5385;
wire n_13841;
wire n_14312;
wire n_11726;
wire n_12346;
wire n_5622;
wire n_14522;
wire n_14110;
wire n_15647;
wire n_10523;
wire n_8618;
wire n_10377;
wire n_10243;
wire n_5635;
wire n_8538;
wire n_8590;
wire n_13883;
wire n_14945;
wire n_7907;
wire n_9204;
wire n_8970;
wire n_4280;
wire n_6034;
wire n_5609;
wire n_15558;
wire n_8791;
wire n_15013;
wire n_14739;
wire n_13724;
wire n_4811;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_10165;
wire n_14776;
wire n_9616;
wire n_5380;
wire n_9708;
wire n_7862;
wire n_10153;
wire n_9130;
wire n_9988;
wire n_8703;
wire n_12265;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_12147;
wire n_7721;
wire n_4524;
wire n_9209;
wire n_15374;
wire n_8061;
wire n_10775;
wire n_10173;
wire n_10585;
wire n_4657;
wire n_5568;
wire n_12075;
wire n_8754;
wire n_15755;
wire n_14996;
wire n_8864;
wire n_5941;
wire n_15478;
wire n_10985;
wire n_4891;
wire n_11300;
wire n_14294;
wire n_8837;
wire n_12108;
wire n_10999;
wire n_13425;
wire n_13791;
wire n_8915;
wire n_15251;
wire n_10587;
wire n_8784;
wire n_11219;
wire n_6604;
wire n_6611;
wire n_5364;
wire n_15833;
wire n_15415;
wire n_11857;
wire n_5597;
wire n_11735;
wire n_11986;
wire n_9086;
wire n_8768;
wire n_12102;
wire n_6999;
wire n_8072;
wire n_8086;
wire n_9014;
wire n_15205;
wire n_5469;
wire n_6019;
wire n_7539;
wire n_14611;
wire n_9010;
wire n_11637;
wire n_13925;
wire n_16100;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_14417;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_11072;
wire n_12183;
wire n_13432;
wire n_15860;
wire n_4876;
wire n_16022;
wire n_15084;
wire n_16193;
wire n_15217;
wire n_5021;
wire n_12519;
wire n_12955;
wire n_9044;
wire n_13538;
wire n_14176;
wire n_5936;
wire n_14650;
wire n_8307;
wire n_14939;
wire n_14789;
wire n_13774;
wire n_5312;
wire n_15290;
wire n_6784;
wire n_9694;
wire n_16237;
wire n_11421;
wire n_13323;
wire n_10718;
wire n_13214;
wire n_10951;
wire n_10412;
wire n_8470;
wire n_15216;
wire n_5928;
wire n_7830;
wire n_8050;
wire n_14980;
wire n_10310;
wire n_4200;
wire n_5785;
wire n_5222;
wire n_10655;
wire n_9633;
wire n_6165;
wire n_10133;
wire n_12793;
wire n_11989;
wire n_15399;
wire n_10942;
wire n_4938;
wire n_6114;
wire n_13192;
wire n_15189;
wire n_13392;
wire n_13433;
wire n_5505;
wire n_14662;
wire n_12865;
wire n_4604;
wire n_9261;
wire n_11331;
wire n_12285;
wire n_5504;
wire n_7348;
wire n_9345;
wire n_14894;
wire n_11953;
wire n_6829;
wire n_11820;
wire n_12478;
wire n_9375;
wire n_4239;
wire n_9472;
wire n_9764;
wire n_10509;
wire n_8010;
wire n_13059;
wire n_12522;
wire n_13451;
wire n_9448;
wire n_6464;
wire n_8802;
wire n_8950;
wire n_5129;
wire n_13199;
wire n_7320;
wire n_4704;
wire n_9487;
wire n_8603;
wire n_15654;
wire n_15691;
wire n_10639;
wire n_13588;
wire n_5494;
wire n_5970;
wire n_15531;
wire n_11358;
wire n_12413;
wire n_6838;
wire n_13191;
wire n_16102;
wire n_6368;
wire n_14133;
wire n_10690;
wire n_12369;
wire n_12681;
wire n_7935;
wire n_11118;
wire n_8143;
wire n_11844;
wire n_9271;
wire n_5663;
wire n_15332;
wire n_12084;
wire n_5161;
wire n_14132;
wire n_7933;
wire n_12152;
wire n_12726;
wire n_12784;
wire n_7155;
wire n_6640;
wire n_9851;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_15281;
wire n_5626;
wire n_4706;
wire n_6850;
wire n_12511;
wire n_4343;
wire n_12520;
wire n_12705;
wire n_7743;
wire n_4764;
wire n_5389;
wire n_11861;
wire n_13899;
wire n_14443;
wire n_4990;
wire n_8584;
wire n_14934;
wire n_11370;
wire n_13017;
wire n_9101;
wire n_15186;
wire n_16266;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_15461;
wire n_8574;
wire n_12832;
wire n_4919;
wire n_15145;
wire n_13422;
wire n_15448;
wire n_15834;
wire n_7043;
wire n_7986;
wire n_8049;
wire n_9927;
wire n_12207;
wire n_13666;
wire n_12782;
wire n_7266;
wire n_13042;
wire n_15875;
wire n_10621;
wire n_11884;
wire n_5653;
wire n_15664;
wire n_14860;
wire n_4835;
wire n_4420;
wire n_15299;
wire n_7996;
wire n_14513;
wire n_12970;
wire n_15507;
wire n_10789;
wire n_4251;
wire n_5266;
wire n_10496;
wire n_12384;
wire n_4559;
wire n_4742;
wire n_12605;
wire n_5038;
wire n_14724;
wire n_15011;
wire n_15679;
wire n_10319;
wire n_15683;
wire n_15871;
wire n_5800;
wire n_14021;
wire n_8509;
wire n_14830;
wire n_12408;
wire n_16223;
wire n_4372;
wire n_5396;
wire n_9850;
wire n_4162;
wire n_5766;
wire n_10499;
wire n_14223;
wire n_11717;
wire n_5293;
wire n_10224;
wire n_13234;
wire n_15155;
wire n_4790;
wire n_7035;
wire n_10970;
wire n_4173;
wire n_8354;
wire n_12651;
wire n_5309;
wire n_15501;
wire n_15059;
wire n_6047;
wire n_9432;
wire n_12160;
wire n_13829;
wire n_11464;
wire n_16263;
wire n_11243;
wire n_9824;
wire n_14582;
wire n_8277;
wire n_10827;
wire n_7442;
wire n_4727;
wire n_14880;
wire n_6568;
wire n_11473;
wire n_14508;
wire n_5627;
wire n_10055;
wire n_12638;
wire n_12698;
wire n_11654;
wire n_13878;
wire n_10783;
wire n_15208;
wire n_14562;
wire n_8583;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_8644;
wire n_10148;
wire n_7939;
wire n_9884;
wire n_7715;
wire n_11534;
wire n_10465;
wire n_14040;
wire n_14361;
wire n_11749;
wire n_7350;
wire n_15972;
wire n_7314;
wire n_6026;
wire n_10610;
wire n_8609;
wire n_13955;
wire n_9144;
wire n_15453;
wire n_8052;
wire n_12481;
wire n_4799;
wire n_8733;
wire n_9758;
wire n_12078;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_12815;
wire n_4534;
wire n_12129;
wire n_5636;
wire n_4960;
wire n_9931;
wire n_7699;
wire n_9693;
wire n_11546;
wire n_12502;
wire n_10830;
wire n_9273;
wire n_15530;
wire n_16126;
wire n_9196;
wire n_5707;
wire n_15474;
wire n_5594;
wire n_9029;
wire n_10086;
wire n_15614;
wire n_5697;
wire n_13763;
wire n_7580;
wire n_5606;
wire n_15737;
wire n_11785;
wire n_6727;
wire n_5911;
wire n_12697;
wire n_7340;
wire n_8080;
wire n_13437;
wire n_10279;
wire n_7303;
wire n_10932;
wire n_11440;
wire n_9967;
wire n_15849;
wire n_12908;
wire n_16078;
wire n_8819;
wire n_7870;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_14799;
wire n_7387;
wire n_8487;
wire n_13293;
wire n_6454;
wire n_11697;
wire n_11545;
wire n_16183;
wire n_13487;
wire n_13555;
wire n_15591;
wire n_13239;
wire n_10487;
wire n_14579;
wire n_14853;
wire n_9881;
wire n_11645;
wire n_12512;
wire n_11263;
wire n_12199;
wire n_15043;
wire n_6333;
wire n_11937;
wire n_7004;
wire n_15538;
wire n_12584;
wire n_13854;
wire n_13361;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_10910;
wire n_5058;
wire n_8382;
wire n_9733;
wire n_16139;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_13558;
wire n_9075;
wire n_11324;
wire n_13954;
wire n_4166;
wire n_5356;
wire n_11763;
wire n_13803;
wire n_7167;
wire n_5849;
wire n_11853;
wire n_12988;
wire n_14537;
wire n_8906;
wire n_5841;
wire n_10109;
wire n_7146;
wire n_7030;
wire n_14542;
wire n_10857;
wire n_4478;
wire n_8203;
wire n_9442;
wire n_15096;
wire n_4246;
wire n_7618;
wire n_14625;
wire n_13244;
wire n_4632;
wire n_13305;
wire n_15741;
wire n_12284;
wire n_11364;
wire n_11941;
wire n_9630;
wire n_11359;
wire n_12031;
wire n_14203;
wire n_9898;
wire n_15926;
wire n_11323;
wire n_11504;
wire n_15146;
wire n_11704;
wire n_11587;
wire n_13697;
wire n_11620;
wire n_12652;
wire n_8340;
wire n_4754;
wire n_9582;
wire n_8268;
wire n_10865;
wire n_15291;
wire n_16029;
wire n_8171;
wire n_4375;
wire n_12850;
wire n_15244;
wire n_9877;
wire n_14578;
wire n_10179;
wire n_12969;
wire n_12379;
wire n_10925;
wire n_12607;
wire n_13743;
wire n_9986;
wire n_13951;
wire n_14222;
wire n_13695;
wire n_8008;
wire n_7633;
wire n_10246;
wire n_9636;
wire n_4684;
wire n_10439;
wire n_13376;
wire n_14377;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_8824;
wire n_11902;
wire n_7280;
wire n_8369;
wire n_5043;
wire n_12701;
wire n_14008;
wire n_7339;
wire n_7597;
wire n_8884;
wire n_12898;
wire n_4241;
wire n_9225;
wire n_4183;
wire n_7768;
wire n_11282;
wire n_5645;
wire n_5020;
wire n_6455;
wire n_13639;
wire n_7615;
wire n_16015;
wire n_12475;
wire n_16208;
wire n_10182;
wire n_14795;
wire n_8271;
wire n_9091;
wire n_6183;
wire n_13772;
wire n_14643;
wire n_12027;
wire n_8392;
wire n_15835;
wire n_8309;
wire n_14986;
wire n_6107;
wire n_15685;
wire n_12218;
wire n_10795;
wire n_13602;
wire n_6476;
wire n_5232;
wire n_16197;
wire n_10046;
wire n_4256;
wire n_9412;
wire n_11834;
wire n_8874;
wire n_8228;
wire n_12174;
wire n_5035;
wire n_11405;
wire n_11028;
wire n_11663;
wire n_5453;
wire n_4333;
wire n_15645;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_15646;
wire n_12385;
wire n_14407;
wire n_15321;
wire n_15882;
wire n_6636;
wire n_9525;
wire n_11071;
wire n_12289;
wire n_11625;
wire n_15626;
wire n_11187;
wire n_12041;
wire n_12565;
wire n_12882;
wire n_13736;
wire n_15075;
wire n_13254;
wire n_12819;
wire n_8172;
wire n_14810;
wire n_4455;
wire n_13341;
wire n_6554;
wire n_9575;
wire n_5631;
wire n_6994;
wire n_7401;
wire n_10413;
wire n_10456;
wire n_11566;
wire n_11271;
wire n_12164;
wire n_12433;
wire n_15383;
wire n_11649;
wire n_12224;
wire n_13061;
wire n_5101;
wire n_9738;
wire n_10735;
wire n_6020;
wire n_13328;
wire n_14908;
wire n_9252;
wire n_16259;
wire n_12550;
wire n_6185;
wire n_8344;
wire n_12800;
wire n_14568;
wire n_15452;
wire n_16012;
wire n_14259;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_12561;
wire n_8936;
wire n_8738;
wire n_10822;
wire n_9739;
wire n_6785;
wire n_14871;
wire n_9727;
wire n_10508;
wire n_4735;
wire n_6870;
wire n_6643;
wire n_13281;
wire n_15323;
wire n_7574;
wire n_5170;
wire n_8226;
wire n_15272;
wire n_14874;
wire n_6695;
wire n_7529;
wire n_5608;
wire n_6501;
wire n_11308;
wire n_11739;
wire n_11593;
wire n_9148;
wire n_10858;
wire n_6466;
wire n_10736;
wire n_11828;
wire n_9958;
wire n_6467;
wire n_14138;
wire n_9323;
wire n_4212;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_9779;
wire n_15074;
wire n_8088;
wire n_5702;
wire n_14244;
wire n_9545;
wire n_8930;
wire n_9155;
wire n_12563;
wire n_8662;
wire n_13114;
wire n_11291;
wire n_11425;
wire n_13566;
wire n_9046;
wire n_9430;
wire n_11890;
wire n_4477;
wire n_5806;
wire n_9625;
wire n_13621;
wire n_8783;
wire n_12398;
wire n_13624;
wire n_5182;
wire n_4217;
wire n_8663;
wire n_14015;
wire n_10928;
wire n_5277;
wire n_6507;
wire n_10842;
wire n_12941;
wire n_6618;
wire n_9447;
wire n_13407;
wire n_15865;
wire n_13404;
wire n_16195;
wire n_6213;
wire n_8364;
wire n_9485;
wire n_4949;
wire n_15857;
wire n_14818;
wire n_8490;
wire n_8981;
wire n_9129;
wire n_12461;
wire n_11832;
wire n_7872;
wire n_6873;
wire n_7958;
wire n_4605;
wire n_8118;
wire n_4649;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_12095;
wire n_15714;
wire n_14191;
wire n_8785;
wire n_11470;
wire n_11744;
wire n_10210;
wire n_11294;
wire n_13994;
wire n_14841;
wire n_15817;
wire n_7843;
wire n_12998;
wire n_9047;
wire n_13219;
wire n_15952;
wire n_10057;
wire n_6063;
wire n_13737;
wire n_16245;
wire n_12630;
wire n_11641;
wire n_15141;
wire n_15464;
wire n_15181;
wire n_7578;
wire n_12789;
wire n_12679;
wire n_14146;
wire n_13372;
wire n_5415;
wire n_14084;
wire n_7261;
wire n_8982;
wire n_10739;
wire n_4592;
wire n_4999;
wire n_12327;
wire n_6993;
wire n_9745;
wire n_14288;
wire n_12038;
wire n_13932;
wire n_10533;
wire n_4820;
wire n_13978;
wire n_11875;
wire n_8100;
wire n_10878;
wire n_15600;
wire n_10988;
wire n_8522;
wire n_13563;
wire n_15733;
wire n_13141;
wire n_12338;
wire n_10993;
wire n_13249;
wire n_8381;
wire n_9320;
wire n_8835;
wire n_6767;
wire n_11014;
wire n_4656;
wire n_4862;
wire n_12030;
wire n_14553;
wire n_15258;
wire n_5687;
wire n_6558;
wire n_13517;
wire n_6755;
wire n_9108;
wire n_9457;
wire n_15001;
wire n_9907;
wire n_10959;
wire n_6153;
wire n_15545;
wire n_11310;
wire n_7263;
wire n_11062;
wire n_10940;
wire n_12067;
wire n_13783;
wire n_12675;
wire n_6608;
wire n_11400;
wire n_11040;
wire n_15797;
wire n_6202;
wire n_15353;
wire n_6780;
wire n_7688;
wire n_13968;
wire n_16073;
wire n_12870;
wire n_14038;
wire n_12291;
wire n_5383;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_9567;
wire n_6359;
wire n_11773;
wire n_14385;
wire n_5690;
wire n_10583;
wire n_14027;
wire n_11332;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_7585;
wire n_8356;
wire n_16146;
wire n_5029;
wire n_13279;
wire n_13731;
wire n_12013;
wire n_13007;
wire n_15818;
wire n_9852;
wire n_10881;
wire n_16037;
wire n_12395;
wire n_16268;
wire n_7418;
wire n_16192;
wire n_6353;
wire n_14049;
wire n_13160;
wire n_11943;
wire n_5218;
wire n_10544;
wire n_12933;
wire n_16271;
wire n_6577;
wire n_7772;
wire n_13895;
wire n_14403;
wire n_13213;
wire n_8736;
wire n_15899;
wire n_12131;
wire n_10491;
wire n_13507;
wire n_6082;
wire n_15625;
wire n_11144;
wire n_13385;
wire n_10926;
wire n_11841;
wire n_8918;
wire n_11766;
wire n_12766;
wire n_10839;
wire n_10603;
wire n_5361;
wire n_7312;
wire n_9022;
wire n_13790;
wire n_7514;
wire n_15985;
wire n_12399;
wire n_8616;
wire n_6105;
wire n_12762;
wire n_10400;
wire n_11518;
wire n_5512;
wire n_13567;
wire n_7738;
wire n_14346;
wire n_14787;
wire n_8838;
wire n_8908;
wire n_13687;
wire n_11960;
wire n_7609;
wire n_13580;
wire n_9161;
wire n_12241;
wire n_10792;
wire n_5898;
wire n_7113;
wire n_15336;
wire n_11274;
wire n_6548;
wire n_8607;
wire n_13779;
wire n_15473;
wire n_16124;
wire n_8213;
wire n_14487;
wire n_13722;
wire n_13225;
wire n_14615;
wire n_15699;
wire n_5923;
wire n_6657;
wire n_10994;
wire n_5617;
wire n_5946;
wire n_13514;
wire n_13806;
wire n_9903;
wire n_9831;
wire n_14595;
wire n_15460;
wire n_10032;
wire n_8436;
wire n_7282;
wire n_13261;
wire n_8551;
wire n_14638;
wire n_13039;
wire n_15524;
wire n_4550;
wire n_14717;
wire n_9238;
wire n_12137;
wire n_14167;
wire n_4347;
wire n_11624;
wire n_10580;
wire n_7921;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_10512;
wire n_9248;
wire n_12495;
wire n_5514;
wire n_11917;
wire n_5611;
wire n_12790;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_4895;
wire n_14924;
wire n_15288;
wire n_9867;
wire n_12106;
wire n_11130;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_10005;
wire n_11053;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_11872;
wire n_5188;
wire n_12434;
wire n_6674;
wire n_15881;
wire n_13669;
wire n_5049;
wire n_12710;
wire n_7489;
wire n_9056;
wire n_6331;
wire n_5308;
wire n_9106;
wire n_4434;
wire n_13303;
wire n_5068;
wire n_12881;
wire n_7863;
wire n_15906;
wire n_6493;
wire n_7363;
wire n_14496;
wire n_7281;
wire n_5739;
wire n_10596;
wire n_12920;
wire n_4199;
wire n_14260;
wire n_7968;
wire n_11220;
wire n_10061;
wire n_10507;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_7833;
wire n_12086;
wire n_11887;
wire n_14189;
wire n_12281;
wire n_15437;
wire n_12991;
wire n_4510;
wire n_14552;
wire n_7750;
wire n_5057;
wire n_9071;
wire n_6196;
wire n_12995;
wire n_16247;
wire n_5425;
wire n_5273;
wire n_10136;
wire n_5839;
wire n_7588;
wire n_10967;
wire n_11551;
wire n_14339;
wire n_13368;
wire n_10369;
wire n_14971;
wire n_7697;
wire n_10025;
wire n_10708;
wire n_11703;
wire n_5887;
wire n_16053;
wire n_13948;
wire n_7808;
wire n_9519;
wire n_15960;
wire n_9027;
wire n_7603;
wire n_13598;
wire n_6321;
wire n_14180;
wire n_5683;
wire n_8704;
wire n_14341;
wire n_8984;
wire n_9786;
wire n_10194;
wire n_7192;
wire n_12807;
wire n_5248;
wire n_4899;
wire n_11153;
wire n_10833;
wire n_10685;
wire n_10513;
wire n_4156;
wire n_8613;
wire n_13611;
wire n_11030;
wire n_14704;
wire n_13178;
wire n_14293;
wire n_10223;
wire n_5880;
wire n_13495;
wire n_15417;
wire n_8012;
wire n_12012;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_16016;
wire n_9404;
wire n_13777;
wire n_5666;
wire n_13301;
wire n_11368;
wire n_12098;
wire n_7988;
wire n_12025;
wire n_12669;
wire n_15468;
wire n_13205;
wire n_15617;
wire n_4448;
wire n_10410;
wire n_13049;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_9370;
wire n_15553;
wire n_6995;
wire n_13009;
wire n_16175;
wire n_4193;
wire n_4579;
wire n_6347;
wire n_14885;
wire n_13748;
wire n_14878;
wire n_13338;
wire n_6496;
wire n_13747;
wire n_4776;
wire n_8387;
wire n_9352;
wire n_14972;
wire n_11716;
wire n_14083;
wire n_8105;
wire n_10984;
wire n_13485;
wire n_10144;
wire n_16167;
wire n_12019;
wire n_6745;
wire n_7943;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_13416;
wire n_12255;
wire n_7377;
wire n_11967;
wire n_8900;
wire n_4392;
wire n_6064;
wire n_9681;
wire n_14439;
wire n_8353;
wire n_12503;
wire n_9051;
wire n_7723;
wire n_4691;
wire n_7904;
wire n_5682;
wire n_5461;
wire n_9098;
wire n_12415;
wire n_7296;
wire n_4397;
wire n_8323;
wire n_13053;
wire n_13752;
wire n_10459;
wire n_12951;
wire n_14125;
wire n_6164;
wire n_11426;
wire n_8711;
wire n_13273;
wire n_15787;
wire n_11628;
wire n_4753;
wire n_12704;
wire n_9484;
wire n_4803;
wire n_8731;
wire n_5730;
wire n_10155;
wire n_11367;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_16020;
wire n_5754;
wire n_11418;
wire n_8597;
wire n_6330;
wire n_15289;
wire n_7178;
wire n_11026;
wire n_15672;
wire n_7045;
wire n_11576;
wire n_9853;
wire n_8534;
wire n_15046;
wire n_8655;
wire n_9210;
wire n_12884;
wire n_16056;
wire n_16165;
wire n_13324;
wire n_4893;
wire n_10915;
wire n_13414;
wire n_13894;
wire n_10949;
wire n_7777;
wire n_12339;
wire n_8302;
wire n_14616;
wire n_4258;
wire n_5756;
wire n_14784;
wire n_14695;
wire n_14455;
wire n_12911;
wire n_15301;
wire n_8496;
wire n_7693;
wire n_11150;
wire n_10156;
wire n_5033;
wire n_11123;
wire n_14414;
wire n_10248;
wire n_14941;
wire n_6015;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_14449;
wire n_16273;
wire n_11733;
wire n_15903;
wire n_10215;
wire n_10624;
wire n_12915;
wire n_7682;
wire n_7300;
wire n_6861;
wire n_10152;
wire n_12888;
wire n_15811;
wire n_4203;
wire n_12105;
wire n_9756;
wire n_16132;
wire n_5789;
wire n_12034;
wire n_5400;
wire n_7558;
wire n_5347;
wire n_14744;
wire n_11188;
wire n_9166;
wire n_8103;
wire n_8719;
wire n_10877;
wire n_15954;
wire n_7798;
wire n_9778;
wire n_8879;
wire n_13906;
wire n_4767;
wire n_15218;
wire n_8969;
wire n_9141;
wire n_4569;
wire n_11209;
wire n_6528;
wire n_14441;
wire n_13159;
wire n_9700;
wire n_10316;
wire n_8896;
wire n_5144;
wire n_11503;
wire n_14769;
wire n_6895;
wire n_10385;
wire n_15192;
wire n_15775;
wire n_14732;
wire n_8335;
wire n_13337;
wire n_4468;
wire n_5509;
wire n_15917;
wire n_15433;
wire n_7400;
wire n_14230;
wire n_11699;
wire n_13145;
wire n_16014;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_12549;
wire n_6523;
wire n_11817;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_14618;
wire n_11469;
wire n_9363;
wire n_11971;
wire n_4698;
wire n_14199;
wire n_16003;
wire n_15497;
wire n_14722;
wire n_5349;
wire n_14101;
wire n_6472;
wire n_9532;
wire n_10823;
wire n_12237;
wire n_14001;
wire n_6389;
wire n_14623;
wire n_14586;
wire n_14635;
wire n_15586;
wire n_10680;
wire n_5534;
wire n_9307;
wire n_13922;
wire n_9876;
wire n_12220;
wire n_12564;
wire n_10814;
wire n_12375;
wire n_13333;
wire n_5183;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_9959;
wire n_8834;
wire n_9989;
wire n_10651;
wire n_14495;
wire n_8286;
wire n_8417;
wire n_13872;
wire n_12809;
wire n_8964;
wire n_10611;
wire n_6869;
wire n_4761;
wire n_4627;
wire n_10549;
wire n_10370;
wire n_11621;
wire n_7672;
wire n_10770;
wire n_14171;
wire n_4556;
wire n_6137;
wire n_9467;
wire n_15635;
wire n_11558;
wire n_12043;
wire n_12513;
wire n_14988;
wire n_5254;
wire n_12337;
wire n_10393;
wire n_5079;
wire n_14975;
wire n_8247;
wire n_9406;
wire n_10089;
wire n_11417;
wire n_11113;
wire n_14182;
wire n_4520;
wire n_10543;
wire n_13355;
wire n_15639;
wire n_8639;
wire n_12504;
wire n_15246;
wire n_11301;
wire n_9160;
wire n_5751;
wire n_11051;
wire n_12489;
wire n_10321;
wire n_12886;
wire n_13308;
wire n_7712;
wire n_4444;
wire n_4263;
wire n_7681;
wire n_6885;
wire n_15173;
wire n_5039;
wire n_6613;
wire n_6580;
wire n_8566;
wire n_8727;
wire n_15492;
wire n_14791;
wire n_4265;
wire n_8482;
wire n_6404;
wire n_6120;
wire n_13905;
wire n_11018;
wire n_13923;
wire n_14884;
wire n_15956;
wire n_10259;
wire n_14927;
wire n_7491;
wire n_15194;
wire n_12836;
wire n_14243;
wire n_13936;
wire n_15419;
wire n_10909;
wire n_10094;
wire n_8599;
wire n_4612;
wire n_14386;
wire n_5997;
wire n_10302;
wire n_11328;
wire n_15243;
wire n_8781;
wire n_5375;
wire n_5438;
wire n_9167;
wire n_11276;
wire n_15796;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_6530;
wire n_6602;
wire n_15845;
wire n_7915;
wire n_4149;
wire n_4958;
wire n_6135;
wire n_12655;
wire n_10623;
wire n_8839;
wire n_11326;
wire n_13627;
wire n_14359;
wire n_14786;
wire n_4538;
wire n_5563;
wire n_13882;
wire n_12779;
wire n_8365;
wire n_15973;
wire n_13144;
wire n_14085;
wire n_6942;
wire n_7860;
wire n_14108;
wire n_6892;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8489;
wire n_13364;
wire n_8859;
wire n_8060;
wire n_9290;
wire n_6782;
wire n_6230;
wire n_4421;
wire n_15319;
wire n_15427;
wire n_8244;
wire n_13134;
wire n_13340;
wire n_6977;
wire n_7229;
wire n_12688;
wire n_11732;
wire n_10485;
wire n_8096;
wire n_11946;
wire n_7336;
wire n_5932;
wire n_11334;
wire n_6598;
wire n_10105;
wire n_6795;
wire n_6121;
wire n_11855;
wire n_12321;
wire n_5919;
wire n_8346;
wire n_6614;
wire n_5012;
wire n_6506;
wire n_11781;
wire n_13310;
wire n_14548;
wire n_14306;
wire n_15765;
wire n_11080;
wire n_9705;
wire n_4967;
wire n_8367;
wire n_4696;
wire n_9113;
wire n_10761;
wire n_12104;
wire n_14074;
wire n_6001;
wire n_14043;
wire n_13445;
wire n_14676;
wire n_4971;
wire n_9521;
wire n_9682;
wire n_7493;
wire n_9278;
wire n_5664;
wire n_15967;
wire n_6406;
wire n_5890;
wire n_14355;
wire n_14025;
wire n_4661;
wire n_5823;
wire n_8898;
wire n_8658;
wire n_9222;
wire n_5944;
wire n_8905;
wire n_5422;
wire n_15174;
wire n_15939;
wire n_6989;
wire n_8145;
wire n_8237;
wire n_6299;
wire n_11445;
wire n_12643;
wire n_10592;
wire n_9813;
wire n_7424;
wire n_10216;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_9863;
wire n_15348;
wire n_10616;
wire n_11350;
wire n_14527;
wire n_12799;
wire n_13833;
wire n_15022;
wire n_12202;
wire n_12694;
wire n_11057;
wire n_9394;
wire n_10170;
wire n_11182;
wire n_4305;
wire n_11140;
wire n_16213;
wire n_11082;
wire n_15754;
wire n_7273;
wire n_9663;
wire n_7901;
wire n_14371;
wire n_15759;
wire n_5725;
wire n_10146;
wire n_5404;
wire n_15378;
wire n_16060;
wire n_15287;
wire n_10175;
wire n_11949;
wire n_13576;
wire n_12055;
wire n_4834;
wire n_9994;
wire n_5332;
wire n_7149;
wire n_9723;
wire n_15095;
wire n_7116;
wire n_16270;
wire n_4692;
wire n_15153;
wire n_11693;
wire n_12506;
wire n_8211;
wire n_8537;
wire n_15670;
wire n_15717;
wire n_8946;
wire n_5616;
wire n_8055;
wire n_10848;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_12788;
wire n_12894;
wire n_6053;
wire n_11024;
wire n_6233;
wire n_10450;
wire n_10918;
wire n_12333;
wire n_13502;
wire n_4299;
wire n_15254;
wire n_14879;
wire n_13131;
wire n_5625;
wire n_13238;
wire n_14597;
wire n_6758;
wire n_14801;
wire n_5367;
wire n_9069;
wire n_12866;
wire n_6629;
wire n_5288;
wire n_16122;
wire n_13247;
wire n_11158;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_4965;
wire n_7601;
wire n_8998;
wire n_13391;
wire n_15561;
wire n_14190;
wire n_11046;
wire n_15529;
wire n_7033;
wire n_16092;
wire n_16009;
wire n_6010;
wire n_4178;
wire n_11390;
wire n_15296;
wire n_12551;
wire n_11224;
wire n_13970;
wire n_10536;
wire n_15604;
wire n_14696;
wire n_8157;
wire n_9284;
wire n_4953;
wire n_10990;
wire n_8484;
wire n_4813;
wire n_12223;
wire n_12390;
wire n_12627;
wire n_15794;
wire n_7147;
wire n_9556;
wire n_7596;
wire n_12226;
wire n_14546;
wire n_5294;
wire n_11380;
wire n_8161;
wire n_5570;
wire n_11101;
wire n_6411;
wire n_11578;
wire n_9337;
wire n_5411;
wire n_5670;
wire n_16041;
wire n_13256;
wire n_11015;
wire n_11214;
wire n_9211;
wire n_12378;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_10278;
wire n_4793;
wire n_4802;
wire n_10482;
wire n_14174;
wire n_6032;
wire n_10996;
wire n_5733;
wire n_8692;
wire n_12794;
wire n_4897;
wire n_9243;
wire n_14046;
wire n_12436;
wire n_6918;
wire n_10733;
wire n_16244;
wire n_9773;
wire n_14158;
wire n_4674;
wire n_15127;
wire n_15724;
wire n_8812;
wire n_14218;
wire n_11033;
wire n_8682;
wire n_13170;
wire n_4796;
wire n_8290;
wire n_7138;
wire n_13664;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_9928;
wire n_10975;
wire n_11950;
wire n_8890;
wire n_10484;
wire n_12962;
wire n_8747;
wire n_7617;
wire n_12094;
wire n_4575;
wire n_9784;
wire n_11115;
wire n_10641;
wire n_12964;
wire n_8062;
wire n_14120;
wire n_7137;
wire n_5061;
wire n_14652;
wire n_14412;
wire n_14499;
wire n_4653;
wire n_7700;
wire n_11709;
wire n_15431;
wire n_15491;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_14938;
wire n_10584;
wire n_16222;
wire n_14609;
wire n_8667;
wire n_4581;
wire n_9192;
wire n_14466;
wire n_10365;
wire n_14427;
wire n_6008;
wire n_10778;
wire n_4625;
wire n_11542;
wire n_11607;
wire n_7098;
wire n_6181;
wire n_14668;
wire n_5070;
wire n_4845;
wire n_13105;
wire n_4148;
wire n_9134;
wire n_12838;
wire n_13964;
wire n_5575;
wire n_6654;
wire n_11491;
wire n_7661;
wire n_4968;
wire n_7801;
wire n_8807;
wire n_9975;
wire n_13766;
wire n_9765;
wire n_11896;
wire n_13525;
wire n_6907;
wire n_4590;
wire n_5177;
wire n_11371;
wire n_11939;
wire n_7876;
wire n_5316;
wire n_14332;
wire n_4214;
wire n_13081;
wire n_10378;
wire n_5290;
wire n_13057;
wire n_15067;
wire n_10324;
wire n_11563;
wire n_7323;
wire n_15223;
wire n_13861;
wire n_10850;
wire n_5048;
wire n_11565;
wire n_13129;
wire n_13257;
wire n_15395;
wire n_5363;
wire n_14583;
wire n_11164;
wire n_12633;
wire n_5665;
wire n_6517;
wire n_11401;
wire n_11414;
wire n_4892;
wire n_6339;
wire n_10330;
wire n_12514;
wire n_15136;
wire n_14408;
wire n_14659;
wire n_16034;
wire n_9564;
wire n_14267;
wire n_9127;
wire n_11199;
wire n_15540;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_14370;
wire n_5607;
wire n_7929;
wire n_14516;
wire n_14840;
wire n_15692;
wire n_11319;
wire n_9306;
wire n_4353;
wire n_8212;
wire n_4950;
wire n_10442;
wire n_7755;
wire n_14970;
wire n_6504;
wire n_9891;
wire n_13865;
wire n_13135;
wire n_10962;
wire n_10022;
wire n_13973;
wire n_4176;
wire n_9078;
wire n_7556;
wire n_11415;
wire n_13553;
wire n_4124;
wire n_4431;
wire n_15005;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_10972;
wire n_6814;
wire n_7216;
wire n_13248;
wire n_4488;
wire n_10127;
wire n_5278;
wire n_15123;
wire n_14278;
wire n_10824;
wire n_5214;
wire n_11128;
wire n_9332;
wire n_12262;
wire n_12391;
wire n_8043;
wire n_8223;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_8868;
wire n_9889;
wire n_4608;
wire n_9294;
wire n_12731;
wire n_6691;
wire n_13623;
wire n_13775;
wire n_12235;
wire n_4839;
wire n_9174;
wire n_5969;
wire n_10375;
wire n_9132;
wire n_13464;
wire n_4454;
wire n_11669;
wire n_4184;
wire n_15609;
wire n_9547;
wire n_6343;
wire n_12406;
wire n_15213;
wire n_6005;
wire n_6686;
wire n_12929;
wire n_16217;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_14067;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_6025;
wire n_12229;
wire n_15252;
wire n_8434;
wire n_14264;
wire n_15969;
wire n_12508;
wire n_5436;
wire n_7962;
wire n_6697;
wire n_11262;
wire n_16121;
wire n_12271;
wire n_11110;
wire n_12803;
wire n_13084;
wire n_14451;
wire n_14614;
wire n_10122;
wire n_6085;
wire n_10898;
wire n_14785;
wire n_9762;
wire n_11849;
wire n_5341;
wire n_8608;
wire n_13583;
wire n_5140;
wire n_13470;
wire n_12245;
wire n_16218;
wire n_6062;
wire n_4541;
wire n_14394;
wire n_15430;
wire n_6715;
wire n_15872;
wire n_16110;
wire n_8656;
wire n_15414;
wire n_5096;
wire n_9183;
wire n_11287;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_11247;
wire n_5847;
wire n_7204;
wire n_12376;
wire n_9461;
wire n_9117;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_12773;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_4665;
wire n_7476;
wire n_10116;
wire n_10991;
wire n_10590;
wire n_11945;
wire n_14743;
wire n_11769;
wire n_4884;
wire n_16185;
wire n_12720;
wire n_12736;
wire n_8249;
wire n_4276;
wire n_5268;
wire n_5050;
wire n_9062;
wire n_5503;
wire n_5718;
wire n_7208;
wire n_5240;
wire n_10265;
wire n_7718;
wire n_9915;
wire n_13006;
wire n_11277;
wire n_12459;
wire n_11075;
wire n_5001;
wire n_12708;
wire n_6567;
wire n_11919;
wire n_16063;
wire n_12387;
wire n_13705;
wire n_5658;
wire n_4174;
wire n_9001;
wire n_13599;
wire n_15211;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_13077;
wire n_9081;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_9156;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_10159;
wire n_15643;
wire n_5174;
wire n_9024;
wire n_9198;
wire n_10178;
wire n_4801;
wire n_10571;
wire n_15516;
wire n_6079;
wire n_6260;
wire n_4582;
wire n_14268;
wire n_4774;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_13892;
wire n_14251;
wire n_15911;
wire n_12239;
wire n_15567;
wire n_14136;
wire n_12636;
wire n_14002;
wire n_6671;
wire n_11085;
wire n_9335;
wire n_4740;
wire n_16047;
wire n_10550;
wire n_9488;
wire n_16090;
wire n_7632;
wire n_4394;
wire n_15850;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_16112;
wire n_11510;
wire n_9725;
wire n_8842;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_10185;
wire n_12648;
wire n_9526;
wire n_4920;
wire n_10809;
wire n_13316;
wire n_4220;
wire n_13140;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_10660;
wire n_13162;
wire n_15308;
wire n_12501;
wire n_5610;
wire n_9962;
wire n_15848;
wire n_8576;
wire n_12755;
wire n_15869;
wire n_6703;
wire n_14262;
wire n_10657;
wire n_10627;
wire n_8799;
wire n_4378;
wire n_9667;
wire n_5166;
wire n_11256;
wire n_6065;
wire n_7265;
wire n_12441;
wire n_14018;
wire n_14805;
wire n_14935;
wire n_4180;
wire n_11516;
wire n_11520;
wire n_15376;
wire n_4459;
wire n_6878;
wire n_11461;
wire n_11137;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_15309;
wire n_6527;
wire n_4594;
wire n_13604;
wire n_14877;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_14029;
wire n_13157;
wire n_11536;
wire n_15790;
wire n_11544;
wire n_14488;
wire n_10897;
wire n_4642;
wire n_13952;
wire n_14234;
wire n_9716;
wire n_6913;
wire n_15502;
wire n_7473;
wire n_7242;
wire n_9253;
wire n_6533;
wire n_11305;
wire n_14126;
wire n_15352;
wire n_7164;
wire n_15890;
wire n_15164;
wire n_15804;
wire n_15959;
wire n_8022;
wire n_10617;
wire n_12011;
wire n_6845;
wire n_10451;
wire n_8227;
wire n_5300;
wire n_14438;
wire n_10768;
wire n_7853;
wire n_11268;
wire n_13707;
wire n_5233;
wire n_12742;
wire n_10309;
wire n_5381;
wire n_15569;
wire n_9796;
wire n_5770;
wire n_7483;
wire n_13868;
wire n_8756;
wire n_5710;
wire n_10021;
wire n_9953;
wire n_7389;
wire n_10053;
wire n_10315;
wire n_16125;
wire n_5333;
wire n_5799;
wire n_10765;
wire n_6265;
wire n_4914;
wire n_12317;
wire n_8604;
wire n_12831;
wire n_8809;
wire n_13092;
wire n_8976;
wire n_11815;
wire n_13694;
wire n_10907;
wire n_7046;
wire n_13928;
wire n_15135;
wire n_7834;
wire n_10312;
wire n_11299;
wire n_16085;
wire n_4587;
wire n_16116;
wire n_11273;
wire n_8940;
wire n_15416;
wire n_5008;
wire n_9077;
wire n_12872;
wire n_15541;
wire n_13147;
wire n_15879;
wire n_12871;
wire n_13212;
wire n_12590;
wire n_14503;
wire n_14325;
wire n_15644;
wire n_11213;
wire n_13519;
wire n_8844;
wire n_14998;
wire n_6148;
wire n_8995;
wire n_8255;
wire n_5538;
wire n_6357;
wire n_8216;
wire n_8693;
wire n_12785;
wire n_14808;
wire n_5499;
wire n_13661;
wire n_9123;
wire n_4150;
wire n_7811;
wire n_6522;
wire n_12545;
wire n_8669;
wire n_15771;
wire n_4285;
wire n_7097;
wire n_12531;
wire n_7000;
wire n_10486;
wire n_11290;
wire n_15228;
wire n_10357;
wire n_9922;
wire n_5582;
wire n_9177;
wire n_14348;
wire n_5675;
wire n_5109;
wire n_7880;
wire n_14130;
wire n_8769;
wire n_9463;
wire n_6713;
wire n_12916;
wire n_8149;
wire n_10067;
wire n_13163;
wire n_12953;
wire n_15198;
wire n_10698;
wire n_5281;
wire n_6087;
wire n_7851;
wire n_13106;
wire n_13874;
wire n_13246;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_10135;
wire n_13776;
wire n_6108;
wire n_12222;
wire n_10260;
wire n_7664;
wire n_12370;
wire n_6100;
wire n_14329;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_11412;
wire n_7332;
wire n_14428;
wire n_14813;
wire n_8990;
wire n_5862;
wire n_7477;
wire n_14617;
wire n_10268;
wire n_8208;
wire n_7468;
wire n_12692;
wire n_11550;
wire n_13640;
wire n_15965;
wire n_5886;
wire n_9451;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_12976;
wire n_6415;
wire n_8479;
wire n_6783;
wire n_14660;
wire n_4861;
wire n_13984;
wire n_12397;
wire n_8512;
wire n_14524;
wire n_13093;
wire n_9843;
wire n_9710;
wire n_12634;
wire n_13288;
wire n_16104;
wire n_9087;
wire n_4621;
wire n_15896;
wire n_14287;
wire n_4451;
wire n_7845;
wire n_5285;
wire n_11619;
wire n_13086;
wire n_14052;
wire n_14216;
wire n_5564;
wire n_15044;
wire n_12613;
wire n_9956;
wire n_9079;
wire n_5162;
wire n_14925;
wire n_15641;
wire n_5442;
wire n_12946;
wire n_5802;
wire n_9782;
wire n_10049;
wire n_4784;
wire n_14206;
wire n_13012;
wire n_13606;
wire n_13449;
wire n_12901;
wire n_10589;
wire n_6340;
wire n_13099;
wire n_14475;
wire n_9950;
wire n_11019;
wire n_14620;
wire n_7858;
wire n_11580;
wire n_13699;
wire n_12683;
wire n_6103;
wire n_15829;
wire n_14837;
wire n_6392;
wire n_6513;
wire n_11642;
wire n_4613;
wire n_13389;
wire n_14978;
wire n_9197;
wire n_6720;
wire n_12286;
wire n_11076;
wire n_11752;
wire n_5883;
wire n_9140;
wire n_14134;
wire n_13995;
wire n_10785;
wire n_14726;
wire n_13439;
wire n_8401;
wire n_6078;
wire n_14122;
wire n_12146;
wire n_7680;
wire n_14415;
wire n_5630;
wire n_6666;
wire n_9364;
wire n_9452;
wire n_5117;
wire n_4979;
wire n_9398;
wire n_9362;
wire n_13675;
wire n_13483;
wire n_14977;
wire n_6815;
wire n_14321;
wire n_15275;
wire n_9203;
wire n_6207;
wire n_6381;
wire n_9712;
wire n_15201;
wire n_14903;
wire n_9536;
wire n_12054;
wire n_8450;
wire n_9848;
wire n_12081;
wire n_13614;
wire n_14095;
wire n_11202;
wire n_5054;
wire n_6571;
wire n_9460;
wire n_5929;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_14080;
wire n_8324;
wire n_16159;
wire n_11227;
wire n_5975;
wire n_4242;
wire n_4751;
wire n_13814;
wire n_10381;
wire n_9841;
wire n_14502;
wire n_15367;
wire n_12557;
wire n_9772;
wire n_10554;
wire n_10147;
wire n_9057;
wire n_14847;
wire n_7061;
wire n_11860;
wire n_8104;
wire n_7066;
wire n_9068;
wire n_5496;
wire n_7485;
wire n_7174;
wire n_8014;
wire n_12213;
wire n_6661;
wire n_16265;
wire n_10919;
wire n_12646;
wire n_14750;
wire n_4522;
wire n_15350;
wire n_10228;
wire n_14159;
wire n_5991;
wire n_8623;
wire n_14077;
wire n_14518;
wire n_4952;
wire n_9634;
wire n_6967;
wire n_4426;
wire n_15704;
wire n_5956;
wire n_5699;
wire n_15766;
wire n_4362;
wire n_6017;
wire n_9348;
wire n_11125;
wire n_15209;
wire n_15554;
wire n_5920;
wire n_13011;
wire n_12737;
wire n_6125;
wire n_8651;
wire n_5000;
wire n_10699;
wire n_4634;
wire n_9632;
wire n_4932;
wire n_14358;
wire n_12092;
wire n_11951;
wire n_5211;
wire n_9257;
wire n_15017;
wire n_11451;
wire n_11816;
wire n_9500;
wire n_5132;
wire n_9747;
wire n_9470;
wire n_11508;
wire n_6414;
wire n_5535;
wire n_4506;
wire n_6097;
wire n_14467;
wire n_7783;
wire n_11232;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_10188;
wire n_14898;
wire n_9591;
wire n_11138;
wire n_14373;
wire n_9049;
wire n_14912;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_4346;
wire n_13585;
wire n_7003;
wire n_10433;
wire n_8137;
wire n_10231;
wire n_8413;
wire n_10841;
wire n_6302;
wire n_10929;
wire n_12642;
wire n_13142;
wire n_15300;
wire n_13974;
wire n_14656;
wire n_9471;
wire n_6922;
wire n_15185;
wire n_14070;
wire n_14909;
wire n_15772;
wire n_16004;
wire n_15294;
wire n_10582;
wire n_13494;
wire n_12601;
wire n_15210;
wire n_10719;
wire n_8300;
wire n_10747;
wire n_8069;
wire n_10934;
wire n_7501;
wire n_11383;
wire n_9409;
wire n_10711;
wire n_10743;
wire n_11088;
wire n_6432;
wire n_12959;
wire n_7984;
wire n_12899;
wire n_15447;
wire n_12616;
wire n_7366;
wire n_8173;
wire n_4359;
wire n_10481;
wire n_13562;
wire n_13540;
wire n_12919;
wire n_15895;
wire n_7589;
wire n_14953;
wire n_13568;
wire n_13642;
wire n_15379;
wire n_4447;
wire n_14764;
wire n_4293;
wire n_6880;
wire n_6223;
wire n_5176;
wire n_9832;
wire n_12010;
wire n_12314;
wire n_5793;
wire n_14632;
wire n_6926;
wire n_8091;
wire n_13751;
wire n_12394;
wire n_12856;
wire n_5761;
wire n_13465;
wire n_6699;
wire n_12797;
wire n_13683;
wire n_16231;
wire n_13630;
wire n_9067;
wire n_8254;
wire n_8400;
wire n_10141;
wire n_11090;
wire n_14661;
wire n_10305;
wire n_7232;
wire n_15372;
wire n_9858;
wire n_7511;
wire n_10936;
wire n_12134;
wire n_13824;
wire n_12730;
wire n_9482;
wire n_9033;
wire n_6957;
wire n_11429;
wire n_15570;
wire n_5074;
wire n_14624;
wire n_12735;
wire n_14510;
wire n_7917;
wire n_11908;
wire n_4942;
wire n_8368;
wire n_15388;
wire n_6694;
wire n_9247;
wire n_8463;
wire n_9965;
wire n_10425;
wire n_15226;
wire n_15927;
wire n_6449;
wire n_10862;
wire n_12254;
wire n_14333;
wire n_4348;
wire n_7422;
wire n_9299;
wire n_13357;
wire n_8889;
wire n_5681;
wire n_9785;
wire n_9244;
wire n_11298;
wire n_14667;
wire n_16232;
wire n_5261;
wire n_12427;
wire n_12124;
wire n_9195;
wire n_8322;
wire n_11353;
wire n_12494;
wire n_15623;
wire n_6591;
wire n_7466;
wire n_8987;
wire n_13454;
wire n_9280;
wire n_7621;
wire n_9911;
wire n_12051;
wire n_8274;
wire n_13958;
wire n_6594;
wire n_6342;
wire n_6195;
wire n_14802;
wire n_10373;
wire n_6441;
wire n_11116;
wire n_7572;
wire n_7158;
wire n_13637;
wire n_11173;
wire n_11660;
wire n_15675;
wire n_7500;
wire n_12355;
wire n_7985;
wire n_9687;
wire n_4240;
wire n_8657;
wire n_11567;
wire n_8954;
wire n_6354;
wire n_11881;
wire n_10563;
wire n_12458;
wire n_8311;
wire n_15786;
wire n_5748;
wire n_4393;
wire n_11363;
wire n_6662;
wire n_7494;
wire n_9088;
wire n_16250;
wire n_14050;
wire n_8728;
wire n_9580;
wire n_11280;
wire n_9569;
wire n_8994;
wire n_4389;
wire n_6433;
wire n_9680;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_12463;
wire n_12612;
wire n_8407;
wire n_8071;
wire n_13423;
wire n_13046;
wire n_4461;
wire n_11636;
wire n_14926;
wire n_10530;
wire n_6902;
wire n_4615;
wire n_12798;
wire n_7197;
wire n_6369;
wire n_8528;
wire n_14088;
wire n_9227;
wire n_13644;
wire n_5657;
wire n_12510;
wire n_11313;
wire n_14364;
wire n_8475;
wire n_9951;
wire n_15182;
wire n_9855;
wire n_9072;
wire n_12635;
wire n_10102;
wire n_13545;
wire n_12537;
wire n_14913;
wire n_13197;
wire n_5244;
wire n_5765;
wire n_12076;
wire n_5114;
wire n_9054;
wire n_4551;
wire n_15836;
wire n_10117;
wire n_4521;
wire n_13252;
wire n_6956;
wire n_13139;
wire n_10126;
wire n_7587;
wire n_6451;
wire n_12874;
wire n_11920;
wire n_7704;
wire n_10604;
wire n_6497;
wire n_8511;
wire n_5420;
wire n_7865;
wire n_5206;
wire n_13356;
wire n_14447;
wire n_16039;
wire n_4387;
wire n_14237;
wire n_14745;
wire n_9584;
wire n_9287;
wire n_10344;
wire n_10568;
wire n_9459;
wire n_6701;
wire n_5298;
wire n_9490;
wire n_10209;
wire n_8867;
wire n_8246;
wire n_8558;
wire n_9655;
wire n_13769;
wire n_9846;
wire n_12048;
wire n_9593;
wire n_4598;
wire n_4464;
wire n_12072;
wire n_8925;
wire n_5106;
wire n_7881;
wire n_11317;
wire n_9147;
wire n_13339;
wire n_15854;
wire n_4789;
wire n_14433;
wire n_12829;
wire n_14672;
wire n_9678;
wire n_10803;
wire n_12132;
wire n_13626;
wire n_11903;
wire n_8641;
wire n_9658;
wire n_10299;
wire n_9560;
wire n_15036;
wire n_12528;
wire n_9578;
wire n_11813;
wire n_14195;
wire n_5080;
wire n_9396;
wire n_7032;
wire n_4565;
wire n_12745;
wire n_16061;
wire n_9303;
wire n_12371;
wire n_11811;
wire n_12841;
wire n_7198;
wire n_12417;
wire n_14866;
wire n_6884;
wire n_7752;
wire n_10618;
wire n_10836;
wire n_11378;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_12180;
wire n_12049;
wire n_7953;
wire n_6106;
wire n_14434;
wire n_16086;
wire n_6876;
wire n_15746;
wire n_9553;
wire n_12603;
wire n_8046;
wire n_4552;
wire n_14964;
wire n_12978;
wire n_7193;
wire n_6287;
wire n_14575;
wire n_10930;
wire n_6172;
wire n_14005;
wire n_9942;
wire n_9805;
wire n_13686;
wire n_4482;
wire n_5957;
wire n_4172;
wire n_12466;
wire n_13842;
wire n_16220;
wire n_8414;
wire n_5567;
wire n_8292;
wire n_9138;
wire n_9879;
wire n_5406;
wire n_8647;
wire n_11936;
wire n_6362;
wire n_9213;
wire n_12071;
wire n_4328;
wire n_12982;
wire n_8543;
wire n_14680;
wire n_13459;
wire n_11543;
wire n_15637;
wire n_11184;
wire n_11795;
wire n_5191;
wire n_11391;
wire n_6067;
wire n_11646;
wire n_6833;
wire n_4940;
wire n_15156;
wire n_9374;
wire n_13649;
wire n_14720;
wire n_14497;
wire n_8331;
wire n_8317;
wire n_7126;
wire n_12578;
wire n_12311;
wire n_11963;
wire n_5867;
wire n_14109;
wire n_13253;
wire n_12985;
wire n_12232;
wire n_15316;
wire n_5085;
wire n_12640;
wire n_7496;
wire n_13729;
wire n_15027;
wire n_6430;
wire n_11435;
wire n_13647;
wire n_9179;
wire n_6296;
wire n_10014;
wire n_11056;
wire n_14241;
wire n_10714;
wire n_5602;
wire n_7196;
wire n_4928;
wire n_14855;
wire n_12101;
wire n_11120;
wire n_11185;
wire n_7360;
wire n_5428;
wire n_10895;
wire n_6325;
wire n_10916;
wire n_14693;
wire n_12197;
wire n_12497;
wire n_4865;
wire n_15611;
wire n_6678;
wire n_7982;
wire n_10838;
wire n_13002;
wire n_6564;
wire n_7268;
wire n_8187;
wire n_8174;
wire n_8929;
wire n_10108;
wire n_14069;
wire n_4436;
wire n_15196;
wire n_5822;
wire n_5786;
wire n_15964;
wire n_10661;
wire n_8846;
wire n_5817;
wire n_9277;
wire n_4160;
wire n_14754;
wire n_15151;
wire n_15111;
wire n_6109;
wire n_9611;
wire n_6385;
wire n_12571;
wire n_9744;
wire n_5798;
wire n_10123;
wire n_4137;
wire n_13022;
wire n_15949;
wire n_8032;
wire n_9504;
wire n_5417;
wire n_14118;
wire n_14445;
wire n_11147;
wire n_10048;
wire n_4545;
wire n_11194;
wire n_8200;
wire n_4758;
wire n_9285;
wire n_8036;
wire n_15068;
wire n_15590;
wire n_5713;
wire n_4840;
wire n_9905;
wire n_10963;
wire n_11016;
wire n_12228;
wire n_11146;
wire n_13088;
wire n_4395;
wire n_4873;
wire n_10788;
wire n_16161;
wire n_14142;
wire n_9190;
wire n_8586;
wire n_15937;
wire n_8524;
wire n_11924;
wire n_12540;
wire n_4535;
wire n_7518;
wire n_8828;
wire n_9639;
wire n_10422;
wire n_4385;
wire n_12001;
wire n_15916;
wire n_7779;
wire n_12059;
wire n_9664;
wire n_13275;
wire n_11830;
wire n_14577;
wire n_4731;
wire n_7575;
wire n_11489;
wire n_7073;
wire n_13026;
wire n_15753;
wire n_8092;
wire n_10471;
wire n_13760;
wire n_12479;
wire n_16087;
wire n_10979;
wire n_6309;
wire n_8370;
wire n_9109;
wire n_10189;
wire n_13820;
wire n_8135;
wire n_12702;
wire n_6519;
wire n_4671;
wire n_14366;
wire n_9741;
wire n_5989;
wire n_5571;
wire n_4766;
wire n_10569;
wire n_4558;
wire n_13116;
wire n_13663;
wire n_10686;
wire n_14055;
wire n_14197;
wire n_16153;
wire n_8764;
wire n_14454;
wire n_7349;
wire n_9875;
wire n_8502;
wire n_10713;
wire n_11411;
wire n_4319;
wire n_9360;
wire n_6585;
wire n_12211;
wire n_14323;
wire n_7786;
wire n_10913;
wire n_9021;
wire n_8454;
wire n_12306;
wire n_4358;
wire n_11145;
wire n_9122;
wire n_7579;
wire n_10099;
wire n_7122;
wire n_12637;
wire n_12335;
wire n_10193;
wire n_14096;
wire n_4874;
wire n_4904;
wire n_10203;
wire n_10140;
wire n_13982;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_11000;
wire n_10149;
wire n_10920;
wire n_11712;
wire n_14068;
wire n_4748;
wire n_14019;
wire n_7624;
wire n_13405;
wire n_9803;
wire n_13828;
wire n_14397;
wire n_15738;
wire n_8776;
wire n_10576;
wire n_8564;
wire n_12114;
wire n_8343;
wire n_7828;
wire n_14319;
wire n_4618;
wire n_6721;
wire n_15106;
wire n_13102;
wire n_8718;
wire n_14301;
wire n_13550;
wire n_14910;
wire n_10682;
wire n_16198;
wire n_5506;
wire n_7543;
wire n_9659;
wire n_12204;
wire n_13643;
wire n_15997;
wire n_15812;
wire n_16252;
wire n_8042;
wire n_5475;
wire n_7727;
wire n_14774;
wire n_5908;
wire n_9013;
wire n_5431;
wire n_9427;
wire n_12325;
wire n_8379;
wire n_8034;
wire n_12143;
wire n_7778;
wire n_5100;
wire n_10225;
wire n_9126;
wire n_7019;
wire n_5315;
wire n_5752;
wire n_9474;
wire n_8441;
wire n_14026;
wire n_14362;
wire n_7702;
wire n_14114;
wire n_5746;
wire n_10368;
wire n_4910;
wire n_4724;
wire n_10237;
wire n_14504;
wire n_9538;
wire n_6685;
wire n_14930;
wire n_8569;
wire n_9574;
wire n_10531;
wire n_12032;
wire n_4666;
wire n_12066;
wire n_14471;
wire n_8592;
wire n_8865;
wire n_7952;
wire n_11170;
wire n_7347;
wire n_9450;
wire n_10031;
wire n_6016;
wire n_4466;
wire n_9998;
wire n_13963;
wire n_15568;
wire n_15948;
wire n_5366;
wire n_11523;
wire n_5322;
wire n_11121;
wire n_12176;
wire n_5414;
wire n_11805;
wire n_13266;
wire n_7791;
wire n_8362;
wire n_6971;
wire n_10847;
wire n_8632;
wire n_10035;
wire n_14242;
wire n_14523;
wire n_15660;
wire n_7739;
wire n_12740;
wire n_7945;
wire n_9372;
wire n_9045;
wire n_15040;
wire n_16233;
wire n_8361;
wire n_9657;
wire n_7656;
wire n_11457;
wire n_14883;
wire n_5903;
wire n_7199;
wire n_10107;
wire n_11725;
wire n_10283;
wire n_5151;
wire n_15731;
wire n_5307;
wire n_9904;
wire n_4721;
wire n_12344;
wire n_14937;
wire n_9924;
wire n_9159;
wire n_8561;
wire n_6549;
wire n_9326;
wire n_8611;
wire n_8410;
wire n_15486;
wire n_16225;
wire n_5003;
wire n_6540;
wire n_7166;
wire n_6658;
wire n_11694;
wire n_5369;
wire n_9476;
wire n_6683;
wire n_15634;
wire n_4921;
wire n_5912;
wire n_11540;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_10050;
wire n_14800;
wire n_11058;
wire n_5156;
wire n_15743;
wire n_5803;
wire n_6327;
wire n_8878;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_5779;
wire n_12203;
wire n_15606;
wire n_16156;
wire n_11403;
wire n_8492;
wire n_9301;
wire n_14099;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_10392;
wire n_14041;
wire n_12769;
wire n_15076;
wire n_8888;
wire n_6820;
wire n_5446;
wire n_11741;
wire n_7610;
wire n_7107;
wire n_11245;
wire n_4561;
wire n_14225;
wire n_7456;
wire n_9382;
wire n_11784;
wire n_8095;
wire n_15426;
wire n_11365;
wire n_13291;
wire n_14756;
wire n_9921;
wire n_7369;
wire n_15559;
wire n_14888;
wire n_9325;
wire n_9945;
wire n_9643;
wire n_7548;
wire n_11005;
wire n_13016;
wire n_12820;
wire n_8735;
wire n_15073;
wire n_7598;
wire n_7250;
wire n_8808;
wire n_9201;
wire n_8902;
wire n_7823;
wire n_9771;
wire n_8833;
wire n_14605;
wire n_12869;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_14413;
wire n_16154;
wire n_4879;
wire n_13435;
wire n_16031;
wire n_8794;
wire n_12689;
wire n_11074;
wire n_5044;
wire n_4536;
wire n_9894;
wire n_9274;
wire n_11141;
wire n_12750;
wire n_14753;
wire n_15936;
wire n_8549;
wire n_14161;
wire n_6676;
wire n_4304;
wire n_10095;
wire n_4927;
wire n_5459;
wire n_14285;
wire n_10716;
wire n_11102;
wire n_12171;
wire n_14812;
wire n_14000;
wire n_10088;
wire n_11238;
wire n_11406;
wire n_16000;
wire n_10443;
wire n_10488;
wire n_7525;
wire n_16251;
wire n_4418;
wire n_7924;
wire n_11103;
wire n_12420;
wire n_9232;
wire n_8690;
wire n_4125;
wire n_5390;
wire n_12954;
wire n_5351;
wire n_5267;
wire n_11852;
wire n_5024;
wire n_7012;
wire n_12500;
wire n_15393;
wire n_8593;
wire n_11837;
wire n_10912;
wire n_13501;
wire n_10469;
wire n_15958;
wire n_13533;
wire n_9649;
wire n_11684;
wire n_5275;
wire n_12112;
wire n_15377;
wire n_15864;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_6923;
wire n_4412;
wire n_7649;
wire n_8195;
wire n_8009;
wire n_8588;
wire n_16027;
wire n_15628;
wire n_9839;
wire n_10887;
wire n_12004;
wire n_6704;
wire n_7634;
wire n_9090;
wire n_7406;
wire n_13520;
wire n_4682;
wire n_9346;
wire n_11012;
wire n_6673;
wire n_14480;
wire n_9696;
wire n_11041;
wire n_14181;
wire n_10742;
wire n_14024;
wire n_11798;
wire n_12614;
wire n_13165;
wire n_15312;
wire n_9996;
wire n_6534;
wire n_9968;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_4957;
wire n_15576;
wire n_6127;
wire n_4855;
wire n_9383;
wire n_9498;
wire n_10405;
wire n_6246;
wire n_10390;
wire n_11978;
wire n_10989;
wire n_9836;
wire n_5005;
wire n_14570;
wire n_14702;
wire n_11827;
wire n_10328;
wire n_16191;
wire n_13315;
wire n_10692;
wire n_15118;
wire n_6126;
wire n_7372;
wire n_8596;
wire n_9938;
wire n_12912;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_15592;
wire n_10867;
wire n_6841;
wire n_11847;
wire n_10206;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_11281;
wire n_12957;
wire n_5624;
wire n_10092;
wire n_4601;
wire n_4518;
wire n_7009;
wire n_5474;
wire n_11772;
wire n_15837;
wire n_9743;
wire n_9121;
wire n_7371;
wire n_13448;
wire n_11237;
wire n_14752;
wire n_9509;
wire n_5447;
wire n_12153;
wire n_12005;
wire n_7463;
wire n_9621;
wire n_15966;
wire n_10738;
wire n_4308;
wire n_5755;
wire n_5700;
wire n_11851;
wire n_9158;
wire n_4325;
wire n_14239;
wire n_14501;
wire n_4711;
wire n_6889;
wire n_16068;
wire n_12586;
wire n_11993;
wire n_5962;
wire n_15710;
wire n_4413;
wire n_11131;
wire n_12221;
wire n_8627;
wire n_14318;
wire n_11432;
wire n_12302;
wire n_8945;
wire n_9142;
wire n_13628;
wire n_9216;
wire n_9189;
wire n_6723;
wire n_7398;
wire n_9563;
wire n_7941;
wire n_4135;
wire n_15229;
wire n_12757;
wire n_13010;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_13251;
wire n_14738;
wire n_8858;
wire n_12107;
wire n_11738;
wire n_11595;
wire n_13504;
wire n_13521;
wire n_14404;
wire n_12695;
wire n_11512;
wire n_5801;
wire n_14163;
wire n_15504;
wire n_12349;
wire n_6054;
wire n_13703;
wire n_4821;
wire n_14758;
wire n_13161;
wire n_7011;
wire n_10813;
wire n_15403;
wire n_14076;
wire n_10986;
wire n_11603;
wire n_15573;
wire n_6393;
wire n_14291;
wire n_14761;
wire n_12380;
wire n_7074;
wire n_10853;
wire n_8916;
wire n_10899;
wire n_11707;
wire n_11728;
wire n_13352;
wire n_11521;
wire n_13309;
wire n_5465;
wire n_16137;
wire n_12577;
wire n_10575;
wire n_8745;
wire n_5154;
wire n_14388;
wire n_5721;
wire n_8169;
wire n_14932;
wire n_6184;
wire n_8018;
wire n_11802;
wire n_9984;
wire n_4138;
wire n_7083;
wire n_15889;
wire n_8260;
wire n_12723;
wire n_10334;
wire n_14153;
wire n_12135;
wire n_14674;
wire n_7143;
wire n_7701;
wire n_11688;
wire n_13484;
wire n_8688;
wire n_9794;
wire n_15761;
wire n_7969;
wire n_16062;
wire n_10726;
wire n_16210;
wire n_8279;
wire n_4384;
wire n_8793;
wire n_4639;
wire n_12864;
wire n_13486;
wire n_10388;
wire n_4577;
wire n_6312;
wire n_13478;
wire n_7683;
wire n_9550;
wire n_13108;
wire n_11042;
wire n_15701;
wire n_12570;
wire n_14124;
wire n_15932;
wire n_10510;
wire n_14344;
wire n_7669;
wire n_8298;
wire n_6711;
wire n_6818;
wire n_11696;
wire n_15802;
wire n_6438;
wire n_11761;
wire n_4481;
wire n_5087;
wire n_10635;
wire n_11681;
wire n_7209;
wire n_13429;
wire n_6193;
wire n_13897;
wire n_8023;
wire n_9319;
wire n_7330;
wire n_6007;
wire n_13374;
wire n_13182;
wire n_6734;
wire n_10852;
wire n_6535;
wire n_14867;
wire n_14893;
wire n_13789;
wire n_8053;
wire n_11407;
wire n_15893;
wire n_8059;
wire n_9871;
wire n_14354;
wire n_6879;
wire n_9562;
wire n_15442;
wire n_15632;
wire n_9896;
wire n_9612;
wire n_6208;
wire n_7190;
wire n_9698;
wire n_6303;
wire n_6014;
wire n_15840;
wire n_4270;
wire n_7692;
wire n_9528;
wire n_10241;
wire n_4620;
wire n_6255;
wire n_6457;
wire n_5397;
wire n_13690;
wire n_9272;
wire n_13055;
wire n_14379;
wire n_9955;
wire n_15451;
wire n_9645;
wire n_15953;
wire n_4924;
wire n_8372;
wire n_6270;
wire n_14283;
wire n_8737;
wire n_9731;
wire n_10026;
wire n_15999;
wire n_5996;
wire n_13577;
wire n_5566;
wire n_9697;
wire n_7288;
wire n_15307;
wire n_10772;
wire n_4388;
wire n_13098;
wire n_10901;
wire n_7362;
wire n_15855;
wire n_14942;
wire n_7082;
wire n_7237;
wire n_8988;
wire n_10664;
wire n_7131;
wire n_6276;
wire n_15661;
wire n_12328;
wire n_13839;
wire n_9642;
wire n_8723;
wire n_11189;
wire n_12559;
wire n_9929;
wire n_9050;
wire n_4406;
wire n_4271;
wire n_12056;
wire n_13898;
wire n_15030;
wire n_16204;
wire n_7042;
wire n_9859;
wire n_8419;
wire n_10767;
wire n_10320;
wire n_5652;
wire n_13380;
wire n_8893;
wire n_5805;
wire n_7304;
wire n_11910;
wire n_16235;
wire n_6266;
wire n_15386;
wire n_12109;
wire n_14457;
wire n_14905;
wire n_9531;
wire n_10521;
wire n_8077;
wire n_5492;
wire n_11242;
wire n_5501;
wire n_12917;
wire n_14711;
wire n_15445;
wire n_6934;
wire n_13188;
wire n_14179;
wire n_13362;
wire n_7386;
wire n_7391;
wire n_15259;
wire n_4401;
wire n_11361;
wire n_7754;
wire n_11894;
wire n_12058;
wire n_8826;
wire n_13819;
wire n_7023;
wire n_10872;
wire n_13990;
wire n_15745;
wire n_9732;
wire n_5758;
wire n_5842;
wire n_12083;
wire n_9685;
wire n_12529;
wire n_15521;
wire n_10374;
wire n_11253;
wire n_13983;
wire n_12045;
wire n_13193;
wire n_14995;
wire n_15856;
wire n_7404;
wire n_10345;
wire n_8959;
wire n_15648;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_12471;
wire n_4973;
wire n_13802;
wire n_13781;
wire n_15887;
wire n_7981;
wire n_4792;
wire n_13037;
wire n_4402;
wire n_14252;
wire n_14736;
wire n_15058;
wire n_15351;
wire n_12188;
wire n_14851;
wire n_5473;
wire n_12575;
wire n_10601;
wire n_14698;
wire n_11623;
wire n_8712;
wire n_12473;
wire n_10372;
wire n_15394;
wire n_6352;
wire n_11124;
wire n_14295;
wire n_4286;
wire n_9378;
wire n_6211;
wire n_10448;
wire n_15100;
wire n_8109;
wire n_10301;
wire n_11977;
wire n_15487;
wire n_10074;
wire n_12040;
wire n_13127;
wire n_9389;
wire n_12598;
wire n_5562;
wire n_4858;
wire n_6093;
wire n_5370;
wire n_10001;
wire n_13561;
wire n_7378;
wire n_15922;
wire n_9623;
wire n_4435;
wire n_5317;
wire n_5458;
wire n_14944;
wire n_15987;
wire n_15562;
wire n_7877;
wire n_14336;
wire n_11351;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_12626;
wire n_11094;
wire n_10960;
wire n_10712;
wire n_8007;
wire n_13911;
wire n_14313;
wire n_15578;
wire n_4318;
wire n_13961;
wire n_13343;
wire n_12546;
wire n_8910;
wire n_16070;
wire n_5227;
wire n_14091;
wire n_14842;
wire n_15981;
wire n_10100;
wire n_5902;
wire n_9164;
wire n_6402;
wire n_5359;
wire n_4673;
wire n_11366;
wire n_5282;
wire n_9387;
wire n_8301;
wire n_6764;
wire n_7871;
wire n_14512;
wire n_13539;
wire n_10162;
wire n_9840;
wire n_15982;
wire n_15471;
wire n_7016;
wire n_4738;
wire n_12100;
wire n_11399;
wire n_8892;
wire n_9637;
wire n_5386;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_10535;
wire n_12676;
wire n_10674;
wire n_13584;
wire n_9491;
wire n_13107;
wire n_6955;
wire n_7563;
wire n_10337;
wire n_10774;
wire n_5952;
wire n_7180;
wire n_14655;
wire n_10407;
wire n_14850;
wire n_16253;
wire n_10577;
wire n_14481;
wire n_13778;
wire n_16171;
wire n_8972;
wire n_14531;
wire n_8494;
wire n_12999;
wire n_14709;
wire n_10264;
wire n_15148;
wire n_6569;
wire n_7919;
wire n_13740;
wire n_15355;
wire n_9992;
wire n_14606;
wire n_14089;
wire n_8278;
wire n_8180;
wire n_11549;
wire n_14437;
wire n_12362;
wire n_13913;
wire n_7031;
wire n_13367;
wire n_5716;
wire n_10313;
wire n_10843;
wire n_12983;
wire n_14003;
wire n_8941;
wire n_10771;
wire n_8891;
wire n_7103;
wire n_12360;
wire n_13570;
wire n_6605;
wire n_10724;
wire n_5888;
wire n_9266;
wire n_14409;
wire n_16182;
wire n_8270;
wire n_16103;
wire n_8231;
wire n_4181;
wire n_12313;
wire n_11983;
wire n_6832;
wire n_12604;
wire n_5980;
wire n_8683;
wire n_15885;
wire n_15114;
wire n_9391;
wire n_12558;
wire n_15503;
wire n_15053;
wire n_10445;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_13284;
wire n_6544;
wire n_8810;
wire n_12596;
wire n_6469;
wire n_12840;
wire n_5036;
wire n_11119;
wire n_12696;
wire n_6332;
wire n_15241;
wire n_10863;
wire n_10958;
wire n_11215;
wire n_13730;
wire n_5790;
wire n_7130;
wire n_10174;
wire n_6680;
wire n_15729;
wire n_4647;
wire n_13960;
wire n_6310;
wire n_8932;
wire n_8264;
wire n_12435;
wire n_9695;
wire n_7134;
wire n_8288;
wire n_13411;
wire n_11954;
wire n_14629;
wire n_14778;
wire n_15891;
wire n_16240;
wire n_11526;
wire n_13438;
wire n_14010;
wire n_11591;
wire n_10403;
wire n_11972;
wire n_4142;
wire n_5118;
wire n_9834;
wire n_5485;
wire n_9901;
wire n_5525;
wire n_7102;
wire n_10015;
wire n_10076;
wire n_6259;
wire n_14432;
wire n_15371;
wire n_5271;
wire n_4849;
wire n_13410;
wire n_7133;
wire n_9800;
wire n_10745;
wire n_6289;
wire n_6651;
wire n_9255;
wire n_8882;
wire n_14308;
wire n_12460;
wire n_6565;
wire n_5194;
wire n_12733;
wire n_15532;
wire n_8388;
wire n_5445;
wire n_8067;
wire n_13600;
wire n_8385;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_15061;
wire n_8670;
wire n_4504;
wire n_10460;
wire n_14299;
wire n_14215;
wire n_7813;
wire n_4917;
wire n_7706;
wire n_13332;
wire n_8142;
wire n_14265;
wire n_15266;
wire n_13942;
wire n_7992;
wire n_9085;
wire n_7643;
wire n_15381;
wire n_15090;
wire n_11204;
wire n_6836;
wire n_12939;
wire n_9120;
wire n_6595;
wire n_10415;
wire n_11302;
wire n_16089;
wire n_9899;
wire n_12374;
wire n_15054;
wire n_15398;
wire n_9136;
wire n_16081;
wire n_12261;
wire n_6186;
wire n_11561;
wire n_10227;
wire n_13490;
wire n_14198;
wire n_14836;
wire n_7628;
wire n_13381;
wire n_5628;
wire n_9436;
wire n_5245;
wire n_4489;
wire n_14013;
wire n_15220;
wire n_11385;
wire n_12065;
wire n_13204;
wire n_5329;
wire n_12275;
wire n_8224;
wire n_6035;
wire n_5472;
wire n_9042;
wire n_10884;
wire n_13375;
wire n_15669;
wire n_9570;
wire n_7236;
wire n_9239;
wire n_4833;
wire n_6405;
wire n_8345;
wire n_11054;
wire n_11777;
wire n_9644;
wire n_5850;
wire n_9343;
wire n_8614;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_9131;
wire n_13286;
wire n_9060;
wire n_9792;
wire n_15826;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_14204;
wire n_13384;
wire n_11325;
wire n_10801;
wire n_6769;
wire n_10325;
wire n_13013;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_8951;
wire n_11217;
wire n_15744;
wire n_13582;
wire n_12752;
wire n_10327;
wire n_8700;
wire n_6766;
wire n_4185;
wire n_5940;
wire n_14157;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_11651;
wire n_6232;
wire n_13255;
wire n_4676;
wire n_15144;
wire n_7802;
wire n_7519;
wire n_10505;
wire n_12979;
wire n_14140;
wire n_7457;
wire n_14723;
wire n_11196;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_14933;
wire n_4756;
wire n_15851;
wire n_5860;
wire n_15262;
wire n_11672;
wire n_11557;
wire n_9982;
wire n_11552;
wire n_6416;
wire n_13682;
wire n_8468;
wire n_9031;
wire n_12715;
wire n_12910;
wire n_7515;
wire n_7639;
wire n_11084;
wire n_12787;
wire n_8933;
wire n_6214;
wire n_8636;
wire n_9006;
wire n_10408;
wire n_11442;
wire n_9221;
wire n_13424;
wire n_4365;
wire n_14102;
wire n_4349;
wire n_10514;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_14603;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_10091;
wire n_11195;
wire n_4198;
wire n_7172;
wire n_10562;
wire n_10586;
wire n_10893;
wire n_8283;
wire n_6225;
wire n_4373;
wire n_7914;
wire n_8860;
wire n_16243;
wire n_15052;
wire n_12401;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_14104;
wire n_4390;
wire n_10593;
wire n_13304;
wire n_11517;
wire n_7892;
wire n_15078;
wire n_12722;
wire n_13716;
wire n_9523;
wire n_10821;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_11918;
wire n_14561;
wire n_13460;
wire n_4453;
wire n_6219;
wire n_15484;
wire n_7674;
wire n_8686;
wire n_13590;
wire n_12712;
wire n_15494;
wire n_10961;
wire n_6175;
wire n_6445;
wire n_9829;
wire n_15778;
wire n_8563;
wire n_11077;
wire n_4571;
wire n_13914;
wire n_11579;
wire n_14887;
wire n_10197;
wire n_16207;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_14119;
wire n_13670;
wire n_13148;
wire n_14962;
wire n_15792;
wire n_10950;
wire n_6499;
wire n_9411;
wire n_12209;
wire n_7983;
wire n_5311;
wire n_8765;
wire n_14168;
wire n_14494;
wire n_15946;
wire n_13452;
wire n_14506;
wire n_5164;
wire n_11640;
wire n_13688;
wire n_4964;
wire n_10180;
wire n_9153;
wire n_6842;
wire n_4700;
wire n_10079;
wire n_7361;
wire n_14825;
wire n_11656;
wire n_4679;
wire n_6397;
wire n_6827;
wire n_11845;
wire n_11679;
wire n_14007;
wire n_13671;
wire n_15839;
wire n_8653;
wire n_5495;
wire n_6281;
wire n_13005;
wire n_4483;
wire n_13313;
wire n_15884;
wire n_5547;
wire n_4693;
wire n_10361;
wire n_15708;
wire n_14154;
wire n_11635;
wire n_8601;
wire n_9675;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_8333;
wire n_9097;
wire n_9571;
wire n_12323;
wire n_12835;
wire n_7079;
wire n_5379;
wire n_15703;
wire n_4487;
wire n_5878;
wire n_10075;
wire n_11572;
wire n_9789;
wire n_13387;
wire n_5820;
wire n_13068;
wire n_11529;
wire n_9925;
wire n_7309;
wire n_7119;
wire n_15139;
wire n_14426;
wire n_7184;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4501;
wire n_4808;
wire n_13173;
wire n_10012;
wire n_14351;
wire n_14957;
wire n_12873;
wire n_12830;
wire n_12015;
wire n_12348;
wire n_12767;
wire n_10939;
wire n_10008;
wire n_11384;
wire n_14382;
wire n_9511;
wire n_15992;
wire n_9795;
wire n_11134;
wire n_8708;
wire n_10503;
wire n_5964;
wire n_6076;
wire n_10111;
wire n_10982;
wire n_10798;
wire n_11630;
wire n_4678;
wire n_12867;
wire n_13479;
wire n_13710;
wire n_5301;
wire n_13263;
wire n_13203;
wire n_14700;
wire n_5126;
wire n_13211;
wire n_8659;
wire n_15469;
wire n_6732;
wire n_8759;
wire n_9622;
wire n_12198;
wire n_9761;
wire n_14707;
wire n_6817;
wire n_5776;
wire n_15408;
wire n_7646;
wire n_14249;
wire n_9954;
wire n_14530;
wire n_14870;
wire n_13848;
wire n_6982;
wire n_12617;
wire n_15184;
wire n_7291;
wire n_10669;
wire n_8790;
wire n_13052;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_8832;
wire n_13282;
wire n_8305;
wire n_14999;
wire n_4303;
wire n_5603;
wire n_8453;
wire n_15800;
wire n_6560;
wire n_6634;
wire n_14275;
wire n_5348;
wire n_12666;
wire n_9847;
wire n_13818;
wire n_4868;
wire n_7017;
wire n_13846;
wire n_12845;
wire n_15961;
wire n_11617;
wire n_7848;
wire n_13312;
wire n_4465;
wire n_14969;
wire n_9640;
wire n_8127;
wire n_13565;
wire n_5217;
wire n_15764;
wire n_8337;
wire n_9115;
wire n_5558;
wire n_7861;
wire n_12047;
wire n_10190;
wire n_12411;
wire n_9534;
wire n_15274;
wire n_13788;
wire n_4245;
wire n_11422;
wire n_5520;
wire n_7889;
wire n_13295;
wire n_12594;
wire n_10542;
wire n_14349;
wire n_5909;
wire n_16127;
wire n_4852;
wire n_7554;
wire n_11289;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_11376;
wire n_5750;
wire n_7648;
wire n_8968;
wire n_10752;
wire n_5654;
wire n_11157;
wire n_16178;
wire n_14718;
wire n_14819;
wire n_10868;
wire n_11013;
wire n_9594;
wire n_11017;
wire n_7653;
wire n_11765;
wire n_6400;
wire n_12885;
wire n_11307;
wire n_7846;
wire n_8347;
wire n_5554;
wire n_9503;
wire n_12811;
wire n_9919;
wire n_15596;
wire n_13346;
wire n_13331;
wire n_5135;
wire n_16071;
wire n_15605;
wire n_7551;
wire n_11793;
wire n_11574;
wire n_4599;
wire n_13307;
wire n_4222;
wire n_6655;
wire n_10017;
wire n_13574;
wire n_12073;
wire n_8093;
wire n_8899;
wire n_9385;
wire n_12913;
wire n_13027;
wire n_14563;
wire n_5448;
wire n_14357;
wire n_15104;
wire n_7737;
wire n_6480;
wire n_5837;
wire n_11836;
wire n_5412;
wire n_8481;
wire n_14169;
wire n_15456;
wire n_15971;
wire n_6851;
wire n_6621;
wire n_11747;
wire n_4701;
wire n_7606;
wire n_9963;
wire n_7420;
wire n_10572;
wire n_11193;
wire n_9885;
wire n_8115;
wire n_4869;
wire n_15914;
wire n_13939;
wire n_5533;
wire n_11670;
wire n_14042;
wire n_10642;
wire n_10115;
wire n_10517;
wire n_14429;
wire n_14098;
wire n_13289;
wire n_10247;
wire n_13851;
wire n_13852;
wire n_5224;
wire n_12451;
wire n_12585;
wire n_12029;
wire n_12963;
wire n_13616;
wire n_6226;
wire n_14490;
wire n_9827;
wire n_12169;
wire n_14748;
wire n_12801;
wire n_9182;
wire n_10620;
wire n_9426;
wire n_8182;
wire n_9293;
wire n_10065;
wire n_15318;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_11762;
wire n_14030;
wire n_14500;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_9581;
wire n_5900;
wire n_8629;
wire n_12657;
wire n_8186;
wire n_7319;
wire n_15721;
wire n_11758;
wire n_15082;
wire n_6158;
wire n_13366;
wire n_9400;
wire n_15028;
wire n_10744;
wire n_9246;
wire n_4342;
wire n_6819;
wire n_6122;
wire n_4903;
wire n_8233;
wire n_4382;
wire n_6898;
wire n_14734;
wire n_14814;
wire n_6570;
wire n_5486;
wire n_9445;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_6843;
wire n_4475;
wire n_5851;
wire n_7516;
wire n_5432;
wire n_14838;
wire n_15620;
wire n_6317;
wire n_6928;
wire n_10609;
wire n_15449;
wire n_13860;
wire n_11958;
wire n_6707;
wire n_10009;
wire n_13847;
wire n_7244;
wire n_11314;
wire n_4626;
wire n_12210;
wire n_10072;
wire n_12443;
wire n_12699;
wire n_7625;
wire n_8750;
wire n_10130;
wire n_4997;
wire n_8183;
wire n_13657;
wire n_5065;
wire n_9104;
wire n_13450;
wire n_6806;
wire n_15752;
wire n_10956;
wire n_7991;
wire n_15389;
wire n_8637;
wire n_9542;
wire n_4638;
wire n_11490;
wire n_11515;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_13610;
wire n_15813;
wire n_6269;
wire n_7857;
wire n_13871;
wire n_7970;
wire n_16021;
wire n_9302;
wire n_8258;
wire n_10829;
wire n_7154;
wire n_11356;
wire n_12781;
wire n_15991;
wire n_10506;
wire n_9960;
wire n_12573;
wire n_13326;
wire n_14843;
wire n_5295;
wire n_8416;
wire n_8390;
wire n_13881;
wire n_11678;
wire n_12744;
wire n_6088;
wire n_10236;
wire n_11374;
wire n_14519;
wire n_11176;
wire n_7194;
wire n_16072;
wire n_4841;
wire n_11402;
wire n_4683;
wire n_5173;
wire n_11162;
wire n_10002;
wire n_8696;
wire n_9185;
wire n_9601;
wire n_13137;
wire n_15698;
wire n_13226;
wire n_11771;
wire n_15951;
wire n_5655;
wire n_5855;
wire n_7175;
wire n_7163;
wire n_13431;
wire n_14402;
wire n_14507;
wire n_14845;
wire n_14020;
wire n_13552;
wire n_13164;
wire n_7027;
wire n_8552;
wire n_12006;
wire n_5861;
wire n_4600;
wire n_6964;
wire n_10855;
wire n_14389;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_9403;
wire n_14558;
wire n_11322;
wire n_6316;
wire n_8619;
wire n_7068;
wire n_11484;
wire n_9972;
wire n_11711;
wire n_13227;
wire n_14541;
wire n_8594;
wire n_9878;
wire n_10139;
wire n_14183;
wire n_9541;
wire n_16055;
wire n_10941;
wire n_14689;
wire n_15667;
wire n_12548;
wire n_8162;
wire n_9735;
wire n_9576;
wire n_14528;
wire n_4549;
wire n_7327;
wire n_16190;
wire n_12727;
wire n_15588;
wire n_12240;
wire n_13045;
wire n_6610;
wire n_13620;
wire n_15919;
wire n_5998;
wire n_8318;
wire n_14742;
wire n_4702;
wire n_5102;
wire n_9974;
wire n_4954;
wire n_15707;
wire n_10992;
wire n_4491;
wire n_8425;
wire n_6752;
wire n_13001;
wire n_6959;
wire n_9704;
wire n_6250;
wire n_13919;
wire n_11392;
wire n_12372;
wire n_11803;
wire n_15597;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_11912;
wire n_13862;
wire n_15066;
wire n_13784;
wire n_7864;
wire n_11139;
wire n_10650;
wire n_8051;
wire n_4734;
wire n_11021;
wire n_6675;
wire n_7955;
wire n_15204;
wire n_5827;
wire n_9039;
wire n_12914;
wire n_16141;
wire n_7384;
wire n_12844;
wire n_5656;
wire n_7218;
wire n_12952;
wire n_15996;
wire n_5678;
wire n_6561;
wire n_11379;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_13271;
wire n_7512;
wire n_7814;
wire n_12276;
wire n_12096;
wire n_8389;
wire n_4515;
wire n_10417;
wire n_10029;
wire n_12150;
wire n_14271;
wire n_13595;
wire n_8620;
wire n_10125;
wire n_5555;
wire n_13757;
wire n_15711;
wire n_8886;
wire n_7152;
wire n_4809;
wire n_14770;
wire n_10253;
wire n_11899;
wire n_16051;
wire n_15533;
wire n_13761;
wire n_15705;
wire n_15574;
wire n_5212;
wire n_4760;
wire n_13190;
wire n_13136;
wire n_6823;
wire n_10693;
wire n_14461;
wire n_7062;
wire n_7090;
wire n_12449;
wire n_8202;
wire n_15261;
wire n_13633;
wire n_11966;
wire n_14205;
wire n_5815;
wire n_4320;
wire n_12118;
wire n_10599;
wire n_5084;
wire n_7223;
wire n_14266;
wire n_12770;
wire n_5251;
wire n_15014;
wire n_8755;
wire n_13174;
wire n_16028;
wire n_8668;
wire n_5965;
wire n_4980;
wire n_10977;
wire n_13528;
wire n_6796;
wire n_8979;
wire n_5407;
wire n_12814;
wire n_11553;
wire n_4560;
wire n_14064;
wire n_14322;
wire n_13220;
wire n_12009;
wire n_15550;
wire n_13456;
wire n_13916;
wire n_7761;
wire n_10947;
wire n_8141;
wire n_10386;
wire n_8199;
wire n_5042;
wire n_12826;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_10267;
wire n_6090;
wire n_5368;
wire n_10401;
wire n_15666;
wire n_15511;
wire n_16160;
wire n_15171;
wire n_15933;
wire n_9908;
wire n_11127;
wire n_11926;
wire n_8004;
wire n_8383;
wire n_14763;
wire n_9688;
wire n_9864;
wire n_12144;
wire n_7388;
wire n_7056;
wire n_10428;
wire n_14585;
wire n_10212;
wire n_7437;
wire n_11460;
wire n_6489;
wire n_11486;
wire n_9023;
wire n_5310;
wire n_8895;
wire n_8680;
wire n_14208;
wire n_6714;
wire n_4987;
wire n_8394;
wire n_7849;
wire n_10539;
wire n_14152;
wire n_7726;
wire n_4572;
wire n_7417;
wire n_12937;
wire n_11148;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_10728;
wire n_12312;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_6791;
wire n_6620;
wire n_4540;
wire n_9220;
wire n_13929;
wire n_6821;
wire n_9317;
wire n_12580;
wire n_13965;
wire n_13796;
wire n_5588;
wire n_8198;
wire n_9993;
wire n_10879;
wire n_13474;
wire n_8665;
wire n_12393;
wire n_16168;
wire n_6583;
wire n_10545;
wire n_12201;
wire n_7859;
wire n_13240;
wire n_13187;
wire n_13594;
wire n_4854;
wire n_9561;
wire n_10516;
wire n_14640;
wire n_9444;
wire n_10497;
wire n_8017;
wire n_16131;
wire n_11675;
wire n_5477;
wire n_10705;
wire n_7523;
wire n_12082;
wire n_13966;
wire n_14936;
wire n_11032;
wire n_5234;
wire n_14035;
wire n_12322;
wire n_6890;
wire n_9184;
wire n_10432;
wire n_11454;
wire n_7559;
wire n_14345;
wire n_9037;
wire n_7576;
wire n_6988;
wire n_8303;
wire n_10779;
wire n_11554;
wire n_5871;
wire n_11988;
wire n_13981;
wire n_4747;
wire n_14647;
wire n_16162;
wire n_8000;
wire n_11197;
wire n_14286;
wire n_14686;
wire n_6052;
wire n_7769;
wire n_15172;
wire n_15305;
wire n_11416;
wire n_9505;
wire n_9193;
wire n_14360;
wire n_7257;
wire n_12986;
wire n_15179;
wire n_6973;
wire n_10869;
wire n_8852;
wire n_5007;
wire n_8709;
wire n_4881;
wire n_10314;
wire n_10504;
wire n_6488;
wire n_4495;
wire n_10687;
wire n_13691;
wire n_4737;
wire n_9218;
wire n_9755;
wire n_4357;
wire n_11341;
wire n_7729;
wire n_4502;
wire n_11045;
wire n_12373;
wire n_7005;
wire n_12741;
wire n_5334;
wire n_15544;
wire n_8782;
wire n_7081;
wire n_10882;
wire n_7742;
wire n_5253;
wire n_10293;
wire n_6280;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_14828;
wire n_15152;
wire n_9162;
wire n_9506;
wire n_13629;
wire n_15264;
wire n_15584;
wire n_7341;
wire n_5792;
wire n_13155;
wire n_14581;
wire n_15493;
wire n_4513;
wire n_11569;
wire n_13152;
wire n_10256;
wire n_4775;
wire n_6256;
wire n_8716;
wire n_12412;
wire n_8250;
wire n_7264;
wire n_12677;
wire n_7842;
wire n_15976;
wire n_16142;
wire n_14315;
wire n_12181;
wire n_12833;
wire n_6648;
wire n_9415;
wire n_10298;
wire n_12631;
wire n_12115;
wire n_14829;
wire n_16091;
wire n_7492;
wire n_13194;
wire n_15331;
wire n_13546;
wire n_6649;
wire n_8714;
wire n_8357;
wire n_12567;
wire n_12175;
wire n_15424;
wire n_15791;
wire n_6910;
wire n_9990;
wire n_14920;
wire n_15687;
wire n_8466;
wire n_4264;
wire n_5954;
wire n_9015;
wire n_10326;
wire n_14827;
wire n_13446;
wire n_15482;
wire n_10235;
wire n_4709;
wire n_6431;
wire n_8589;
wire n_12754;
wire n_4223;
wire n_14141;
wire n_12455;
wire n_13363;
wire n_11990;
wire n_8266;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_4718;
wire n_10725;
wire n_6324;
wire n_5489;
wire n_15653;
wire n_10274;
wire n_13728;
wire n_13601;
wire n_8876;
wire n_11541;
wire n_9214;
wire n_14780;
wire n_4206;
wire n_12340;
wire n_10799;
wire n_8922;
wire n_11680;
wire n_10090;
wire n_6512;
wire n_12686;
wire n_5342;
wire n_9070;
wire n_15993;
wire n_8498;
wire n_4794;
wire n_9933;
wire n_4843;
wire n_12734;
wire n_5580;
wire n_15108;
wire n_5215;
wire n_15870;
wire n_12331;
wire n_4763;
wire n_10874;
wire n_9339;
wire n_11596;
wire n_9991;
wire n_12880;
wire n_9486;
wire n_8457;
wire n_6243;
wire n_14113;
wire n_5795;
wire n_10763;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_10266;
wire n_8267;
wire n_12184;
wire n_12425;
wire n_7051;
wire n_13918;
wire n_14997;
wire n_11180;
wire n_6773;
wire n_10290;
wire n_6231;
wire n_15758;
wire n_12472;
wire n_13048;
wire n_12266;
wire n_7503;
wire n_12432;
wire n_4838;
wire n_4795;
wire n_8124;
wire n_8545;
wire n_5430;
wire n_6041;
wire n_8526;
wire n_12300;
wire n_13593;
wire n_8319;
wire n_7997;
wire n_12527;
wire n_5659;
wire n_11839;
wire n_9279;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_10732;
wire n_5195;
wire n_12110;
wire n_15354;
wire n_15310;
wire n_13744;
wire n_9790;
wire n_11404;
wire n_7950;
wire n_11548;
wire n_6323;
wire n_13515;
wire n_5720;
wire n_4267;
wire n_8581;
wire n_12122;
wire n_14889;
wire n_10873;
wire n_16026;
wire n_8214;
wire n_15583;
wire n_7793;
wire n_9053;
wire n_8516;
wire n_12310;
wire n_5598;
wire n_11343;
wire n_8989;
wire n_13028;
wire n_7746;
wire n_11362;
wire n_15941;
wire n_4352;
wire n_11007;
wire n_7570;
wire n_9650;
wire n_16119;
wire n_9880;
wire n_11497;
wire n_15859;
wire n_10720;
wire n_6912;
wire n_14574;
wire n_7425;
wire n_15050;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_14014;
wire n_12827;
wire n_14078;
wire n_10220;
wire n_9217;
wire n_9499;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_15696;
wire n_13467;
wire n_13245;
wire n_6747;
wire n_5303;
wire n_10081;
wire n_12804;
wire n_6916;
wire n_9282;
wire n_7894;
wire n_10145;
wire n_11347;
wire n_7957;
wire n_8262;
wire n_10167;
wire n_5530;
wire n_12892;
wire n_12656;
wire n_6718;
wire n_8289;
wire n_13804;
wire n_5809;
wire n_10447;
wire n_12418;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_12448;
wire n_15180;
wire n_12219;
wire n_12729;
wire n_13549;
wire n_13921;
wire n_6473;
wire n_8087;
wire n_10238;
wire n_13345;
wire n_4806;
wire n_11029;
wire n_7961;
wire n_9920;
wire n_5993;
wire n_15129;
wire n_6574;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_9948;
wire n_5299;
wire n_4462;
wire n_13216;
wire n_4219;
wire n_4723;
wire n_4484;
wire n_11226;
wire n_8863;
wire n_9371;
wire n_15396;
wire n_4517;
wire n_8701;
wire n_15551;
wire n_13036;
wire n_15603;
wire n_9237;
wire n_15038;
wire n_13398;
wire n_6857;
wire n_8705;
wire n_14148;
wire n_9815;
wire n_10292;
wire n_12644;
wire n_6975;
wire n_15413;
wire n_10820;
wire n_7763;
wire n_13258;
wire n_6290;
wire n_6646;
wire n_7703;
wire n_11760;
wire n_15781;
wire n_13827;
wire n_7928;
wire n_4234;
wire n_10395;
wire n_12576;
wire n_10168;
wire n_14350;
wire n_8722;
wire n_11664;
wire n_5821;
wire n_15306;
wire n_6622;
wire n_12187;
wire n_7665;
wire n_4836;
wire n_5522;
wire n_7677;
wire n_5262;
wire n_13169;
wire n_14782;
wire n_15978;
wire n_10366;
wire n_5319;
wire n_10287;
wire n_14017;
wire n_15358;
wire n_13940;
wire n_7469;
wire n_10163;
wire n_6118;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_14145;
wire n_11006;
wire n_6532;
wire n_13406;
wire n_10431;
wire n_8622;
wire n_8099;
wire n_8729;
wire n_9479;
wire n_10876;
wire n_11485;
wire n_15092;
wire n_6267;
wire n_15397;
wire n_6682;
wire n_9480;
wire n_12453;
wire n_12593;
wire n_4207;
wire n_11449;
wire n_8085;
wire n_15984;
wire n_4725;
wire n_9597;
wire n_10614;
wire n_10786;
wire n_13873;
wire n_13335;
wire n_14273;
wire n_9173;
wire n_10352;
wire n_15458;
wire n_16067;
wire n_7203;
wire n_8947;
wire n_9641;
wire n_13714;
wire n_7797;
wire n_9983;
wire n_9267;
wire n_14565;
wire n_5943;
wire n_6556;
wire n_10039;
wire n_15079;
wire n_4880;
wire n_15784;
wire n_13070;
wire n_6216;
wire n_13866;
wire n_4563;
wire n_7128;
wire n_9849;
wire n_15231;
wire n_11831;
wire n_15454;
wire n_5335;
wire n_6365;
wire n_8459;
wire n_7111;
wire n_11096;
wire n_4334;
wire n_8478;
wire n_5284;
wire n_12288;
wire n_8786;
wire n_9414;
wire n_4978;
wire n_11677;
wire n_13025;
wire n_14256;
wire n_5771;
wire n_9419;
wire n_8887;
wire n_12091;
wire n_14922;
wire n_11898;
wire n_4707;
wire n_14749;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_15168;
wire n_15716;
wire n_8540;
wire n_8276;
wire n_7284;
wire n_5516;
wire n_7057;
wire n_14862;
wire n_13457;
wire n_9823;
wire n_5168;
wire n_9152;
wire n_15915;
wire n_8706;
wire n_6167;
wire n_12357;
wire n_4274;
wire n_5583;
wire n_11826;
wire n_7064;
wire n_12629;
wire n_8532;
wire n_9533;
wire n_10750;
wire n_5433;
wire n_11825;
wire n_7278;
wire n_5429;
wire n_12893;
wire n_9281;
wire n_9103;
wire n_9111;
wire n_6772;
wire n_15499;
wire n_7088;
wire n_7799;
wire n_9618;
wire n_10383;
wire n_16134;
wire n_5698;
wire n_10856;
wire n_5731;
wire n_14532;
wire n_14105;
wire n_10883;
wire n_12935;
wire n_8871;
wire n_8433;
wire n_9065;
wire n_10429;
wire n_14627;
wire n_15552;
wire n_14463;
wire n_15727;
wire n_14735;
wire n_15808;
wire n_15103;
wire n_6159;
wire n_12732;
wire n_5857;
wire n_7048;
wire n_7979;
wire n_12569;
wire n_9674;
wire n_6617;
wire n_7725;
wire n_13547;
wire n_10859;
wire n_5120;
wire n_8371;
wire n_8547;
wire n_11538;
wire n_10815;
wire n_11008;
wire n_8467;
wire n_12980;
wire n_11093;
wire n_11585;
wire n_16205;
wire n_8409;
wire n_6217;
wire n_11616;
wire n_10303;
wire n_9157;
wire n_5560;
wire n_16093;
wire n_15071;
wire n_14831;
wire n_9170;
wire n_4441;
wire n_10424;
wire n_6777;
wire n_5455;
wire n_11001;
wire n_8640;
wire n_15500;
wire n_10196;
wire n_6742;
wire n_15543;
wire n_14823;
wire n_7447;
wire n_5209;
wire n_15807;
wire n_10684;
wire n_13154;
wire n_6307;
wire n_5704;
wire n_14129;
wire n_16074;
wire n_4458;
wire n_4889;
wire n_8431;
wire n_16049;
wire n_14547;
wire n_4523;
wire n_13280;
wire n_5916;
wire n_8415;
wire n_10184;
wire n_13904;
wire n_10421;
wire n_13944;
wire n_15935;
wire n_13359;
wire n_6479;
wire n_11472;
wire n_14376;
wire n_13855;
wire n_13073;
wire n_5099;
wire n_11063;
wire n_5781;
wire n_11179;
wire n_5619;
wire n_14777;
wire n_9416;
wire n_11885;
wire n_9368;
wire n_7365;
wire n_8329;
wire n_13083;
wire n_14201;
wire n_7792;
wire n_9208;
wire n_8089;
wire n_5022;
wire n_11657;
wire n_13124;
wire n_6370;
wire n_9223;
wire n_13771;
wire n_10329;
wire n_10924;
wire n_13845;
wire n_11921;
wire n_15443;
wire n_14224;
wire n_10285;
wire n_7275;
wire n_15039;
wire n_5353;
wire n_4771;
wire n_12099;
wire n_14991;
wire n_6856;
wire n_9781;
wire n_13609;
wire n_13572;
wire n_13817;
wire n_8633;
wire n_12897;
wire n_9392;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_9422;
wire n_15338;
wire n_8541;
wire n_10084;
wire n_12924;
wire n_8762;
wire n_15866;
wire n_14162;
wire n_12619;
wire n_12541;
wire n_5518;
wire n_9970;
wire n_14882;
wire n_13428;
wire n_15880;
wire n_4261;
wire n_15488;
wire n_15508;
wire n_7037;
wire n_13104;
wire n_15292;
wire n_9338;
wire n_15176;
wire n_11647;
wire n_8125;
wire n_6240;
wire n_15222;
wire n_5236;
wire n_4236;
wire n_10077;
wire n_10964;
wire n_14367;
wire n_9492;
wire n_14566;
wire n_6693;
wire n_15694;
wire n_10759;
wire n_9226;
wire n_6712;
wire n_7530;
wire n_10129;
wire n_10101;
wire n_13844;
wire n_11757;
wire n_10566;
wire n_7471;
wire n_9328;
wire n_6465;
wire n_8188;
wire n_10192;
wire n_5673;
wire n_14363;
wire n_11846;
wire n_11519;
wire n_14571;
wire n_8615;
wire n_5814;
wire n_6586;
wire n_7058;
wire n_14857;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_12191;
wire n_10207;
wire n_6730;
wire n_11530;
wire n_13526;
wire n_13998;
wire n_6367;
wire n_8923;
wire n_11488;
wire n_11389;
wire n_8624;
wire n_8222;
wire n_11928;
wire n_15150;
wire n_12429;
wire n_12825;
wire n_6069;
wire n_6515;
wire n_8206;
wire n_15547;
wire n_15907;
wire n_6077;
wire n_9513;
wire n_11315;
wire n_9393;
wire n_13267;
wire n_15249;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_13506;
wire n_8065;
wire n_9914;
wire n_14833;
wire n_14398;
wire n_7008;
wire n_12318;
wire n_12918;
wire n_14731;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_7540;
wire n_10886;
wire n_12923;
wire n_15112;
wire n_13632;
wire n_14600;
wire n_10804;
wire n_7581;
wire n_12077;
wire n_15132;
wire n_10362;
wire n_7139;
wire n_10437;
wire n_10384;
wire n_13834;
wire n_8935;
wire n_14213;
wire n_15081;
wire n_16158;
wire n_16044;
wire n_13444;
wire n_10885;
wire n_11962;
wire n_11002;
wire n_5239;
wire n_13885;
wire n_12805;
wire n_14928;
wire n_7782;
wire n_7432;
wire n_4913;
wire n_13067;
wire n_8155;
wire n_9334;
wire n_14059;
wire n_11648;
wire n_10093;
wire n_13924;
wire n_14289;
wire n_4428;
wire n_12808;
wire n_6483;
wire n_7770;
wire n_12853;
wire n_9684;
wire n_12591;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_10600;
wire n_10480;
wire n_11994;
wire n_8175;
wire n_5357;
wire n_7173;
wire n_10892;
wire n_9254;
wire n_6576;
wire n_6810;
wire n_10003;
wire n_11050;
wire n_5421;
wire n_9083;
wire n_11250;
wire n_12645;
wire n_16106;
wire n_11316;
wire n_14727;
wire n_14485;
wire n_15277;
wire n_12987;
wire n_4396;
wire n_15938;
wire n_13717;
wire n_6708;
wire n_12251;
wire n_10252;
wire n_16229;
wire n_12948;
wire n_8026;
wire n_6667;
wire n_9175;
wire n_9838;
wire n_15636;
wire n_11428;
wire n_12467;
wire n_12756;
wire n_11463;
wire n_15280;
wire n_6040;
wire n_10495;
wire n_6847;
wire n_8974;
wire n_6305;
wire n_8836;
wire n_10812;
wire n_12678;
wire n_14211;
wire n_4228;
wire n_14641;
wire n_12700;
wire n_11674;
wire n_11097;
wire n_11069;
wire n_7251;
wire n_10894;
wire n_12602;
wire n_14155;
wire n_12194;
wire n_15751;
wire n_7356;
wire n_7412;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_15465;
wire n_11318;
wire n_7751;
wire n_12351;
wire n_7951;
wire n_12965;
wire n_7060;
wire n_14184;
wire n_9336;
wire n_12367;
wire n_13603;
wire n_8873;
wire n_14111;
wire n_10311;
wire n_7591;
wire n_10490;
wire n_6750;
wire n_5769;
wire n_7444;
wire n_10702;
wire n_15207;
wire n_7911;
wire n_7595;
wire n_4931;
wire n_7790;
wire n_11586;
wire n_7426;
wire n_11786;
wire n_13571;
wire n_4400;
wire n_7502;
wire n_13492;
wire n_5434;
wire n_10906;
wire n_10891;
wire n_6855;
wire n_10840;
wire n_8170;
wire n_14257;
wire n_15019;
wire n_5181;
wire n_6239;
wire n_10181;
wire n_13673;
wire n_12036;
wire n_9554;
wire n_14589;
wire n_15950;
wire n_5768;
wire n_11330;
wire n_6199;
wire n_12263;
wire n_8120;
wire n_9116;
wire n_9315;
wire n_9830;
wire n_8825;
wire n_14416;
wire n_9169;
wire n_7252;
wire n_11201;
wire n_5963;
wire n_9999;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_14899;
wire n_12703;
wire n_4192;
wire n_8003;
wire n_11979;
wire n_12253;
wire n_9215;
wire n_15380;
wire n_6789;
wire n_5972;
wire n_8395;
wire n_13986;
wire n_7065;
wire n_8083;
wire n_14963;
wire n_11888;
wire n_6177;
wire n_14596;
wire n_8057;
wire n_5937;
wire n_15902;
wire n_9259;
wire n_5146;
wire n_7367;
wire n_10755;
wire n_14274;
wire n_11835;
wire n_11537;
wire n_8164;
wire n_10525;
wire n_11583;
wire n_12776;
wire n_14714;
wire n_15897;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_15069;
wire n_4221;
wire n_12445;
wire n_8877;
wire n_6825;
wire n_15282;
wire n_7614;
wire n_6460;
wire n_9150;
wire n_6952;
wire n_9595;
wire n_11420;
wire n_8366;
wire n_14907;
wire n_6173;
wire n_8476;
wire n_4190;
wire n_11527;
wire n_6218;
wire n_10435;
wire n_10342;
wire n_11048;
wire n_7685;
wire n_14584;
wire n_11933;
wire n_6486;
wire n_15133;
wire n_13826;
wire n_11900;
wire n_12620;
wire n_7619;
wire n_11106;
wire n_15237;
wire n_15832;
wire n_12299;
wire n_13078;
wire n_5013;
wire n_4145;
wire n_10983;
wire n_11266;
wire n_6852;
wire n_11340;
wire n_11929;
wire n_15659;
wire n_15709;
wire n_5577;
wire n_12673;
wire n_13557;
wire n_9100;
wire n_5872;
wire n_7883;
wire n_13516;
wire n_10397;
wire n_15007;
wire n_6692;
wire n_15337;
wire n_13208;
wire n_9707;
wire n_5017;
wire n_16010;
wire n_8854;
wire n_13523;
wire n_12834;
wire n_10202;
wire n_14549;
wire n_12821;
wire n_10677;
wire n_7220;
wire n_7560;
wire n_10648;
wire n_9262;
wire n_5976;
wire n_4717;
wire n_9249;
wire n_6888;
wire n_4739;
wire n_14798;
wire n_11964;
wire n_12247;
wire n_15023;
wire n_13030;
wire n_8256;
wire n_4312;
wire n_5424;
wire n_13065;
wire n_7270;
wire n_14751;
wire n_10273;
wire n_12927;
wire n_12324;
wire n_12817;
wire n_15627;
wire n_11255;
wire n_8621;
wire n_13753;
wire n_11751;
wire n_4750;
wire n_10978;
wire n_9806;
wire n_10834;
wire n_13430;
wire n_8577;
wire n_9019;
wire n_10097;
wire n_13880;
wire n_14796;
wire n_9361;
wire n_7731;
wire n_6626;
wire n_13175;
wire n_4537;
wire n_13050;
wire n_10890;
wire n_5838;
wire n_13732;
wire n_7034;
wire n_10816;
wire n_8654;
wire n_12887;
wire n_13133;
wire n_6854;
wire n_7940;
wire n_15496;
wire n_16256;
wire n_6793;
wire n_14188;
wire n_5456;
wire n_4847;
wire n_5846;
wire n_9814;
wire n_11930;
wire n_15361;
wire n_5930;
wire n_11269;
wire n_10462;
wire n_12316;
wire n_12539;
wire n_13358;
wire n_8952;
wire n_13823;
wire n_12758;
wire n_12414;
wire n_9438;
wire n_7537;
wire n_12600;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_14875;
wire n_15920;
wire n_15506;
wire n_11985;
wire n_4427;
wire n_7458;
wire n_7740;
wire n_4705;
wire n_15572;
wire n_15149;
wire n_6794;
wire n_12949;
wire n_11205;
wire n_9856;
wire n_8421;
wire n_7179;
wire n_10832;
wire n_7433;
wire n_13499;
wire n_14057;
wire n_4279;
wire n_9327;
wire n_9313;
wire n_4330;
wire n_6334;
wire n_13560;
wire n_6257;
wire n_16219;
wire n_10142;
wire n_4152;
wire n_6874;
wire n_14073;
wire n_14079;
wire n_10300;
wire n_15489;
wire n_8911;
wire n_15340;
wire n_5537;
wire n_9518;
wire n_5572;
wire n_15693;
wire n_4783;
wire n_7658;
wire n_10335;
wire n_10753;
wire n_5409;
wire n_14220;
wire n_15783;
wire n_4539;
wire n_12783;
wire n_13658;
wire n_5142;
wire n_12431;
wire n_10921;
wire n_10177;
wire n_8971;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_10567;
wire n_6286;
wire n_4603;
wire n_5010;
wire n_15677;
wire n_4332;
wire n_7226;
wire n_11915;
wire n_7987;
wire n_9291;
wire n_7217;
wire n_9009;
wire n_9882;
wire n_6377;
wire n_10492;
wire n_14137;
wire n_15385;
wire n_12061;
wire n_5401;
wire n_16176;
wire n_4595;
wire n_7272;
wire n_11873;
wire n_15505;
wire n_8215;
wire n_16048;
wire n_5201;
wire n_5816;
wire n_12628;
wire n_5551;
wire n_9722;
wire n_5416;
wire n_14175;
wire n_4404;
wire n_15373;
wire n_14644;
wire n_7906;
wire n_11260;
wire n_5498;
wire n_16172;
wire n_5543;
wire n_12359;
wire n_15328;
wire n_9760;
wire n_6018;
wire n_7765;
wire n_14320;
wire n_6021;
wire n_11880;
wire n_11605;
wire n_13615;
wire n_4617;
wire n_14022;
wire n_12974;
wire n_13156;
wire n_10741;
wire n_4611;
wire n_10037;
wire n_8949;
wire n_12136;
wire n_5797;
wire n_9454;
wire n_10760;
wire n_6511;
wire n_13849;
wire n_12121;
wire n_7815;
wire n_12658;
wire n_11838;
wire n_13956;
wire n_4732;
wire n_14768;
wire n_10607;
wire n_5942;
wire n_5764;
wire n_13702;
wire n_8983;
wire n_4969;
wire n_11089;
wire n_14314;
wire n_8121;
wire n_15088;
wire n_5252;
wire n_11629;
wire n_11259;
wire n_5777;
wire n_11100;
wire n_15283;
wire n_13119;
wire n_8942;
wire n_7785;
wire n_11608;
wire n_13756;
wire n_4641;
wire n_5063;
wire n_15564;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_12364;
wire n_14628;
wire n_13867;
wire n_8280;
wire n_7728;
wire n_11632;
wire n_16094;
wire n_4712;
wire n_7255;
wire n_7181;
wire n_12156;
wire n_11443;
wire n_13409;
wire n_13832;
wire n_5393;
wire n_10658;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_8427;
wire n_11161;
wire n_11770;
wire n_13509;
wire n_14399;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_6322;
wire n_7359;
wire n_5643;
wire n_11466;
wire n_15931;
wire n_10489;
wire n_15270;
wire n_9826;
wire n_9937;
wire n_10347;
wire n_12632;
wire n_11810;
wire n_7825;
wire n_13168;
wire n_4437;
wire n_6419;
wire n_7916;
wire n_16170;
wire n_13581;
wire n_10952;
wire n_8194;
wire n_15862;
wire n_10758;
wire n_15798;
wire n_5346;
wire n_7283;
wire n_9453;
wire n_7903;
wire n_9900;
wire n_12033;
wire n_7089;
wire n_16128;
wire n_14954;
wire n_8217;
wire n_14534;
wire n_14890;
wire n_10518;
wire n_9331;
wire n_7604;
wire n_11789;
wire n_7647;
wire n_13447;
wire n_12465;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_15649;
wire n_14164;
wire n_14771;
wire n_5868;
wire n_6417;
wire n_8521;
wire n_8285;
wire n_7145;
wire n_10808;
wire n_12358;
wire n_4867;
wire n_12446;
wire n_9178;
wire n_7803;
wire n_9689;
wire n_13999;
wire n_8448;
wire n_14526;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_11690;
wire n_5986;
wire n_12684;
wire n_9355;
wire n_12851;
wire n_13725;
wire n_16206;
wire n_9489;
wire n_13319;
wire n_6932;
wire n_12307;
wire n_10971;
wire n_15757;
wire n_7258;
wire n_13019;
wire n_5104;
wire n_16236;
wire n_12341;
wire n_13807;
wire n_6961;
wire n_8732;
wire n_13297;
wire n_7622;
wire n_14610;
wire n_11968;
wire n_9359;
wire n_13395;
wire n_7839;
wire n_11854;
wire n_6792;
wire n_7720;
wire n_4368;
wire n_16152;
wire n_5794;
wire n_8136;
wire n_10404;
wire n_5272;
wire n_6919;
wire n_11797;
wire n_8420;
wire n_13672;
wire n_4430;
wire n_8386;
wire n_16097;
wire n_6123;
wire n_5338;
wire n_10802;
wire n_7440;
wire n_15317;
wire n_9568;
wire n_6831;
wire n_4544;
wire n_14302;
wire n_5578;
wire n_12654;
wire n_4191;
wire n_4409;
wire n_12921;
wire n_11991;
wire n_7809;
wire n_16140;
wire n_10340;
wire n_5722;
wire n_16043;
wire n_5811;
wire n_14170;
wire n_7072;
wire n_10681;
wire n_14303;
wire n_15077;
wire n_4961;
wire n_11618;
wire n_15202;
wire n_11502;
wire n_10452;
wire n_10221;
wire n_8746;
wire n_10051;
wire n_5395;
wire n_4531;
wire n_12498;
wire n_6458;
wire n_11465;
wire n_12768;
wire n_9401;
wire n_8857;
wire n_11335;
wire n_6986;
wire n_9495;
wire n_12625;
wire n_13221;
wire n_10987;
wire n_4532;
wire n_15409;
wire n_10551;
wire n_7564;
wire n_12063;
wire n_10396;
wire n_10646;
wire n_13471;
wire n_13021;
wire n_15589;
wire n_15322;
wire n_10955;
wire n_5863;
wire n_8185;
wire n_8313;
wire n_6633;
wire n_11382;
wire n_13062;
wire n_14298;
wire n_14931;
wire n_7775;
wire n_7118;
wire n_9234;
wire n_7960;
wire n_14967;
wire n_6152;
wire n_9431;
wire n_5734;
wire n_15831;
wire n_10308;
wire n_10023;
wire n_8281;
wire n_12347;
wire n_12543;
wire n_12958;
wire n_11254;
wire n_5095;
wire n_14797;
wire n_10538;
wire n_6169;
wire n_5774;
wire n_12532;
wire n_15974;
wire n_7069;
wire n_11388;
wire n_5199;
wire n_13347;
wire n_6546;
wire n_15557;
wire n_14051;
wire n_4257;
wire n_15548;
wire n_4282;
wire n_11043;
wire n_7636;
wire n_4341;
wire n_10199;
wire n_6925;
wire n_10673;
wire n_7186;
wire n_10467;
wire n_8766;
wire n_13976;
wire n_12334;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_12876;
wire n_4944;
wire n_8066;
wire n_11252;
wire n_9340;
wire n_12774;
wire n_12544;
wire n_13793;
wire n_9380;
wire n_7666;
wire n_15892;
wire n_12353;
wire n_6425;
wire n_12653;
wire n_11824;
wire n_10581;
wire n_14594;
wire n_15816;
wire n_14369;
wire n_9976;
wire n_4994;
wire n_10818;
wire n_10226;
wire n_7967;
wire n_5977;
wire n_14515;
wire n_16052;
wire n_15998;
wire n_8314;
wire n_5175;
wire n_7246;
wire n_11724;
wire n_12052;
wire n_11507;
wire n_11086;
wire n_10647;
wire n_13184;
wire n_9064;
wire n_15311;
wire n_4381;
wire n_8239;
wire n_9092;
wire n_14968;
wire n_14721;
wire n_11533;
wire n_4316;
wire n_15900;
wire n_7301;
wire n_11905;
wire n_14160;
wire n_4860;
wire n_4469;
wire n_16017;
wire n_9746;
wire n_12994;
wire n_4930;
wire n_8497;
wire n_5352;
wire n_10637;
wire n_15824;
wire n_7262;
wire n_5959;
wire n_15089;
wire n_13856;
wire n_8056;
wire n_8210;
wire n_10769;
wire n_5945;
wire n_4423;
wire n_12215;
wire n_10519;
wire n_13218;
wire n_7584;
wire n_7748;
wire n_9066;
wire n_14637;
wire n_6301;
wire n_14965;
wire n_15988;
wire n_13298;
wire n_5668;
wire n_12535;
wire n_14248;
wire n_4209;
wire n_12582;
wire n_15175;
wire n_14982;
wire n_7686;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_11800;
wire n_9870;
wire n_14391;
wire n_9817;
wire n_12505;
wire n_13396;
wire n_13988;
wire n_14648;
wire n_7059;
wire n_15349;
wire n_14947;
wire n_15725;
wire n_6985;
wire n_4350;
wire n_5600;
wire n_13132;
wire n_15546;
wire n_6737;
wire n_10723;
wire n_12875;
wire n_9857;
wire n_13794;
wire n_4804;
wire n_8404;
wire n_4888;
wire n_5767;
wire n_9455;
wire n_10056;
wire n_6459;
wire n_15126;
wire n_7670;
wire n_13400;
wire n_13813;
wire n_14307;
wire n_4936;
wire n_8505;
wire n_10653;
wire n_6384;
wire n_4669;
wire n_15345;
wire n_15509;
wire n_5228;
wire n_15571;
wire n_15678;
wire n_15777;
wire n_9916;
wire n_10157;
wire n_8606;
wire n_13542;
wire n_7443;
wire n_10701;
wire n_10470;
wire n_10923;
wire n_12828;
wire n_5973;
wire n_7484;
wire n_12402;
wire n_14387;
wire n_9440;
wire n_4759;
wire n_10038;
wire n_9059;
wire n_11691;
wire n_9812;
wire n_14666;
wire n_5869;
wire n_5914;
wire n_6753;
wire n_9690;
wire n_13879;
wire n_11594;
wire n_9912;
wire n_11687;
wire n_14793;
wire n_4887;
wire n_15913;
wire n_9002;
wire n_11513;
wire n_16057;
wire n_9620;
wire n_10619;
wire n_13522;
wire n_6448;
wire n_9229;
wire n_12524;
wire n_14535;
wire n_15051;
wire n_5186;
wire n_14196;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_13403;
wire n_10454;
wire n_11655;
wire n_13241;
wire n_4218;
wire n_9464;
wire n_11386;
wire n_4687;
wire n_7077;
wire n_14060;
wire n_10656;
wire n_10871;
wire n_15406;
wire n_8518;
wire n_11111;
wire n_13270;
wire n_4720;
wire n_15037;
wire n_11938;
wire n_6043;
wire n_6268;
wire n_12670;
wire n_9497;
wire n_14923;
wire n_14543;
wire n_5604;
wire n_7663;
wire n_8350;
wire n_8741;
wire n_10444;
wire n_11866;
wire n_7024;
wire n_8148;
wire n_5221;
wire n_11833;
wire n_8408;
wire n_6145;
wire n_12308;
wire n_15523;
wire n_10846;
wire n_12659;
wire n_13934;
wire n_14854;
wire n_13024;
wire n_5925;
wire n_6529;
wire n_5591;
wire n_4762;
wire n_13223;
wire n_8236;
wire n_14202;
wire n_11192;
wire n_15970;
wire n_11229;
wire n_7214;
wire n_11244;
wire n_8806;
wire n_14352;
wire n_4490;
wire n_8295;
wire n_9587;
wire n_13888;
wire n_7977;
wire n_15370;
wire n_15166;
wire n_14719;
wire n_15260;
wire n_5387;
wire n_13529;
wire n_12452;
wire n_6311;
wire n_8167;
wire n_11848;
wire n_8377;
wire n_13530;
wire n_7652;
wire n_13591;
wire n_10558;
wire n_9783;
wire n_4644;
wire n_8956;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_7566;
wire n_14631;
wire n_4131;
wire n_11876;
wire n_16120;
wire n_12667;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_15032;
wire n_15121;
wire n_12707;
wire n_6134;
wire n_16246;
wire n_4158;
wire n_6812;
wire n_10466;
wire n_14824;
wire n_10546;
wire n_10044;
wire n_12878;
wire n_14919;
wire n_5190;
wire n_15886;
wire n_6733;
wire n_11666;
wire n_5325;
wire n_13354;
wire n_10527;
wire n_4231;
wire n_8960;
wire n_8957;
wire n_9008;
wire n_10143;
wire n_12361;
wire n_5047;
wire n_5004;
wire n_10233;
wire n_14856;
wire n_6262;
wire n_4926;
wire n_8207;
wire n_6938;
wire n_4872;
wire n_12709;
wire n_4778;
wire n_5876;
wire n_10461;
wire n_5344;
wire n_15827;
wire n_10186;
wire n_6160;
wire n_12721;
wire n_4667;
wire n_5813;
wire n_10113;
wire n_6235;
wire n_13023;
wire n_6212;
wire n_16150;
wire n_9381;
wire n_9194;
wire n_6816;
wire n_8904;
wire n_12264;
wire n_14683;
wire n_7374;
wire n_12464;
wire n_13268;
wire n_12753;
wire n_13887;
wire n_12968;
wire n_15107;
wire n_10120;
wire n_5892;
wire n_9549;
wire n_7678;
wire n_15402;
wire n_4837;
wire n_14848;
wire n_4210;
wire n_15539;
wire n_11248;
wire n_13660;
wire n_7110;
wire n_15712;
wire n_5714;
wire n_12111;
wire n_6953;
wire n_9652;
wire n_7975;
wire n_9957;
wire n_13481;
wire n_15485;
wire n_12609;
wire n_13143;
wire n_12482;
wire n_8451;
wire n_6089;
wire n_10591;
wire n_11780;
wire n_5634;
wire n_12966;
wire n_5133;
wire n_14607;
wire n_7553;
wire n_8527;
wire n_5990;
wire n_7086;
wire n_7732;
wire n_5305;
wire n_5689;
wire n_7891;
wire n_13383;
wire n_13419;
wire n_9089;
wire n_4578;
wire n_8840;
wire n_11424;
wire n_11467;
wire n_5644;
wire n_9137;
wire n_9390;
wire n_11995;
wire n_12178;
wire n_8038;
wire n_8190;
wire n_9439;
wire n_11701;
wire n_15803;
wire n_15405;
wire n_6138;
wire n_15621;
wire n_9080;
wire n_14773;
wire n_15706;
wire n_15878;
wire n_13351;
wire n_9296;
wire n_12997;
wire n_16169;
wire n_10625;
wire n_13544;
wire n_16180;
wire n_4877;
wire n_15060;
wire n_14173;
wire n_9312;
wire n_10662;
wire n_12818;
wire n_9151;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_9883;
wire n_13420;
wire n_14576;
wire n_8287;
wire n_10697;
wire n_14981;
wire n_8111;
wire n_8341;
wire n_13527;
wire n_16006;
wire n_8830;
wire n_13206;
wire n_13235;
wire n_4998;
wire n_10200;
wire n_14436;
wire n_5576;
wire n_13399;
wire n_10935;
wire n_7345;
wire n_9324;
wire n_13317;
wire n_9631;
wire n_8308;
wire n_10547;
wire n_6070;
wire n_15432;
wire n_5852;
wire n_5918;
wire n_8021;
wire n_11092;
wire n_13622;
wire n_10933;
wire n_14790;
wire n_8965;
wire n_9736;
wire n_7041;
wire n_9365;
wire n_10632;
wire n_6717;
wire n_14651;
wire n_16083;
wire n_7593;
wire n_8265;
wire n_13564;
wire n_11166;
wire n_6881;
wire n_10085;
wire n_14881;
wire n_9600;
wire n_6871;
wire n_15629;
wire n_9816;
wire n_6672;
wire n_5343;
wire n_9869;
wire n_7757;
wire n_8251;
wire n_9402;
wire n_7866;
wire n_7334;
wire n_6518;
wire n_13276;
wire n_6396;
wire n_7028;
wire n_14383;
wire n_4379;
wire n_8773;
wire n_12195;
wire n_14400;
wire n_5947;
wire n_6242;
wire n_14143;
wire n_6601;
wire n_8570;
wire n_12536;
wire n_10645;
wire n_10041;
wire n_15392;
wire n_12168;
wire n_14858;
wire n_5835;
wire n_10096;
wire n_12533;
wire n_8579;
wire n_15333;
wire n_15762;
wire n_8079;
wire n_5542;
wire n_9615;
wire n_11869;
wire n_14106;
wire n_5015;
wire n_13792;
wire n_12560;
wire n_5527;
wire n_9759;
wire n_9711;
wire n_4812;
wire n_8506;
wire n_8973;
wire n_13171;
wire n_6606;
wire n_4497;
wire n_13764;
wire n_8291;
wire n_14725;
wire n_4300;
wire n_16077;
wire n_11264;
wire n_10336;
wire n_16018;
wire n_9820;
wire n_8635;
wire n_7758;
wire n_8320;
wire n_12477;
wire n_9703;
wire n_4472;
wire n_12516;
wire n_9819;
wire n_15422;
wire n_9118;
wire n_11060;
wire n_15722;
wire n_9321;
wire n_12523;
wire n_11493;
wire n_11562;
wire n_13698;
wire n_5819;
wire n_5180;
wire n_10703;
wire n_8375;
wire n_11575;
wire n_13462;
wire n_10449;
wire n_14959;
wire n_16114;
wire n_14806;
wire n_10280;
wire n_9428;
wire n_8612;
wire n_10198;
wire n_8778;
wire n_11065;
wire n_5893;
wire n_9292;
wire n_11452;
wire n_15366;
wire n_7705;
wire n_6092;
wire n_12486;
wire n_6462;
wire n_15977;
wire n_11345;
wire n_4519;
wire n_15989;
wire n_9018;
wire n_13741;
wire n_5025;
wire n_8872;
wire n_12743;
wire n_10371;
wire n_7333;
wire n_12246;
wire n_12297;
wire n_4197;
wire n_13440;
wire n_6669;
wire n_8006;
wire n_11495;
wire n_9565;
wire n_13325;
wire n_6251;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_13089;
wire n_13578;
wire n_7337;
wire n_5726;
wire n_4310;
wire n_4566;
wire n_7439;
wire n_4371;
wire n_12610;
wire n_14006;
wire n_14901;
wire n_14757;
wire n_10483;
wire n_12771;
wire n_5828;
wire n_7744;
wire n_7210;
wire n_10346;
wire n_11864;
wire n_6228;
wire n_15619;
wire n_16030;
wire n_10805;
wire n_14107;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_10059;
wire n_9961;
wire n_15990;
wire n_4749;
wire n_12763;
wire n_16038;
wire n_7707;
wire n_5924;
wire n_7733;
wire n_13496;
wire n_14536;
wire n_5545;
wire n_16174;
wire n_8458;
wire n_9603;
wire n_8853;
wire n_11293;
wire n_14950;
wire n_5083;
wire n_15122;
wire n_15341;
wire n_15159;
wire n_7684;
wire n_14834;
wire n_10700;
wire n_11984;
wire n_11961;
wire n_8306;
wire n_11981;
wire n_14599;
wire n_6997;
wire n_9692;
wire n_4238;
wire n_6371;
wire n_13222;
wire n_11559;
wire n_7673;
wire n_15391;
wire n_14642;
wire n_15674;
wire n_12172;
wire n_11942;
wire n_11207;
wire n_11686;
wire n_14809;
wire n_12280;
wire n_12883;
wire n_7187;
wire n_8013;
wire n_14897;
wire n_14476;
wire n_8342;
wire n_10502;
wire n_12064;
wire n_12480;
wire n_10974;
wire n_7313;
wire n_16212;
wire n_5899;
wire n_11239;
wire n_14221;
wire n_10511;
wire n_10250;
wire n_9012;
wire n_11482;
wire n_12682;
wire n_10831;
wire n_5122;
wire n_11992;
wire n_4189;
wire n_12621;
wire n_15843;
wire n_4479;
wire n_13754;
wire n_10613;
wire n_16254;
wire n_6641;
wire n_12283;
wire n_6463;
wire n_10351;
wire n_10172;
wire n_13285;
wire n_4986;
wire n_10333;
wire n_4668;
wire n_9868;
wire n_6264;
wire n_15789;
wire n_5782;
wire n_8119;
wire n_9264;
wire n_4168;
wire n_8582;
wire n_7036;
wire n_11479;
wire n_4298;
wire n_10594;
wire n_11814;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_13181;
wire n_11622;
wire n_8445;
wire n_12225;
wire n_9720;
wire n_4250;
wire n_15245;
wire n_13004;
wire n_11067;
wire n_8044;
wire n_13413;
wire n_5864;
wire n_8464;
wire n_8363;
wire n_8921;
wire n_12208;
wire n_14072;
wire n_13608;
wire n_15858;
wire n_12126;
wire n_13397;
wire n_15003;
wire n_11083;
wire n_14282;
wire n_10010;
wire n_10588;
wire n_11907;
wire n_12396;
wire n_12984;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_11952;
wire n_9646;
wire n_16109;
wire n_7480;
wire n_13997;
wire n_12158;
wire n_8843;
wire n_13513;
wire n_5185;
wire n_8405;
wire n_13232;
wire n_13296;
wire n_13816;
wire n_14713;
wire n_8376;
wire n_13859;
wire n_5032;
wire n_11506;
wire n_6990;
wire n_7071;
wire n_5034;
wire n_10797;
wire n_8694;
wire n_8848;
wire n_6288;
wire n_13989;
wire n_14573;
wire n_10643;
wire n_8752;
wire n_8894;
wire n_8625;
wire n_7380;
wire n_14058;
wire n_16118;
wire n_8813;
wire n_7708;
wire n_12690;
wire n_12813;
wire n_11524;
wire n_10905;
wire n_9842;
wire n_11859;
wire n_4128;
wire n_11228;
wire n_12725;
wire n_9671;
wire n_5269;
wire n_15025;
wire n_8430;
wire n_5709;
wire n_11035;
wire n_10784;
wire n_4807;
wire n_11023;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_14009;
wire n_5115;
wire n_12474;
wire n_7376;
wire n_11174;
wire n_8411;
wire n_13759;
wire n_8817;
wire n_8461;
wire n_10438;
wire n_15056;
wire n_14911;
wire n_10234;
wire n_10946;
wire n_11582;
wire n_9230;
wire n_5324;
wire n_4915;
wire n_4383;
wire n_4830;
wire n_11705;
wire n_4391;
wire n_11796;
wire n_12484;
wire n_9893;
wire n_6409;
wire n_8391;
wire n_8507;
wire n_12021;
wire n_5927;
wire n_8691;
wire n_9188;
wire n_11003;
wire n_4485;
wire n_9032;
wire n_7657;
wire n_6388;
wire n_10275;
wire n_15279;
wire n_6839;
wire n_14284;
wire n_5163;
wire n_9614;
wire n_8967;
wire n_12990;
wire n_4356;
wire n_9628;
wire n_9231;
wire n_10854;
wire n_6864;
wire n_14309;
wire n_13652;
wire n_13207;
wire n_4890;
wire n_10204;
wire n_8084;
wire n_8856;
wire n_15963;
wire n_12685;
wire n_12778;
wire n_6679;
wire n_12862;
wire n_11528;
wire n_10734;
wire n_13442;
wire n_10201;
wire n_8631;
wire n_16144;
wire n_6051;
wire n_15128;
wire n_4224;
wire n_8219;
wire n_16008;
wire n_9730;
wire n_5507;
wire n_15898;
wire n_10608;
wire n_4573;
wire n_10746;
wire n_4943;
wire n_10676;
wire n_6599;
wire n_14423;
wire n_12177;
wire n_13128;
wire n_7504;
wire n_14086;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_5642;
wire n_12672;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_8428;
wire n_9172;
wire n_12141;
wire n_14665;
wire n_14342;
wire n_9926;
wire n_14634;
wire n_6738;
wire n_12665;
wire n_13719;
wire n_5226;
wire n_11615;
wire n_11079;
wire n_8338;
wire n_14772;
wire n_7602;
wire n_9180;
wire n_9017;
wire n_12024;
wire n_12795;
wire n_9269;
wire n_6566;
wire n_9026;
wire n_13453;
wire n_9462;
wire n_10900;
wire n_5696;
wire n_7998;
wire n_13370;
wire n_8666;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_11438;
wire n_11700;
wire n_7557;
wire n_12940;
wire n_7408;
wire n_12555;
wire n_16123;
wire n_14539;
wire n_7026;
wire n_4335;
wire n_10052;
wire n_16215;
wire n_13656;
wire n_11668;
wire n_15286;
wire n_6146;
wire n_13667;
wire n_5677;
wire n_13641;
wire n_4277;
wire n_12487;
wire n_4614;
wire n_4629;
wire n_7394;
wire n_11387;
wire n_9515;
wire n_10560;
wire n_9502;
wire n_13103;
wire n_4516;
wire n_5235;
wire n_13183;
wire n_13720;
wire n_13971;
wire n_15650;
wire n_11099;
wire n_7627;
wire n_15929;
wire n_6436;
wire n_12305;
wire n_7719;
wire n_10773;
wire n_7450;
wire n_9316;
wire n_11996;
wire n_15962;
wire n_8938;
wire n_6081;
wire n_13436;
wire n_14479;
wire n_16098;
wire n_10455;
wire n_14410;
wire n_16148;
wire n_7852;
wire n_5724;
wire n_12526;
wire n_12622;
wire n_7462;
wire n_12456;
wire n_7780;
wire n_8523;
wire n_10391;
wire n_12857;
wire n_5979;
wire n_10476;
wire n_10559;
wire n_10630;
wire n_13797;
wire n_6027;
wire n_13321;
wire n_10911;
wire n_11547;
wire n_10121;
wire n_11064;
wire n_12439;
wire n_4467;
wire n_15785;
wire n_13809;
wire n_7582;
wire n_15522;
wire n_10540;
wire n_5521;
wire n_15140;
wire n_7421;
wire n_13575;
wire n_16239;
wire n_11104;
wire n_9873;
wire n_10473;
wire n_15120;
wire n_15234;
wire n_12287;
wire n_10828;
wire n_12182;
wire n_13390;
wire n_8924;
wire n_12366;
wire n_4955;
wire n_7555;
wire n_11112;
wire n_14915;
wire n_10114;
wire n_5410;
wire n_12552;
wire n_6110;
wire n_14123;
wire n_10269;
wire n_14258;
wire n_6238;
wire n_7025;
wire n_8380;
wire n_13371;
wire n_12777;
wire n_9978;
wire n_5241;
wire n_12492;
wire n_10418;
wire n_4248;
wire n_4645;
wire n_15235;
wire n_13231;
wire n_5331;
wire n_7478;
wire n_6326;
wire n_10672;
wire n_7451;
wire n_9494;
wire n_15918;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_14601;
wire n_11850;
wire n_12437;
wire n_6612;
wire n_10922;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g4123 ( 
.A(n_3925),
.Y(n_4123)
);

CKINVDCx5p33_ASAP7_75t_R g4124 ( 
.A(n_3360),
.Y(n_4124)
);

CKINVDCx5p33_ASAP7_75t_R g4125 ( 
.A(n_1965),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_872),
.Y(n_4126)
);

BUFx2_ASAP7_75t_L g4127 ( 
.A(n_3954),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_2146),
.Y(n_4128)
);

CKINVDCx20_ASAP7_75t_R g4129 ( 
.A(n_1933),
.Y(n_4129)
);

CKINVDCx5p33_ASAP7_75t_R g4130 ( 
.A(n_483),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_106),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3961),
.Y(n_4132)
);

CKINVDCx5p33_ASAP7_75t_R g4133 ( 
.A(n_861),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_1523),
.Y(n_4134)
);

CKINVDCx5p33_ASAP7_75t_R g4135 ( 
.A(n_904),
.Y(n_4135)
);

INVx2_ASAP7_75t_SL g4136 ( 
.A(n_4065),
.Y(n_4136)
);

CKINVDCx5p33_ASAP7_75t_R g4137 ( 
.A(n_358),
.Y(n_4137)
);

CKINVDCx5p33_ASAP7_75t_R g4138 ( 
.A(n_1845),
.Y(n_4138)
);

CKINVDCx5p33_ASAP7_75t_R g4139 ( 
.A(n_3390),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_575),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_2532),
.Y(n_4141)
);

CKINVDCx5p33_ASAP7_75t_R g4142 ( 
.A(n_2077),
.Y(n_4142)
);

CKINVDCx5p33_ASAP7_75t_R g4143 ( 
.A(n_3252),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_227),
.Y(n_4144)
);

CKINVDCx5p33_ASAP7_75t_R g4145 ( 
.A(n_1077),
.Y(n_4145)
);

CKINVDCx5p33_ASAP7_75t_R g4146 ( 
.A(n_3520),
.Y(n_4146)
);

CKINVDCx5p33_ASAP7_75t_R g4147 ( 
.A(n_2192),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_2630),
.Y(n_4148)
);

CKINVDCx5p33_ASAP7_75t_R g4149 ( 
.A(n_4039),
.Y(n_4149)
);

CKINVDCx5p33_ASAP7_75t_R g4150 ( 
.A(n_3834),
.Y(n_4150)
);

CKINVDCx5p33_ASAP7_75t_R g4151 ( 
.A(n_326),
.Y(n_4151)
);

BUFx8_ASAP7_75t_SL g4152 ( 
.A(n_289),
.Y(n_4152)
);

CKINVDCx5p33_ASAP7_75t_R g4153 ( 
.A(n_3212),
.Y(n_4153)
);

CKINVDCx5p33_ASAP7_75t_R g4154 ( 
.A(n_208),
.Y(n_4154)
);

CKINVDCx5p33_ASAP7_75t_R g4155 ( 
.A(n_4072),
.Y(n_4155)
);

CKINVDCx5p33_ASAP7_75t_R g4156 ( 
.A(n_3256),
.Y(n_4156)
);

CKINVDCx5p33_ASAP7_75t_R g4157 ( 
.A(n_3608),
.Y(n_4157)
);

BUFx3_ASAP7_75t_L g4158 ( 
.A(n_3097),
.Y(n_4158)
);

CKINVDCx5p33_ASAP7_75t_R g4159 ( 
.A(n_4060),
.Y(n_4159)
);

CKINVDCx5p33_ASAP7_75t_R g4160 ( 
.A(n_3988),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_1531),
.Y(n_4161)
);

CKINVDCx5p33_ASAP7_75t_R g4162 ( 
.A(n_89),
.Y(n_4162)
);

CKINVDCx5p33_ASAP7_75t_R g4163 ( 
.A(n_1434),
.Y(n_4163)
);

BUFx3_ASAP7_75t_L g4164 ( 
.A(n_1740),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_1958),
.Y(n_4165)
);

BUFx3_ASAP7_75t_L g4166 ( 
.A(n_1895),
.Y(n_4166)
);

CKINVDCx5p33_ASAP7_75t_R g4167 ( 
.A(n_2117),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_623),
.Y(n_4168)
);

CKINVDCx5p33_ASAP7_75t_R g4169 ( 
.A(n_3936),
.Y(n_4169)
);

CKINVDCx5p33_ASAP7_75t_R g4170 ( 
.A(n_636),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_736),
.Y(n_4171)
);

INVx2_ASAP7_75t_SL g4172 ( 
.A(n_4002),
.Y(n_4172)
);

CKINVDCx20_ASAP7_75t_R g4173 ( 
.A(n_166),
.Y(n_4173)
);

CKINVDCx5p33_ASAP7_75t_R g4174 ( 
.A(n_1194),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_1251),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_1286),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_1528),
.Y(n_4177)
);

INVx1_ASAP7_75t_SL g4178 ( 
.A(n_1699),
.Y(n_4178)
);

CKINVDCx5p33_ASAP7_75t_R g4179 ( 
.A(n_2802),
.Y(n_4179)
);

CKINVDCx5p33_ASAP7_75t_R g4180 ( 
.A(n_1135),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_548),
.Y(n_4181)
);

CKINVDCx5p33_ASAP7_75t_R g4182 ( 
.A(n_733),
.Y(n_4182)
);

BUFx2_ASAP7_75t_L g4183 ( 
.A(n_1091),
.Y(n_4183)
);

CKINVDCx5p33_ASAP7_75t_R g4184 ( 
.A(n_3913),
.Y(n_4184)
);

CKINVDCx5p33_ASAP7_75t_R g4185 ( 
.A(n_687),
.Y(n_4185)
);

CKINVDCx16_ASAP7_75t_R g4186 ( 
.A(n_819),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3433),
.Y(n_4187)
);

CKINVDCx5p33_ASAP7_75t_R g4188 ( 
.A(n_2180),
.Y(n_4188)
);

CKINVDCx5p33_ASAP7_75t_R g4189 ( 
.A(n_3898),
.Y(n_4189)
);

CKINVDCx5p33_ASAP7_75t_R g4190 ( 
.A(n_3387),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_169),
.Y(n_4191)
);

CKINVDCx5p33_ASAP7_75t_R g4192 ( 
.A(n_1661),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_422),
.Y(n_4193)
);

BUFx5_ASAP7_75t_L g4194 ( 
.A(n_708),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_2569),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_3070),
.Y(n_4196)
);

CKINVDCx5p33_ASAP7_75t_R g4197 ( 
.A(n_4037),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4064),
.Y(n_4198)
);

CKINVDCx5p33_ASAP7_75t_R g4199 ( 
.A(n_2898),
.Y(n_4199)
);

CKINVDCx5p33_ASAP7_75t_R g4200 ( 
.A(n_1119),
.Y(n_4200)
);

INVx1_ASAP7_75t_SL g4201 ( 
.A(n_2091),
.Y(n_4201)
);

CKINVDCx5p33_ASAP7_75t_R g4202 ( 
.A(n_3108),
.Y(n_4202)
);

INVx2_ASAP7_75t_SL g4203 ( 
.A(n_2580),
.Y(n_4203)
);

CKINVDCx16_ASAP7_75t_R g4204 ( 
.A(n_3930),
.Y(n_4204)
);

BUFx10_ASAP7_75t_L g4205 ( 
.A(n_3524),
.Y(n_4205)
);

CKINVDCx16_ASAP7_75t_R g4206 ( 
.A(n_1686),
.Y(n_4206)
);

CKINVDCx5p33_ASAP7_75t_R g4207 ( 
.A(n_2237),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_2199),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_686),
.Y(n_4209)
);

CKINVDCx5p33_ASAP7_75t_R g4210 ( 
.A(n_1679),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3302),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_893),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_1303),
.Y(n_4213)
);

BUFx5_ASAP7_75t_L g4214 ( 
.A(n_3683),
.Y(n_4214)
);

CKINVDCx5p33_ASAP7_75t_R g4215 ( 
.A(n_2832),
.Y(n_4215)
);

CKINVDCx5p33_ASAP7_75t_R g4216 ( 
.A(n_3042),
.Y(n_4216)
);

CKINVDCx5p33_ASAP7_75t_R g4217 ( 
.A(n_3080),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_2247),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_1525),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3983),
.Y(n_4220)
);

CKINVDCx20_ASAP7_75t_R g4221 ( 
.A(n_325),
.Y(n_4221)
);

CKINVDCx5p33_ASAP7_75t_R g4222 ( 
.A(n_2729),
.Y(n_4222)
);

CKINVDCx5p33_ASAP7_75t_R g4223 ( 
.A(n_4010),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_2564),
.Y(n_4224)
);

CKINVDCx5p33_ASAP7_75t_R g4225 ( 
.A(n_2259),
.Y(n_4225)
);

CKINVDCx5p33_ASAP7_75t_R g4226 ( 
.A(n_4014),
.Y(n_4226)
);

CKINVDCx16_ASAP7_75t_R g4227 ( 
.A(n_4083),
.Y(n_4227)
);

CKINVDCx5p33_ASAP7_75t_R g4228 ( 
.A(n_3212),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3907),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_1938),
.Y(n_4230)
);

CKINVDCx5p33_ASAP7_75t_R g4231 ( 
.A(n_2641),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_2524),
.Y(n_4232)
);

CKINVDCx14_ASAP7_75t_R g4233 ( 
.A(n_3927),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_326),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_1980),
.Y(n_4235)
);

CKINVDCx5p33_ASAP7_75t_R g4236 ( 
.A(n_4043),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_2363),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_381),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_1375),
.Y(n_4239)
);

CKINVDCx5p33_ASAP7_75t_R g4240 ( 
.A(n_834),
.Y(n_4240)
);

BUFx10_ASAP7_75t_L g4241 ( 
.A(n_172),
.Y(n_4241)
);

CKINVDCx20_ASAP7_75t_R g4242 ( 
.A(n_1709),
.Y(n_4242)
);

BUFx3_ASAP7_75t_L g4243 ( 
.A(n_2674),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_947),
.Y(n_4244)
);

CKINVDCx5p33_ASAP7_75t_R g4245 ( 
.A(n_62),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_2633),
.Y(n_4246)
);

CKINVDCx16_ASAP7_75t_R g4247 ( 
.A(n_1793),
.Y(n_4247)
);

CKINVDCx5p33_ASAP7_75t_R g4248 ( 
.A(n_2553),
.Y(n_4248)
);

CKINVDCx5p33_ASAP7_75t_R g4249 ( 
.A(n_670),
.Y(n_4249)
);

CKINVDCx5p33_ASAP7_75t_R g4250 ( 
.A(n_4094),
.Y(n_4250)
);

CKINVDCx5p33_ASAP7_75t_R g4251 ( 
.A(n_3369),
.Y(n_4251)
);

CKINVDCx5p33_ASAP7_75t_R g4252 ( 
.A(n_1306),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_1675),
.Y(n_4253)
);

CKINVDCx5p33_ASAP7_75t_R g4254 ( 
.A(n_3917),
.Y(n_4254)
);

CKINVDCx5p33_ASAP7_75t_R g4255 ( 
.A(n_3228),
.Y(n_4255)
);

CKINVDCx5p33_ASAP7_75t_R g4256 ( 
.A(n_237),
.Y(n_4256)
);

CKINVDCx5p33_ASAP7_75t_R g4257 ( 
.A(n_3031),
.Y(n_4257)
);

CKINVDCx5p33_ASAP7_75t_R g4258 ( 
.A(n_3724),
.Y(n_4258)
);

CKINVDCx5p33_ASAP7_75t_R g4259 ( 
.A(n_795),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3162),
.Y(n_4260)
);

CKINVDCx5p33_ASAP7_75t_R g4261 ( 
.A(n_3650),
.Y(n_4261)
);

CKINVDCx5p33_ASAP7_75t_R g4262 ( 
.A(n_476),
.Y(n_4262)
);

CKINVDCx5p33_ASAP7_75t_R g4263 ( 
.A(n_2364),
.Y(n_4263)
);

CKINVDCx5p33_ASAP7_75t_R g4264 ( 
.A(n_945),
.Y(n_4264)
);

CKINVDCx5p33_ASAP7_75t_R g4265 ( 
.A(n_1678),
.Y(n_4265)
);

CKINVDCx20_ASAP7_75t_R g4266 ( 
.A(n_3844),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3459),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_3092),
.Y(n_4268)
);

CKINVDCx5p33_ASAP7_75t_R g4269 ( 
.A(n_345),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_647),
.Y(n_4270)
);

INVx2_ASAP7_75t_SL g4271 ( 
.A(n_3912),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_2194),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_2421),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_2827),
.Y(n_4274)
);

CKINVDCx5p33_ASAP7_75t_R g4275 ( 
.A(n_1891),
.Y(n_4275)
);

INVxp67_ASAP7_75t_L g4276 ( 
.A(n_3985),
.Y(n_4276)
);

BUFx6f_ASAP7_75t_L g4277 ( 
.A(n_4046),
.Y(n_4277)
);

CKINVDCx5p33_ASAP7_75t_R g4278 ( 
.A(n_2197),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_3645),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_2808),
.Y(n_4280)
);

CKINVDCx5p33_ASAP7_75t_R g4281 ( 
.A(n_1847),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_1088),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3977),
.Y(n_4283)
);

CKINVDCx5p33_ASAP7_75t_R g4284 ( 
.A(n_3420),
.Y(n_4284)
);

CKINVDCx5p33_ASAP7_75t_R g4285 ( 
.A(n_2844),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_537),
.Y(n_4286)
);

INVx1_ASAP7_75t_SL g4287 ( 
.A(n_569),
.Y(n_4287)
);

CKINVDCx5p33_ASAP7_75t_R g4288 ( 
.A(n_3627),
.Y(n_4288)
);

CKINVDCx5p33_ASAP7_75t_R g4289 ( 
.A(n_461),
.Y(n_4289)
);

CKINVDCx20_ASAP7_75t_R g4290 ( 
.A(n_178),
.Y(n_4290)
);

CKINVDCx5p33_ASAP7_75t_R g4291 ( 
.A(n_502),
.Y(n_4291)
);

CKINVDCx20_ASAP7_75t_R g4292 ( 
.A(n_3795),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_1044),
.Y(n_4293)
);

CKINVDCx5p33_ASAP7_75t_R g4294 ( 
.A(n_2436),
.Y(n_4294)
);

CKINVDCx5p33_ASAP7_75t_R g4295 ( 
.A(n_3757),
.Y(n_4295)
);

CKINVDCx5p33_ASAP7_75t_R g4296 ( 
.A(n_2588),
.Y(n_4296)
);

BUFx3_ASAP7_75t_L g4297 ( 
.A(n_772),
.Y(n_4297)
);

CKINVDCx5p33_ASAP7_75t_R g4298 ( 
.A(n_4090),
.Y(n_4298)
);

INVx2_ASAP7_75t_SL g4299 ( 
.A(n_3923),
.Y(n_4299)
);

CKINVDCx5p33_ASAP7_75t_R g4300 ( 
.A(n_3793),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_112),
.Y(n_4301)
);

CKINVDCx5p33_ASAP7_75t_R g4302 ( 
.A(n_2684),
.Y(n_4302)
);

CKINVDCx5p33_ASAP7_75t_R g4303 ( 
.A(n_1204),
.Y(n_4303)
);

BUFx2_ASAP7_75t_L g4304 ( 
.A(n_3616),
.Y(n_4304)
);

CKINVDCx5p33_ASAP7_75t_R g4305 ( 
.A(n_618),
.Y(n_4305)
);

CKINVDCx5p33_ASAP7_75t_R g4306 ( 
.A(n_539),
.Y(n_4306)
);

CKINVDCx5p33_ASAP7_75t_R g4307 ( 
.A(n_2665),
.Y(n_4307)
);

CKINVDCx5p33_ASAP7_75t_R g4308 ( 
.A(n_2918),
.Y(n_4308)
);

BUFx10_ASAP7_75t_L g4309 ( 
.A(n_1946),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_192),
.Y(n_4310)
);

CKINVDCx5p33_ASAP7_75t_R g4311 ( 
.A(n_3070),
.Y(n_4311)
);

CKINVDCx16_ASAP7_75t_R g4312 ( 
.A(n_3969),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3732),
.Y(n_4313)
);

CKINVDCx20_ASAP7_75t_R g4314 ( 
.A(n_1111),
.Y(n_4314)
);

CKINVDCx5p33_ASAP7_75t_R g4315 ( 
.A(n_1749),
.Y(n_4315)
);

CKINVDCx5p33_ASAP7_75t_R g4316 ( 
.A(n_554),
.Y(n_4316)
);

BUFx3_ASAP7_75t_L g4317 ( 
.A(n_3967),
.Y(n_4317)
);

CKINVDCx5p33_ASAP7_75t_R g4318 ( 
.A(n_3057),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_1701),
.Y(n_4319)
);

CKINVDCx5p33_ASAP7_75t_R g4320 ( 
.A(n_196),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_537),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_735),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3928),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_3131),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_559),
.Y(n_4325)
);

BUFx3_ASAP7_75t_L g4326 ( 
.A(n_3073),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_721),
.Y(n_4327)
);

CKINVDCx20_ASAP7_75t_R g4328 ( 
.A(n_2805),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_1164),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_2840),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_2383),
.Y(n_4331)
);

BUFx3_ASAP7_75t_L g4332 ( 
.A(n_310),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_515),
.Y(n_4333)
);

CKINVDCx5p33_ASAP7_75t_R g4334 ( 
.A(n_206),
.Y(n_4334)
);

CKINVDCx20_ASAP7_75t_R g4335 ( 
.A(n_4056),
.Y(n_4335)
);

CKINVDCx20_ASAP7_75t_R g4336 ( 
.A(n_727),
.Y(n_4336)
);

CKINVDCx5p33_ASAP7_75t_R g4337 ( 
.A(n_1490),
.Y(n_4337)
);

CKINVDCx20_ASAP7_75t_R g4338 ( 
.A(n_1506),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_3362),
.Y(n_4339)
);

CKINVDCx5p33_ASAP7_75t_R g4340 ( 
.A(n_2158),
.Y(n_4340)
);

CKINVDCx20_ASAP7_75t_R g4341 ( 
.A(n_878),
.Y(n_4341)
);

CKINVDCx5p33_ASAP7_75t_R g4342 ( 
.A(n_909),
.Y(n_4342)
);

CKINVDCx5p33_ASAP7_75t_R g4343 ( 
.A(n_108),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3842),
.Y(n_4344)
);

CKINVDCx5p33_ASAP7_75t_R g4345 ( 
.A(n_3362),
.Y(n_4345)
);

CKINVDCx5p33_ASAP7_75t_R g4346 ( 
.A(n_1199),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_3800),
.Y(n_4347)
);

CKINVDCx5p33_ASAP7_75t_R g4348 ( 
.A(n_2298),
.Y(n_4348)
);

CKINVDCx5p33_ASAP7_75t_R g4349 ( 
.A(n_10),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_1938),
.Y(n_4350)
);

CKINVDCx5p33_ASAP7_75t_R g4351 ( 
.A(n_2361),
.Y(n_4351)
);

INVx1_ASAP7_75t_SL g4352 ( 
.A(n_141),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_3468),
.Y(n_4353)
);

CKINVDCx5p33_ASAP7_75t_R g4354 ( 
.A(n_663),
.Y(n_4354)
);

CKINVDCx5p33_ASAP7_75t_R g4355 ( 
.A(n_2695),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_2391),
.Y(n_4356)
);

CKINVDCx5p33_ASAP7_75t_R g4357 ( 
.A(n_3996),
.Y(n_4357)
);

CKINVDCx5p33_ASAP7_75t_R g4358 ( 
.A(n_2216),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_1375),
.Y(n_4359)
);

BUFx2_ASAP7_75t_L g4360 ( 
.A(n_1424),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_2345),
.Y(n_4361)
);

CKINVDCx5p33_ASAP7_75t_R g4362 ( 
.A(n_1522),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_1922),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_93),
.Y(n_4364)
);

CKINVDCx5p33_ASAP7_75t_R g4365 ( 
.A(n_1406),
.Y(n_4365)
);

BUFx8_ASAP7_75t_SL g4366 ( 
.A(n_2904),
.Y(n_4366)
);

CKINVDCx20_ASAP7_75t_R g4367 ( 
.A(n_1457),
.Y(n_4367)
);

CKINVDCx5p33_ASAP7_75t_R g4368 ( 
.A(n_621),
.Y(n_4368)
);

BUFx2_ASAP7_75t_L g4369 ( 
.A(n_501),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_2217),
.Y(n_4370)
);

CKINVDCx5p33_ASAP7_75t_R g4371 ( 
.A(n_3261),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_494),
.Y(n_4372)
);

CKINVDCx5p33_ASAP7_75t_R g4373 ( 
.A(n_2265),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_2626),
.Y(n_4374)
);

CKINVDCx5p33_ASAP7_75t_R g4375 ( 
.A(n_3897),
.Y(n_4375)
);

CKINVDCx5p33_ASAP7_75t_R g4376 ( 
.A(n_39),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_2186),
.Y(n_4377)
);

CKINVDCx5p33_ASAP7_75t_R g4378 ( 
.A(n_3456),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_1165),
.Y(n_4379)
);

CKINVDCx5p33_ASAP7_75t_R g4380 ( 
.A(n_3790),
.Y(n_4380)
);

CKINVDCx5p33_ASAP7_75t_R g4381 ( 
.A(n_3864),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_1307),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_1762),
.Y(n_4383)
);

CKINVDCx5p33_ASAP7_75t_R g4384 ( 
.A(n_3932),
.Y(n_4384)
);

CKINVDCx5p33_ASAP7_75t_R g4385 ( 
.A(n_3726),
.Y(n_4385)
);

CKINVDCx5p33_ASAP7_75t_R g4386 ( 
.A(n_3945),
.Y(n_4386)
);

CKINVDCx5p33_ASAP7_75t_R g4387 ( 
.A(n_3286),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_1907),
.Y(n_4388)
);

CKINVDCx20_ASAP7_75t_R g4389 ( 
.A(n_4036),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_3980),
.Y(n_4390)
);

INVx1_ASAP7_75t_SL g4391 ( 
.A(n_3943),
.Y(n_4391)
);

INVx2_ASAP7_75t_SL g4392 ( 
.A(n_3710),
.Y(n_4392)
);

CKINVDCx5p33_ASAP7_75t_R g4393 ( 
.A(n_2837),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_1851),
.Y(n_4394)
);

CKINVDCx5p33_ASAP7_75t_R g4395 ( 
.A(n_3051),
.Y(n_4395)
);

CKINVDCx5p33_ASAP7_75t_R g4396 ( 
.A(n_529),
.Y(n_4396)
);

CKINVDCx5p33_ASAP7_75t_R g4397 ( 
.A(n_4068),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_1877),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_2044),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_551),
.Y(n_4400)
);

CKINVDCx5p33_ASAP7_75t_R g4401 ( 
.A(n_296),
.Y(n_4401)
);

CKINVDCx5p33_ASAP7_75t_R g4402 ( 
.A(n_1969),
.Y(n_4402)
);

CKINVDCx5p33_ASAP7_75t_R g4403 ( 
.A(n_3028),
.Y(n_4403)
);

CKINVDCx5p33_ASAP7_75t_R g4404 ( 
.A(n_2250),
.Y(n_4404)
);

CKINVDCx5p33_ASAP7_75t_R g4405 ( 
.A(n_3444),
.Y(n_4405)
);

CKINVDCx16_ASAP7_75t_R g4406 ( 
.A(n_65),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_627),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_815),
.Y(n_4408)
);

CKINVDCx5p33_ASAP7_75t_R g4409 ( 
.A(n_2263),
.Y(n_4409)
);

BUFx2_ASAP7_75t_SL g4410 ( 
.A(n_2984),
.Y(n_4410)
);

CKINVDCx5p33_ASAP7_75t_R g4411 ( 
.A(n_4031),
.Y(n_4411)
);

CKINVDCx5p33_ASAP7_75t_R g4412 ( 
.A(n_2800),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_349),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_2085),
.Y(n_4414)
);

CKINVDCx5p33_ASAP7_75t_R g4415 ( 
.A(n_1311),
.Y(n_4415)
);

CKINVDCx5p33_ASAP7_75t_R g4416 ( 
.A(n_1721),
.Y(n_4416)
);

CKINVDCx5p33_ASAP7_75t_R g4417 ( 
.A(n_3950),
.Y(n_4417)
);

CKINVDCx20_ASAP7_75t_R g4418 ( 
.A(n_2134),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_2161),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_2565),
.Y(n_4420)
);

CKINVDCx5p33_ASAP7_75t_R g4421 ( 
.A(n_2051),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_3888),
.Y(n_4422)
);

INVx1_ASAP7_75t_SL g4423 ( 
.A(n_3443),
.Y(n_4423)
);

INVx2_ASAP7_75t_SL g4424 ( 
.A(n_2070),
.Y(n_4424)
);

CKINVDCx5p33_ASAP7_75t_R g4425 ( 
.A(n_2096),
.Y(n_4425)
);

CKINVDCx5p33_ASAP7_75t_R g4426 ( 
.A(n_3174),
.Y(n_4426)
);

CKINVDCx20_ASAP7_75t_R g4427 ( 
.A(n_4023),
.Y(n_4427)
);

CKINVDCx5p33_ASAP7_75t_R g4428 ( 
.A(n_249),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_2230),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_1934),
.Y(n_4430)
);

CKINVDCx5p33_ASAP7_75t_R g4431 ( 
.A(n_1020),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_3850),
.Y(n_4432)
);

CKINVDCx20_ASAP7_75t_R g4433 ( 
.A(n_3251),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_2285),
.Y(n_4434)
);

CKINVDCx5p33_ASAP7_75t_R g4435 ( 
.A(n_1067),
.Y(n_4435)
);

CKINVDCx5p33_ASAP7_75t_R g4436 ( 
.A(n_3867),
.Y(n_4436)
);

CKINVDCx5p33_ASAP7_75t_R g4437 ( 
.A(n_2596),
.Y(n_4437)
);

CKINVDCx5p33_ASAP7_75t_R g4438 ( 
.A(n_789),
.Y(n_4438)
);

CKINVDCx5p33_ASAP7_75t_R g4439 ( 
.A(n_758),
.Y(n_4439)
);

CKINVDCx5p33_ASAP7_75t_R g4440 ( 
.A(n_3964),
.Y(n_4440)
);

CKINVDCx5p33_ASAP7_75t_R g4441 ( 
.A(n_2075),
.Y(n_4441)
);

CKINVDCx5p33_ASAP7_75t_R g4442 ( 
.A(n_3301),
.Y(n_4442)
);

BUFx5_ASAP7_75t_L g4443 ( 
.A(n_3972),
.Y(n_4443)
);

CKINVDCx5p33_ASAP7_75t_R g4444 ( 
.A(n_2774),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_3952),
.Y(n_4445)
);

CKINVDCx20_ASAP7_75t_R g4446 ( 
.A(n_3356),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_2778),
.Y(n_4447)
);

CKINVDCx5p33_ASAP7_75t_R g4448 ( 
.A(n_1573),
.Y(n_4448)
);

CKINVDCx20_ASAP7_75t_R g4449 ( 
.A(n_2469),
.Y(n_4449)
);

CKINVDCx20_ASAP7_75t_R g4450 ( 
.A(n_2309),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_3030),
.Y(n_4451)
);

CKINVDCx5p33_ASAP7_75t_R g4452 ( 
.A(n_3514),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_1129),
.Y(n_4453)
);

CKINVDCx20_ASAP7_75t_R g4454 ( 
.A(n_1699),
.Y(n_4454)
);

CKINVDCx5p33_ASAP7_75t_R g4455 ( 
.A(n_556),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_1808),
.Y(n_4456)
);

CKINVDCx5p33_ASAP7_75t_R g4457 ( 
.A(n_4069),
.Y(n_4457)
);

CKINVDCx5p33_ASAP7_75t_R g4458 ( 
.A(n_4035),
.Y(n_4458)
);

BUFx2_ASAP7_75t_L g4459 ( 
.A(n_1829),
.Y(n_4459)
);

CKINVDCx5p33_ASAP7_75t_R g4460 ( 
.A(n_1361),
.Y(n_4460)
);

CKINVDCx5p33_ASAP7_75t_R g4461 ( 
.A(n_3481),
.Y(n_4461)
);

CKINVDCx5p33_ASAP7_75t_R g4462 ( 
.A(n_1103),
.Y(n_4462)
);

CKINVDCx5p33_ASAP7_75t_R g4463 ( 
.A(n_1022),
.Y(n_4463)
);

CKINVDCx5p33_ASAP7_75t_R g4464 ( 
.A(n_2870),
.Y(n_4464)
);

BUFx2_ASAP7_75t_SL g4465 ( 
.A(n_1417),
.Y(n_4465)
);

CKINVDCx5p33_ASAP7_75t_R g4466 ( 
.A(n_3986),
.Y(n_4466)
);

CKINVDCx5p33_ASAP7_75t_R g4467 ( 
.A(n_1670),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_42),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_3412),
.Y(n_4469)
);

INVx1_ASAP7_75t_SL g4470 ( 
.A(n_2797),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_1261),
.Y(n_4471)
);

CKINVDCx5p33_ASAP7_75t_R g4472 ( 
.A(n_4053),
.Y(n_4472)
);

CKINVDCx5p33_ASAP7_75t_R g4473 ( 
.A(n_3966),
.Y(n_4473)
);

BUFx3_ASAP7_75t_L g4474 ( 
.A(n_3257),
.Y(n_4474)
);

CKINVDCx5p33_ASAP7_75t_R g4475 ( 
.A(n_3626),
.Y(n_4475)
);

CKINVDCx5p33_ASAP7_75t_R g4476 ( 
.A(n_2879),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_3176),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_2852),
.Y(n_4478)
);

CKINVDCx5p33_ASAP7_75t_R g4479 ( 
.A(n_2851),
.Y(n_4479)
);

CKINVDCx5p33_ASAP7_75t_R g4480 ( 
.A(n_1602),
.Y(n_4480)
);

CKINVDCx5p33_ASAP7_75t_R g4481 ( 
.A(n_4063),
.Y(n_4481)
);

CKINVDCx5p33_ASAP7_75t_R g4482 ( 
.A(n_1341),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3738),
.Y(n_4483)
);

CKINVDCx5p33_ASAP7_75t_R g4484 ( 
.A(n_3992),
.Y(n_4484)
);

BUFx3_ASAP7_75t_L g4485 ( 
.A(n_207),
.Y(n_4485)
);

CKINVDCx5p33_ASAP7_75t_R g4486 ( 
.A(n_685),
.Y(n_4486)
);

CKINVDCx20_ASAP7_75t_R g4487 ( 
.A(n_466),
.Y(n_4487)
);

CKINVDCx20_ASAP7_75t_R g4488 ( 
.A(n_4052),
.Y(n_4488)
);

CKINVDCx5p33_ASAP7_75t_R g4489 ( 
.A(n_3064),
.Y(n_4489)
);

CKINVDCx5p33_ASAP7_75t_R g4490 ( 
.A(n_443),
.Y(n_4490)
);

CKINVDCx5p33_ASAP7_75t_R g4491 ( 
.A(n_4109),
.Y(n_4491)
);

CKINVDCx5p33_ASAP7_75t_R g4492 ( 
.A(n_2294),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_3636),
.Y(n_4493)
);

CKINVDCx5p33_ASAP7_75t_R g4494 ( 
.A(n_2771),
.Y(n_4494)
);

INVx2_ASAP7_75t_SL g4495 ( 
.A(n_913),
.Y(n_4495)
);

BUFx3_ASAP7_75t_L g4496 ( 
.A(n_2002),
.Y(n_4496)
);

CKINVDCx5p33_ASAP7_75t_R g4497 ( 
.A(n_4098),
.Y(n_4497)
);

CKINVDCx5p33_ASAP7_75t_R g4498 ( 
.A(n_1104),
.Y(n_4498)
);

CKINVDCx5p33_ASAP7_75t_R g4499 ( 
.A(n_3990),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_4009),
.Y(n_4500)
);

CKINVDCx5p33_ASAP7_75t_R g4501 ( 
.A(n_4067),
.Y(n_4501)
);

CKINVDCx5p33_ASAP7_75t_R g4502 ( 
.A(n_2558),
.Y(n_4502)
);

CKINVDCx5p33_ASAP7_75t_R g4503 ( 
.A(n_3991),
.Y(n_4503)
);

CKINVDCx14_ASAP7_75t_R g4504 ( 
.A(n_1890),
.Y(n_4504)
);

CKINVDCx5p33_ASAP7_75t_R g4505 ( 
.A(n_703),
.Y(n_4505)
);

CKINVDCx5p33_ASAP7_75t_R g4506 ( 
.A(n_1261),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_2869),
.Y(n_4507)
);

CKINVDCx5p33_ASAP7_75t_R g4508 ( 
.A(n_858),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_2242),
.Y(n_4509)
);

BUFx2_ASAP7_75t_L g4510 ( 
.A(n_2323),
.Y(n_4510)
);

CKINVDCx5p33_ASAP7_75t_R g4511 ( 
.A(n_1420),
.Y(n_4511)
);

CKINVDCx5p33_ASAP7_75t_R g4512 ( 
.A(n_53),
.Y(n_4512)
);

CKINVDCx5p33_ASAP7_75t_R g4513 ( 
.A(n_2071),
.Y(n_4513)
);

HB1xp67_ASAP7_75t_L g4514 ( 
.A(n_3917),
.Y(n_4514)
);

CKINVDCx5p33_ASAP7_75t_R g4515 ( 
.A(n_1020),
.Y(n_4515)
);

CKINVDCx5p33_ASAP7_75t_R g4516 ( 
.A(n_3464),
.Y(n_4516)
);

INVx2_ASAP7_75t_SL g4517 ( 
.A(n_86),
.Y(n_4517)
);

CKINVDCx5p33_ASAP7_75t_R g4518 ( 
.A(n_4080),
.Y(n_4518)
);

CKINVDCx5p33_ASAP7_75t_R g4519 ( 
.A(n_4011),
.Y(n_4519)
);

CKINVDCx5p33_ASAP7_75t_R g4520 ( 
.A(n_2373),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_805),
.Y(n_4521)
);

CKINVDCx5p33_ASAP7_75t_R g4522 ( 
.A(n_2533),
.Y(n_4522)
);

CKINVDCx5p33_ASAP7_75t_R g4523 ( 
.A(n_1851),
.Y(n_4523)
);

CKINVDCx5p33_ASAP7_75t_R g4524 ( 
.A(n_753),
.Y(n_4524)
);

INVx2_ASAP7_75t_SL g4525 ( 
.A(n_1423),
.Y(n_4525)
);

CKINVDCx20_ASAP7_75t_R g4526 ( 
.A(n_3170),
.Y(n_4526)
);

CKINVDCx5p33_ASAP7_75t_R g4527 ( 
.A(n_2834),
.Y(n_4527)
);

CKINVDCx5p33_ASAP7_75t_R g4528 ( 
.A(n_2758),
.Y(n_4528)
);

CKINVDCx5p33_ASAP7_75t_R g4529 ( 
.A(n_3150),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_92),
.Y(n_4530)
);

CKINVDCx5p33_ASAP7_75t_R g4531 ( 
.A(n_1881),
.Y(n_4531)
);

CKINVDCx5p33_ASAP7_75t_R g4532 ( 
.A(n_1617),
.Y(n_4532)
);

CKINVDCx5p33_ASAP7_75t_R g4533 ( 
.A(n_3924),
.Y(n_4533)
);

CKINVDCx20_ASAP7_75t_R g4534 ( 
.A(n_527),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_510),
.Y(n_4535)
);

CKINVDCx5p33_ASAP7_75t_R g4536 ( 
.A(n_3757),
.Y(n_4536)
);

CKINVDCx5p33_ASAP7_75t_R g4537 ( 
.A(n_3718),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_4026),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_810),
.Y(n_4539)
);

INVx1_ASAP7_75t_SL g4540 ( 
.A(n_1937),
.Y(n_4540)
);

CKINVDCx5p33_ASAP7_75t_R g4541 ( 
.A(n_1566),
.Y(n_4541)
);

CKINVDCx5p33_ASAP7_75t_R g4542 ( 
.A(n_1642),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_520),
.Y(n_4543)
);

CKINVDCx5p33_ASAP7_75t_R g4544 ( 
.A(n_1914),
.Y(n_4544)
);

CKINVDCx5p33_ASAP7_75t_R g4545 ( 
.A(n_388),
.Y(n_4545)
);

CKINVDCx5p33_ASAP7_75t_R g4546 ( 
.A(n_4077),
.Y(n_4546)
);

CKINVDCx5p33_ASAP7_75t_R g4547 ( 
.A(n_3991),
.Y(n_4547)
);

BUFx2_ASAP7_75t_L g4548 ( 
.A(n_1683),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_3091),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_3361),
.Y(n_4550)
);

CKINVDCx5p33_ASAP7_75t_R g4551 ( 
.A(n_57),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4036),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_1704),
.Y(n_4553)
);

CKINVDCx5p33_ASAP7_75t_R g4554 ( 
.A(n_1107),
.Y(n_4554)
);

INVx1_ASAP7_75t_SL g4555 ( 
.A(n_1988),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_3971),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_3352),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_334),
.Y(n_4558)
);

CKINVDCx20_ASAP7_75t_R g4559 ( 
.A(n_3736),
.Y(n_4559)
);

CKINVDCx5p33_ASAP7_75t_R g4560 ( 
.A(n_1352),
.Y(n_4560)
);

CKINVDCx5p33_ASAP7_75t_R g4561 ( 
.A(n_743),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_3031),
.Y(n_4562)
);

CKINVDCx5p33_ASAP7_75t_R g4563 ( 
.A(n_1299),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_3939),
.Y(n_4564)
);

CKINVDCx5p33_ASAP7_75t_R g4565 ( 
.A(n_2304),
.Y(n_4565)
);

CKINVDCx5p33_ASAP7_75t_R g4566 ( 
.A(n_2455),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_3955),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_739),
.Y(n_4568)
);

BUFx5_ASAP7_75t_L g4569 ( 
.A(n_1916),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_2168),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_550),
.Y(n_4571)
);

CKINVDCx5p33_ASAP7_75t_R g4572 ( 
.A(n_2671),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_3014),
.Y(n_4573)
);

CKINVDCx5p33_ASAP7_75t_R g4574 ( 
.A(n_829),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4023),
.Y(n_4575)
);

CKINVDCx5p33_ASAP7_75t_R g4576 ( 
.A(n_1576),
.Y(n_4576)
);

BUFx8_ASAP7_75t_SL g4577 ( 
.A(n_164),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_1709),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_3935),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_1580),
.Y(n_4580)
);

CKINVDCx20_ASAP7_75t_R g4581 ( 
.A(n_4029),
.Y(n_4581)
);

CKINVDCx5p33_ASAP7_75t_R g4582 ( 
.A(n_3944),
.Y(n_4582)
);

CKINVDCx20_ASAP7_75t_R g4583 ( 
.A(n_1840),
.Y(n_4583)
);

CKINVDCx5p33_ASAP7_75t_R g4584 ( 
.A(n_2105),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_3457),
.Y(n_4585)
);

CKINVDCx5p33_ASAP7_75t_R g4586 ( 
.A(n_2974),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_25),
.Y(n_4587)
);

INVx2_ASAP7_75t_SL g4588 ( 
.A(n_2615),
.Y(n_4588)
);

CKINVDCx5p33_ASAP7_75t_R g4589 ( 
.A(n_1104),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_1137),
.Y(n_4590)
);

CKINVDCx5p33_ASAP7_75t_R g4591 ( 
.A(n_2),
.Y(n_4591)
);

CKINVDCx5p33_ASAP7_75t_R g4592 ( 
.A(n_764),
.Y(n_4592)
);

INVx1_ASAP7_75t_SL g4593 ( 
.A(n_3054),
.Y(n_4593)
);

CKINVDCx5p33_ASAP7_75t_R g4594 ( 
.A(n_1978),
.Y(n_4594)
);

CKINVDCx5p33_ASAP7_75t_R g4595 ( 
.A(n_3144),
.Y(n_4595)
);

CKINVDCx5p33_ASAP7_75t_R g4596 ( 
.A(n_3133),
.Y(n_4596)
);

CKINVDCx5p33_ASAP7_75t_R g4597 ( 
.A(n_4084),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_2390),
.Y(n_4598)
);

BUFx3_ASAP7_75t_L g4599 ( 
.A(n_1081),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_2364),
.Y(n_4600)
);

CKINVDCx20_ASAP7_75t_R g4601 ( 
.A(n_1461),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4007),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_2229),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_522),
.Y(n_4604)
);

CKINVDCx5p33_ASAP7_75t_R g4605 ( 
.A(n_4003),
.Y(n_4605)
);

CKINVDCx5p33_ASAP7_75t_R g4606 ( 
.A(n_1614),
.Y(n_4606)
);

CKINVDCx5p33_ASAP7_75t_R g4607 ( 
.A(n_604),
.Y(n_4607)
);

CKINVDCx5p33_ASAP7_75t_R g4608 ( 
.A(n_2251),
.Y(n_4608)
);

CKINVDCx5p33_ASAP7_75t_R g4609 ( 
.A(n_1915),
.Y(n_4609)
);

CKINVDCx5p33_ASAP7_75t_R g4610 ( 
.A(n_1069),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_3272),
.Y(n_4611)
);

INVx2_ASAP7_75t_SL g4612 ( 
.A(n_304),
.Y(n_4612)
);

INVxp67_ASAP7_75t_SL g4613 ( 
.A(n_1863),
.Y(n_4613)
);

INVx1_ASAP7_75t_SL g4614 ( 
.A(n_887),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_1600),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_2855),
.Y(n_4616)
);

INVx2_ASAP7_75t_SL g4617 ( 
.A(n_925),
.Y(n_4617)
);

CKINVDCx5p33_ASAP7_75t_R g4618 ( 
.A(n_3151),
.Y(n_4618)
);

CKINVDCx20_ASAP7_75t_R g4619 ( 
.A(n_1270),
.Y(n_4619)
);

CKINVDCx5p33_ASAP7_75t_R g4620 ( 
.A(n_1911),
.Y(n_4620)
);

CKINVDCx5p33_ASAP7_75t_R g4621 ( 
.A(n_1527),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_2313),
.Y(n_4622)
);

CKINVDCx5p33_ASAP7_75t_R g4623 ( 
.A(n_2434),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_3817),
.Y(n_4624)
);

BUFx3_ASAP7_75t_L g4625 ( 
.A(n_229),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_3100),
.Y(n_4626)
);

CKINVDCx5p33_ASAP7_75t_R g4627 ( 
.A(n_662),
.Y(n_4627)
);

CKINVDCx20_ASAP7_75t_R g4628 ( 
.A(n_3204),
.Y(n_4628)
);

BUFx6f_ASAP7_75t_L g4629 ( 
.A(n_1237),
.Y(n_4629)
);

CKINVDCx5p33_ASAP7_75t_R g4630 ( 
.A(n_1753),
.Y(n_4630)
);

CKINVDCx20_ASAP7_75t_R g4631 ( 
.A(n_3004),
.Y(n_4631)
);

CKINVDCx5p33_ASAP7_75t_R g4632 ( 
.A(n_3830),
.Y(n_4632)
);

CKINVDCx5p33_ASAP7_75t_R g4633 ( 
.A(n_3683),
.Y(n_4633)
);

INVxp67_ASAP7_75t_SL g4634 ( 
.A(n_3116),
.Y(n_4634)
);

CKINVDCx20_ASAP7_75t_R g4635 ( 
.A(n_4032),
.Y(n_4635)
);

CKINVDCx5p33_ASAP7_75t_R g4636 ( 
.A(n_1318),
.Y(n_4636)
);

INVx1_ASAP7_75t_SL g4637 ( 
.A(n_4000),
.Y(n_4637)
);

CKINVDCx20_ASAP7_75t_R g4638 ( 
.A(n_3317),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_10),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4011),
.Y(n_4640)
);

INVx1_ASAP7_75t_SL g4641 ( 
.A(n_2701),
.Y(n_4641)
);

CKINVDCx5p33_ASAP7_75t_R g4642 ( 
.A(n_931),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_60),
.Y(n_4643)
);

CKINVDCx5p33_ASAP7_75t_R g4644 ( 
.A(n_912),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_1563),
.Y(n_4645)
);

CKINVDCx5p33_ASAP7_75t_R g4646 ( 
.A(n_2425),
.Y(n_4646)
);

CKINVDCx5p33_ASAP7_75t_R g4647 ( 
.A(n_340),
.Y(n_4647)
);

CKINVDCx20_ASAP7_75t_R g4648 ( 
.A(n_937),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_4029),
.Y(n_4649)
);

CKINVDCx5p33_ASAP7_75t_R g4650 ( 
.A(n_3798),
.Y(n_4650)
);

CKINVDCx5p33_ASAP7_75t_R g4651 ( 
.A(n_2365),
.Y(n_4651)
);

CKINVDCx5p33_ASAP7_75t_R g4652 ( 
.A(n_2640),
.Y(n_4652)
);

CKINVDCx5p33_ASAP7_75t_R g4653 ( 
.A(n_3987),
.Y(n_4653)
);

CKINVDCx20_ASAP7_75t_R g4654 ( 
.A(n_2109),
.Y(n_4654)
);

BUFx6f_ASAP7_75t_L g4655 ( 
.A(n_3946),
.Y(n_4655)
);

CKINVDCx5p33_ASAP7_75t_R g4656 ( 
.A(n_2818),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_2534),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_1156),
.Y(n_4658)
);

CKINVDCx20_ASAP7_75t_R g4659 ( 
.A(n_3958),
.Y(n_4659)
);

CKINVDCx5p33_ASAP7_75t_R g4660 ( 
.A(n_2059),
.Y(n_4660)
);

CKINVDCx5p33_ASAP7_75t_R g4661 ( 
.A(n_1361),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_498),
.Y(n_4662)
);

INVx1_ASAP7_75t_SL g4663 ( 
.A(n_1403),
.Y(n_4663)
);

CKINVDCx5p33_ASAP7_75t_R g4664 ( 
.A(n_2856),
.Y(n_4664)
);

CKINVDCx5p33_ASAP7_75t_R g4665 ( 
.A(n_2630),
.Y(n_4665)
);

CKINVDCx5p33_ASAP7_75t_R g4666 ( 
.A(n_242),
.Y(n_4666)
);

CKINVDCx5p33_ASAP7_75t_R g4667 ( 
.A(n_49),
.Y(n_4667)
);

CKINVDCx20_ASAP7_75t_R g4668 ( 
.A(n_748),
.Y(n_4668)
);

BUFx10_ASAP7_75t_L g4669 ( 
.A(n_638),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_511),
.Y(n_4670)
);

CKINVDCx5p33_ASAP7_75t_R g4671 ( 
.A(n_3978),
.Y(n_4671)
);

CKINVDCx20_ASAP7_75t_R g4672 ( 
.A(n_2623),
.Y(n_4672)
);

CKINVDCx5p33_ASAP7_75t_R g4673 ( 
.A(n_1499),
.Y(n_4673)
);

INVx1_ASAP7_75t_SL g4674 ( 
.A(n_272),
.Y(n_4674)
);

CKINVDCx5p33_ASAP7_75t_R g4675 ( 
.A(n_2098),
.Y(n_4675)
);

CKINVDCx5p33_ASAP7_75t_R g4676 ( 
.A(n_2425),
.Y(n_4676)
);

CKINVDCx5p33_ASAP7_75t_R g4677 ( 
.A(n_2933),
.Y(n_4677)
);

CKINVDCx5p33_ASAP7_75t_R g4678 ( 
.A(n_1638),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_1026),
.Y(n_4679)
);

CKINVDCx5p33_ASAP7_75t_R g4680 ( 
.A(n_3607),
.Y(n_4680)
);

CKINVDCx20_ASAP7_75t_R g4681 ( 
.A(n_3923),
.Y(n_4681)
);

CKINVDCx5p33_ASAP7_75t_R g4682 ( 
.A(n_428),
.Y(n_4682)
);

CKINVDCx5p33_ASAP7_75t_R g4683 ( 
.A(n_253),
.Y(n_4683)
);

CKINVDCx5p33_ASAP7_75t_R g4684 ( 
.A(n_2318),
.Y(n_4684)
);

CKINVDCx5p33_ASAP7_75t_R g4685 ( 
.A(n_4073),
.Y(n_4685)
);

CKINVDCx5p33_ASAP7_75t_R g4686 ( 
.A(n_3913),
.Y(n_4686)
);

CKINVDCx5p33_ASAP7_75t_R g4687 ( 
.A(n_4057),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_2510),
.Y(n_4688)
);

CKINVDCx5p33_ASAP7_75t_R g4689 ( 
.A(n_2075),
.Y(n_4689)
);

CKINVDCx5p33_ASAP7_75t_R g4690 ( 
.A(n_1565),
.Y(n_4690)
);

CKINVDCx5p33_ASAP7_75t_R g4691 ( 
.A(n_2691),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_3054),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4030),
.Y(n_4693)
);

BUFx10_ASAP7_75t_L g4694 ( 
.A(n_1869),
.Y(n_4694)
);

CKINVDCx5p33_ASAP7_75t_R g4695 ( 
.A(n_990),
.Y(n_4695)
);

BUFx10_ASAP7_75t_L g4696 ( 
.A(n_3968),
.Y(n_4696)
);

INVx4_ASAP7_75t_R g4697 ( 
.A(n_4071),
.Y(n_4697)
);

CKINVDCx20_ASAP7_75t_R g4698 ( 
.A(n_919),
.Y(n_4698)
);

CKINVDCx5p33_ASAP7_75t_R g4699 ( 
.A(n_15),
.Y(n_4699)
);

CKINVDCx5p33_ASAP7_75t_R g4700 ( 
.A(n_1046),
.Y(n_4700)
);

CKINVDCx5p33_ASAP7_75t_R g4701 ( 
.A(n_935),
.Y(n_4701)
);

CKINVDCx20_ASAP7_75t_R g4702 ( 
.A(n_4020),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_2927),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_2806),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_293),
.Y(n_4705)
);

CKINVDCx5p33_ASAP7_75t_R g4706 ( 
.A(n_1729),
.Y(n_4706)
);

CKINVDCx5p33_ASAP7_75t_R g4707 ( 
.A(n_2744),
.Y(n_4707)
);

BUFx6f_ASAP7_75t_L g4708 ( 
.A(n_779),
.Y(n_4708)
);

CKINVDCx5p33_ASAP7_75t_R g4709 ( 
.A(n_1918),
.Y(n_4709)
);

BUFx8_ASAP7_75t_SL g4710 ( 
.A(n_3890),
.Y(n_4710)
);

CKINVDCx5p33_ASAP7_75t_R g4711 ( 
.A(n_3270),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_717),
.Y(n_4712)
);

XOR2xp5_ASAP7_75t_L g4713 ( 
.A(n_1141),
.B(n_2235),
.Y(n_4713)
);

CKINVDCx5p33_ASAP7_75t_R g4714 ( 
.A(n_912),
.Y(n_4714)
);

CKINVDCx5p33_ASAP7_75t_R g4715 ( 
.A(n_882),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_553),
.Y(n_4716)
);

CKINVDCx5p33_ASAP7_75t_R g4717 ( 
.A(n_4059),
.Y(n_4717)
);

CKINVDCx5p33_ASAP7_75t_R g4718 ( 
.A(n_3078),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_3965),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_2160),
.Y(n_4720)
);

BUFx10_ASAP7_75t_L g4721 ( 
.A(n_1522),
.Y(n_4721)
);

CKINVDCx5p33_ASAP7_75t_R g4722 ( 
.A(n_2584),
.Y(n_4722)
);

INVx1_ASAP7_75t_SL g4723 ( 
.A(n_1245),
.Y(n_4723)
);

CKINVDCx5p33_ASAP7_75t_R g4724 ( 
.A(n_879),
.Y(n_4724)
);

CKINVDCx5p33_ASAP7_75t_R g4725 ( 
.A(n_1010),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_2184),
.Y(n_4726)
);

BUFx3_ASAP7_75t_L g4727 ( 
.A(n_2619),
.Y(n_4727)
);

CKINVDCx5p33_ASAP7_75t_R g4728 ( 
.A(n_3779),
.Y(n_4728)
);

CKINVDCx5p33_ASAP7_75t_R g4729 ( 
.A(n_798),
.Y(n_4729)
);

CKINVDCx5p33_ASAP7_75t_R g4730 ( 
.A(n_2073),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_3592),
.Y(n_4731)
);

CKINVDCx5p33_ASAP7_75t_R g4732 ( 
.A(n_2885),
.Y(n_4732)
);

CKINVDCx5p33_ASAP7_75t_R g4733 ( 
.A(n_3941),
.Y(n_4733)
);

BUFx10_ASAP7_75t_L g4734 ( 
.A(n_28),
.Y(n_4734)
);

CKINVDCx5p33_ASAP7_75t_R g4735 ( 
.A(n_97),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_3139),
.Y(n_4736)
);

CKINVDCx5p33_ASAP7_75t_R g4737 ( 
.A(n_2085),
.Y(n_4737)
);

CKINVDCx5p33_ASAP7_75t_R g4738 ( 
.A(n_3442),
.Y(n_4738)
);

CKINVDCx5p33_ASAP7_75t_R g4739 ( 
.A(n_665),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_2714),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_1209),
.Y(n_4741)
);

CKINVDCx20_ASAP7_75t_R g4742 ( 
.A(n_1328),
.Y(n_4742)
);

CKINVDCx16_ASAP7_75t_R g4743 ( 
.A(n_985),
.Y(n_4743)
);

CKINVDCx5p33_ASAP7_75t_R g4744 ( 
.A(n_3769),
.Y(n_4744)
);

CKINVDCx5p33_ASAP7_75t_R g4745 ( 
.A(n_2923),
.Y(n_4745)
);

BUFx2_ASAP7_75t_L g4746 ( 
.A(n_3904),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_2666),
.Y(n_4747)
);

CKINVDCx20_ASAP7_75t_R g4748 ( 
.A(n_3364),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_3577),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_2627),
.Y(n_4750)
);

CKINVDCx5p33_ASAP7_75t_R g4751 ( 
.A(n_440),
.Y(n_4751)
);

BUFx5_ASAP7_75t_L g4752 ( 
.A(n_260),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_2953),
.Y(n_4753)
);

CKINVDCx5p33_ASAP7_75t_R g4754 ( 
.A(n_1302),
.Y(n_4754)
);

BUFx3_ASAP7_75t_L g4755 ( 
.A(n_1752),
.Y(n_4755)
);

BUFx6f_ASAP7_75t_L g4756 ( 
.A(n_3059),
.Y(n_4756)
);

BUFx10_ASAP7_75t_L g4757 ( 
.A(n_3942),
.Y(n_4757)
);

CKINVDCx5p33_ASAP7_75t_R g4758 ( 
.A(n_1136),
.Y(n_4758)
);

CKINVDCx5p33_ASAP7_75t_R g4759 ( 
.A(n_232),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_3321),
.Y(n_4760)
);

BUFx10_ASAP7_75t_L g4761 ( 
.A(n_4074),
.Y(n_4761)
);

CKINVDCx5p33_ASAP7_75t_R g4762 ( 
.A(n_3847),
.Y(n_4762)
);

CKINVDCx5p33_ASAP7_75t_R g4763 ( 
.A(n_3231),
.Y(n_4763)
);

CKINVDCx5p33_ASAP7_75t_R g4764 ( 
.A(n_2524),
.Y(n_4764)
);

HB1xp67_ASAP7_75t_L g4765 ( 
.A(n_2251),
.Y(n_4765)
);

CKINVDCx5p33_ASAP7_75t_R g4766 ( 
.A(n_483),
.Y(n_4766)
);

CKINVDCx5p33_ASAP7_75t_R g4767 ( 
.A(n_879),
.Y(n_4767)
);

INVxp67_ASAP7_75t_SL g4768 ( 
.A(n_4093),
.Y(n_4768)
);

CKINVDCx5p33_ASAP7_75t_R g4769 ( 
.A(n_4054),
.Y(n_4769)
);

BUFx2_ASAP7_75t_L g4770 ( 
.A(n_1215),
.Y(n_4770)
);

CKINVDCx5p33_ASAP7_75t_R g4771 ( 
.A(n_2431),
.Y(n_4771)
);

BUFx3_ASAP7_75t_L g4772 ( 
.A(n_3602),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_809),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4073),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_192),
.Y(n_4775)
);

CKINVDCx5p33_ASAP7_75t_R g4776 ( 
.A(n_2591),
.Y(n_4776)
);

CKINVDCx5p33_ASAP7_75t_R g4777 ( 
.A(n_2282),
.Y(n_4777)
);

CKINVDCx5p33_ASAP7_75t_R g4778 ( 
.A(n_1521),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_1435),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_3896),
.Y(n_4780)
);

CKINVDCx16_ASAP7_75t_R g4781 ( 
.A(n_1899),
.Y(n_4781)
);

CKINVDCx5p33_ASAP7_75t_R g4782 ( 
.A(n_353),
.Y(n_4782)
);

CKINVDCx5p33_ASAP7_75t_R g4783 ( 
.A(n_1264),
.Y(n_4783)
);

CKINVDCx5p33_ASAP7_75t_R g4784 ( 
.A(n_3733),
.Y(n_4784)
);

BUFx10_ASAP7_75t_L g4785 ( 
.A(n_4082),
.Y(n_4785)
);

CKINVDCx5p33_ASAP7_75t_R g4786 ( 
.A(n_486),
.Y(n_4786)
);

CKINVDCx5p33_ASAP7_75t_R g4787 ( 
.A(n_575),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_2166),
.Y(n_4788)
);

CKINVDCx5p33_ASAP7_75t_R g4789 ( 
.A(n_3466),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_3955),
.Y(n_4790)
);

CKINVDCx5p33_ASAP7_75t_R g4791 ( 
.A(n_4006),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_871),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_1529),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_776),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_3139),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_3708),
.Y(n_4796)
);

BUFx10_ASAP7_75t_L g4797 ( 
.A(n_3956),
.Y(n_4797)
);

CKINVDCx5p33_ASAP7_75t_R g4798 ( 
.A(n_1039),
.Y(n_4798)
);

INVx1_ASAP7_75t_SL g4799 ( 
.A(n_1004),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_486),
.Y(n_4800)
);

CKINVDCx5p33_ASAP7_75t_R g4801 ( 
.A(n_3230),
.Y(n_4801)
);

CKINVDCx5p33_ASAP7_75t_R g4802 ( 
.A(n_3884),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_3989),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_2565),
.Y(n_4804)
);

CKINVDCx5p33_ASAP7_75t_R g4805 ( 
.A(n_1427),
.Y(n_4805)
);

CKINVDCx5p33_ASAP7_75t_R g4806 ( 
.A(n_3618),
.Y(n_4806)
);

CKINVDCx5p33_ASAP7_75t_R g4807 ( 
.A(n_1703),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_659),
.Y(n_4808)
);

CKINVDCx5p33_ASAP7_75t_R g4809 ( 
.A(n_3648),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_3581),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_49),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_1314),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_2462),
.Y(n_4813)
);

CKINVDCx20_ASAP7_75t_R g4814 ( 
.A(n_3951),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_3022),
.Y(n_4815)
);

INVxp67_ASAP7_75t_L g4816 ( 
.A(n_3818),
.Y(n_4816)
);

CKINVDCx5p33_ASAP7_75t_R g4817 ( 
.A(n_534),
.Y(n_4817)
);

CKINVDCx5p33_ASAP7_75t_R g4818 ( 
.A(n_3365),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_2288),
.Y(n_4819)
);

CKINVDCx5p33_ASAP7_75t_R g4820 ( 
.A(n_4027),
.Y(n_4820)
);

CKINVDCx5p33_ASAP7_75t_R g4821 ( 
.A(n_284),
.Y(n_4821)
);

CKINVDCx16_ASAP7_75t_R g4822 ( 
.A(n_1404),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_3769),
.Y(n_4823)
);

INVxp67_ASAP7_75t_L g4824 ( 
.A(n_311),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4026),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_1213),
.Y(n_4826)
);

CKINVDCx5p33_ASAP7_75t_R g4827 ( 
.A(n_4042),
.Y(n_4827)
);

HB1xp67_ASAP7_75t_L g4828 ( 
.A(n_1520),
.Y(n_4828)
);

CKINVDCx5p33_ASAP7_75t_R g4829 ( 
.A(n_2053),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_3364),
.Y(n_4830)
);

CKINVDCx20_ASAP7_75t_R g4831 ( 
.A(n_3162),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_2114),
.Y(n_4832)
);

CKINVDCx5p33_ASAP7_75t_R g4833 ( 
.A(n_4050),
.Y(n_4833)
);

CKINVDCx14_ASAP7_75t_R g4834 ( 
.A(n_553),
.Y(n_4834)
);

CKINVDCx5p33_ASAP7_75t_R g4835 ( 
.A(n_754),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_393),
.Y(n_4836)
);

BUFx10_ASAP7_75t_L g4837 ( 
.A(n_2842),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_2785),
.Y(n_4838)
);

CKINVDCx5p33_ASAP7_75t_R g4839 ( 
.A(n_2807),
.Y(n_4839)
);

CKINVDCx5p33_ASAP7_75t_R g4840 ( 
.A(n_3931),
.Y(n_4840)
);

INVx2_ASAP7_75t_L g4841 ( 
.A(n_1596),
.Y(n_4841)
);

CKINVDCx5p33_ASAP7_75t_R g4842 ( 
.A(n_970),
.Y(n_4842)
);

INVx1_ASAP7_75t_SL g4843 ( 
.A(n_3814),
.Y(n_4843)
);

CKINVDCx5p33_ASAP7_75t_R g4844 ( 
.A(n_3312),
.Y(n_4844)
);

CKINVDCx5p33_ASAP7_75t_R g4845 ( 
.A(n_9),
.Y(n_4845)
);

CKINVDCx5p33_ASAP7_75t_R g4846 ( 
.A(n_1120),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_1741),
.Y(n_4847)
);

INVx1_ASAP7_75t_SL g4848 ( 
.A(n_70),
.Y(n_4848)
);

CKINVDCx16_ASAP7_75t_R g4849 ( 
.A(n_3934),
.Y(n_4849)
);

CKINVDCx5p33_ASAP7_75t_R g4850 ( 
.A(n_2899),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_166),
.Y(n_4851)
);

CKINVDCx20_ASAP7_75t_R g4852 ( 
.A(n_2830),
.Y(n_4852)
);

CKINVDCx20_ASAP7_75t_R g4853 ( 
.A(n_1647),
.Y(n_4853)
);

CKINVDCx5p33_ASAP7_75t_R g4854 ( 
.A(n_656),
.Y(n_4854)
);

CKINVDCx5p33_ASAP7_75t_R g4855 ( 
.A(n_432),
.Y(n_4855)
);

CKINVDCx5p33_ASAP7_75t_R g4856 ( 
.A(n_64),
.Y(n_4856)
);

INVx1_ASAP7_75t_SL g4857 ( 
.A(n_4027),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_3970),
.Y(n_4858)
);

CKINVDCx5p33_ASAP7_75t_R g4859 ( 
.A(n_3396),
.Y(n_4859)
);

CKINVDCx5p33_ASAP7_75t_R g4860 ( 
.A(n_459),
.Y(n_4860)
);

CKINVDCx5p33_ASAP7_75t_R g4861 ( 
.A(n_1132),
.Y(n_4861)
);

CKINVDCx5p33_ASAP7_75t_R g4862 ( 
.A(n_3548),
.Y(n_4862)
);

CKINVDCx5p33_ASAP7_75t_R g4863 ( 
.A(n_2301),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_2721),
.Y(n_4864)
);

CKINVDCx5p33_ASAP7_75t_R g4865 ( 
.A(n_10),
.Y(n_4865)
);

INVx2_ASAP7_75t_L g4866 ( 
.A(n_4066),
.Y(n_4866)
);

CKINVDCx5p33_ASAP7_75t_R g4867 ( 
.A(n_225),
.Y(n_4867)
);

CKINVDCx5p33_ASAP7_75t_R g4868 ( 
.A(n_252),
.Y(n_4868)
);

BUFx3_ASAP7_75t_L g4869 ( 
.A(n_580),
.Y(n_4869)
);

CKINVDCx20_ASAP7_75t_R g4870 ( 
.A(n_2035),
.Y(n_4870)
);

CKINVDCx5p33_ASAP7_75t_R g4871 ( 
.A(n_2999),
.Y(n_4871)
);

INVx1_ASAP7_75t_SL g4872 ( 
.A(n_336),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_3289),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_2419),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_3350),
.Y(n_4875)
);

CKINVDCx16_ASAP7_75t_R g4876 ( 
.A(n_3954),
.Y(n_4876)
);

CKINVDCx20_ASAP7_75t_R g4877 ( 
.A(n_4076),
.Y(n_4877)
);

CKINVDCx5p33_ASAP7_75t_R g4878 ( 
.A(n_1512),
.Y(n_4878)
);

CKINVDCx5p33_ASAP7_75t_R g4879 ( 
.A(n_2801),
.Y(n_4879)
);

CKINVDCx5p33_ASAP7_75t_R g4880 ( 
.A(n_557),
.Y(n_4880)
);

CKINVDCx20_ASAP7_75t_R g4881 ( 
.A(n_3922),
.Y(n_4881)
);

CKINVDCx5p33_ASAP7_75t_R g4882 ( 
.A(n_3361),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_3210),
.Y(n_4883)
);

BUFx2_ASAP7_75t_L g4884 ( 
.A(n_2974),
.Y(n_4884)
);

BUFx10_ASAP7_75t_L g4885 ( 
.A(n_2757),
.Y(n_4885)
);

INVx2_ASAP7_75t_L g4886 ( 
.A(n_1323),
.Y(n_4886)
);

INVx1_ASAP7_75t_SL g4887 ( 
.A(n_1890),
.Y(n_4887)
);

CKINVDCx5p33_ASAP7_75t_R g4888 ( 
.A(n_3894),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4030),
.Y(n_4889)
);

BUFx10_ASAP7_75t_L g4890 ( 
.A(n_3900),
.Y(n_4890)
);

INVx1_ASAP7_75t_L g4891 ( 
.A(n_3583),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_3745),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_2877),
.Y(n_4893)
);

BUFx10_ASAP7_75t_L g4894 ( 
.A(n_188),
.Y(n_4894)
);

CKINVDCx5p33_ASAP7_75t_R g4895 ( 
.A(n_3513),
.Y(n_4895)
);

CKINVDCx5p33_ASAP7_75t_R g4896 ( 
.A(n_853),
.Y(n_4896)
);

BUFx10_ASAP7_75t_L g4897 ( 
.A(n_2782),
.Y(n_4897)
);

INVxp67_ASAP7_75t_L g4898 ( 
.A(n_4081),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_3654),
.Y(n_4899)
);

INVx2_ASAP7_75t_L g4900 ( 
.A(n_3542),
.Y(n_4900)
);

INVx2_ASAP7_75t_L g4901 ( 
.A(n_1996),
.Y(n_4901)
);

BUFx3_ASAP7_75t_L g4902 ( 
.A(n_1164),
.Y(n_4902)
);

CKINVDCx5p33_ASAP7_75t_R g4903 ( 
.A(n_778),
.Y(n_4903)
);

INVx1_ASAP7_75t_SL g4904 ( 
.A(n_364),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4101),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_2725),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_1997),
.Y(n_4907)
);

CKINVDCx5p33_ASAP7_75t_R g4908 ( 
.A(n_1099),
.Y(n_4908)
);

CKINVDCx5p33_ASAP7_75t_R g4909 ( 
.A(n_3916),
.Y(n_4909)
);

CKINVDCx5p33_ASAP7_75t_R g4910 ( 
.A(n_3981),
.Y(n_4910)
);

CKINVDCx20_ASAP7_75t_R g4911 ( 
.A(n_2674),
.Y(n_4911)
);

CKINVDCx5p33_ASAP7_75t_R g4912 ( 
.A(n_2379),
.Y(n_4912)
);

CKINVDCx5p33_ASAP7_75t_R g4913 ( 
.A(n_481),
.Y(n_4913)
);

CKINVDCx5p33_ASAP7_75t_R g4914 ( 
.A(n_2995),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_958),
.Y(n_4915)
);

CKINVDCx5p33_ASAP7_75t_R g4916 ( 
.A(n_2879),
.Y(n_4916)
);

INVx2_ASAP7_75t_SL g4917 ( 
.A(n_651),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_146),
.Y(n_4918)
);

HB1xp67_ASAP7_75t_L g4919 ( 
.A(n_589),
.Y(n_4919)
);

CKINVDCx20_ASAP7_75t_R g4920 ( 
.A(n_14),
.Y(n_4920)
);

CKINVDCx5p33_ASAP7_75t_R g4921 ( 
.A(n_31),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_1567),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_354),
.Y(n_4923)
);

INVx2_ASAP7_75t_SL g4924 ( 
.A(n_1288),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_3143),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_1516),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_419),
.Y(n_4927)
);

CKINVDCx5p33_ASAP7_75t_R g4928 ( 
.A(n_2101),
.Y(n_4928)
);

BUFx3_ASAP7_75t_L g4929 ( 
.A(n_2868),
.Y(n_4929)
);

CKINVDCx5p33_ASAP7_75t_R g4930 ( 
.A(n_3722),
.Y(n_4930)
);

CKINVDCx20_ASAP7_75t_R g4931 ( 
.A(n_3973),
.Y(n_4931)
);

CKINVDCx5p33_ASAP7_75t_R g4932 ( 
.A(n_443),
.Y(n_4932)
);

CKINVDCx20_ASAP7_75t_R g4933 ( 
.A(n_1467),
.Y(n_4933)
);

CKINVDCx5p33_ASAP7_75t_R g4934 ( 
.A(n_357),
.Y(n_4934)
);

CKINVDCx5p33_ASAP7_75t_R g4935 ( 
.A(n_827),
.Y(n_4935)
);

INVx2_ASAP7_75t_SL g4936 ( 
.A(n_3987),
.Y(n_4936)
);

CKINVDCx20_ASAP7_75t_R g4937 ( 
.A(n_805),
.Y(n_4937)
);

CKINVDCx5p33_ASAP7_75t_R g4938 ( 
.A(n_2873),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_1663),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_3244),
.Y(n_4940)
);

CKINVDCx20_ASAP7_75t_R g4941 ( 
.A(n_4046),
.Y(n_4941)
);

CKINVDCx5p33_ASAP7_75t_R g4942 ( 
.A(n_1149),
.Y(n_4942)
);

CKINVDCx5p33_ASAP7_75t_R g4943 ( 
.A(n_3114),
.Y(n_4943)
);

BUFx6f_ASAP7_75t_L g4944 ( 
.A(n_1779),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_2335),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_3854),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_936),
.Y(n_4947)
);

BUFx10_ASAP7_75t_L g4948 ( 
.A(n_3249),
.Y(n_4948)
);

CKINVDCx5p33_ASAP7_75t_R g4949 ( 
.A(n_4087),
.Y(n_4949)
);

INVx1_ASAP7_75t_SL g4950 ( 
.A(n_4049),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_119),
.Y(n_4951)
);

CKINVDCx5p33_ASAP7_75t_R g4952 ( 
.A(n_1784),
.Y(n_4952)
);

INVx2_ASAP7_75t_L g4953 ( 
.A(n_1488),
.Y(n_4953)
);

BUFx2_ASAP7_75t_L g4954 ( 
.A(n_574),
.Y(n_4954)
);

INVxp67_ASAP7_75t_L g4955 ( 
.A(n_1838),
.Y(n_4955)
);

INVxp67_ASAP7_75t_SL g4956 ( 
.A(n_4019),
.Y(n_4956)
);

CKINVDCx5p33_ASAP7_75t_R g4957 ( 
.A(n_1669),
.Y(n_4957)
);

CKINVDCx5p33_ASAP7_75t_R g4958 ( 
.A(n_1802),
.Y(n_4958)
);

CKINVDCx5p33_ASAP7_75t_R g4959 ( 
.A(n_586),
.Y(n_4959)
);

CKINVDCx5p33_ASAP7_75t_R g4960 ( 
.A(n_1237),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_2500),
.Y(n_4961)
);

CKINVDCx5p33_ASAP7_75t_R g4962 ( 
.A(n_2562),
.Y(n_4962)
);

CKINVDCx5p33_ASAP7_75t_R g4963 ( 
.A(n_4017),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_1391),
.Y(n_4964)
);

CKINVDCx5p33_ASAP7_75t_R g4965 ( 
.A(n_2337),
.Y(n_4965)
);

CKINVDCx20_ASAP7_75t_R g4966 ( 
.A(n_2819),
.Y(n_4966)
);

CKINVDCx5p33_ASAP7_75t_R g4967 ( 
.A(n_3544),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_1790),
.Y(n_4968)
);

CKINVDCx14_ASAP7_75t_R g4969 ( 
.A(n_1391),
.Y(n_4969)
);

CKINVDCx5p33_ASAP7_75t_R g4970 ( 
.A(n_1203),
.Y(n_4970)
);

BUFx6f_ASAP7_75t_L g4971 ( 
.A(n_2637),
.Y(n_4971)
);

CKINVDCx5p33_ASAP7_75t_R g4972 ( 
.A(n_4040),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_634),
.Y(n_4973)
);

CKINVDCx5p33_ASAP7_75t_R g4974 ( 
.A(n_4018),
.Y(n_4974)
);

CKINVDCx5p33_ASAP7_75t_R g4975 ( 
.A(n_420),
.Y(n_4975)
);

BUFx3_ASAP7_75t_L g4976 ( 
.A(n_84),
.Y(n_4976)
);

CKINVDCx16_ASAP7_75t_R g4977 ( 
.A(n_3926),
.Y(n_4977)
);

CKINVDCx5p33_ASAP7_75t_R g4978 ( 
.A(n_2548),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_3979),
.Y(n_4979)
);

CKINVDCx5p33_ASAP7_75t_R g4980 ( 
.A(n_4005),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_132),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_1060),
.Y(n_4982)
);

CKINVDCx5p33_ASAP7_75t_R g4983 ( 
.A(n_71),
.Y(n_4983)
);

CKINVDCx5p33_ASAP7_75t_R g4984 ( 
.A(n_3919),
.Y(n_4984)
);

CKINVDCx20_ASAP7_75t_R g4985 ( 
.A(n_2811),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_1690),
.Y(n_4986)
);

CKINVDCx5p33_ASAP7_75t_R g4987 ( 
.A(n_2220),
.Y(n_4987)
);

CKINVDCx5p33_ASAP7_75t_R g4988 ( 
.A(n_1574),
.Y(n_4988)
);

BUFx10_ASAP7_75t_L g4989 ( 
.A(n_3458),
.Y(n_4989)
);

INVx2_ASAP7_75t_SL g4990 ( 
.A(n_1930),
.Y(n_4990)
);

CKINVDCx5p33_ASAP7_75t_R g4991 ( 
.A(n_98),
.Y(n_4991)
);

CKINVDCx5p33_ASAP7_75t_R g4992 ( 
.A(n_748),
.Y(n_4992)
);

INVx3_ASAP7_75t_L g4993 ( 
.A(n_3341),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_3716),
.Y(n_4994)
);

CKINVDCx5p33_ASAP7_75t_R g4995 ( 
.A(n_33),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_347),
.Y(n_4996)
);

CKINVDCx14_ASAP7_75t_R g4997 ( 
.A(n_2485),
.Y(n_4997)
);

CKINVDCx5p33_ASAP7_75t_R g4998 ( 
.A(n_767),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_1935),
.Y(n_4999)
);

CKINVDCx5p33_ASAP7_75t_R g5000 ( 
.A(n_4088),
.Y(n_5000)
);

CKINVDCx5p33_ASAP7_75t_R g5001 ( 
.A(n_1369),
.Y(n_5001)
);

CKINVDCx5p33_ASAP7_75t_R g5002 ( 
.A(n_1953),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_143),
.Y(n_5003)
);

CKINVDCx5p33_ASAP7_75t_R g5004 ( 
.A(n_4070),
.Y(n_5004)
);

CKINVDCx5p33_ASAP7_75t_R g5005 ( 
.A(n_1138),
.Y(n_5005)
);

BUFx2_ASAP7_75t_L g5006 ( 
.A(n_1529),
.Y(n_5006)
);

INVxp67_ASAP7_75t_L g5007 ( 
.A(n_965),
.Y(n_5007)
);

BUFx2_ASAP7_75t_SL g5008 ( 
.A(n_143),
.Y(n_5008)
);

CKINVDCx5p33_ASAP7_75t_R g5009 ( 
.A(n_826),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_2334),
.Y(n_5010)
);

CKINVDCx5p33_ASAP7_75t_R g5011 ( 
.A(n_1218),
.Y(n_5011)
);

CKINVDCx5p33_ASAP7_75t_R g5012 ( 
.A(n_3138),
.Y(n_5012)
);

CKINVDCx5p33_ASAP7_75t_R g5013 ( 
.A(n_3479),
.Y(n_5013)
);

CKINVDCx16_ASAP7_75t_R g5014 ( 
.A(n_1031),
.Y(n_5014)
);

CKINVDCx5p33_ASAP7_75t_R g5015 ( 
.A(n_457),
.Y(n_5015)
);

BUFx2_ASAP7_75t_R g5016 ( 
.A(n_1637),
.Y(n_5016)
);

CKINVDCx5p33_ASAP7_75t_R g5017 ( 
.A(n_3646),
.Y(n_5017)
);

BUFx2_ASAP7_75t_SL g5018 ( 
.A(n_2801),
.Y(n_5018)
);

INVx1_ASAP7_75t_SL g5019 ( 
.A(n_3172),
.Y(n_5019)
);

CKINVDCx20_ASAP7_75t_R g5020 ( 
.A(n_3967),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_2155),
.Y(n_5021)
);

CKINVDCx5p33_ASAP7_75t_R g5022 ( 
.A(n_3184),
.Y(n_5022)
);

CKINVDCx5p33_ASAP7_75t_R g5023 ( 
.A(n_2492),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_3178),
.Y(n_5024)
);

CKINVDCx5p33_ASAP7_75t_R g5025 ( 
.A(n_3962),
.Y(n_5025)
);

INVx1_ASAP7_75t_SL g5026 ( 
.A(n_2985),
.Y(n_5026)
);

BUFx2_ASAP7_75t_L g5027 ( 
.A(n_3956),
.Y(n_5027)
);

CKINVDCx5p33_ASAP7_75t_R g5028 ( 
.A(n_2726),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_2576),
.Y(n_5029)
);

CKINVDCx5p33_ASAP7_75t_R g5030 ( 
.A(n_3921),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_2925),
.Y(n_5031)
);

CKINVDCx5p33_ASAP7_75t_R g5032 ( 
.A(n_3616),
.Y(n_5032)
);

CKINVDCx5p33_ASAP7_75t_R g5033 ( 
.A(n_57),
.Y(n_5033)
);

CKINVDCx5p33_ASAP7_75t_R g5034 ( 
.A(n_3370),
.Y(n_5034)
);

CKINVDCx5p33_ASAP7_75t_R g5035 ( 
.A(n_2144),
.Y(n_5035)
);

CKINVDCx5p33_ASAP7_75t_R g5036 ( 
.A(n_2215),
.Y(n_5036)
);

CKINVDCx20_ASAP7_75t_R g5037 ( 
.A(n_1834),
.Y(n_5037)
);

HB1xp67_ASAP7_75t_L g5038 ( 
.A(n_347),
.Y(n_5038)
);

CKINVDCx20_ASAP7_75t_R g5039 ( 
.A(n_170),
.Y(n_5039)
);

CKINVDCx5p33_ASAP7_75t_R g5040 ( 
.A(n_2723),
.Y(n_5040)
);

CKINVDCx5p33_ASAP7_75t_R g5041 ( 
.A(n_1854),
.Y(n_5041)
);

CKINVDCx5p33_ASAP7_75t_R g5042 ( 
.A(n_2494),
.Y(n_5042)
);

INVx2_ASAP7_75t_SL g5043 ( 
.A(n_2330),
.Y(n_5043)
);

BUFx5_ASAP7_75t_L g5044 ( 
.A(n_1985),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_1630),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_2328),
.Y(n_5046)
);

INVx1_ASAP7_75t_SL g5047 ( 
.A(n_3334),
.Y(n_5047)
);

CKINVDCx5p33_ASAP7_75t_R g5048 ( 
.A(n_1877),
.Y(n_5048)
);

CKINVDCx5p33_ASAP7_75t_R g5049 ( 
.A(n_2199),
.Y(n_5049)
);

CKINVDCx5p33_ASAP7_75t_R g5050 ( 
.A(n_2330),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_2239),
.Y(n_5051)
);

CKINVDCx5p33_ASAP7_75t_R g5052 ( 
.A(n_3245),
.Y(n_5052)
);

CKINVDCx20_ASAP7_75t_R g5053 ( 
.A(n_2753),
.Y(n_5053)
);

BUFx6f_ASAP7_75t_L g5054 ( 
.A(n_3337),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_2766),
.Y(n_5055)
);

INVxp67_ASAP7_75t_SL g5056 ( 
.A(n_3906),
.Y(n_5056)
);

CKINVDCx5p33_ASAP7_75t_R g5057 ( 
.A(n_1991),
.Y(n_5057)
);

CKINVDCx20_ASAP7_75t_R g5058 ( 
.A(n_1942),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_40),
.Y(n_5059)
);

INVx1_ASAP7_75t_SL g5060 ( 
.A(n_555),
.Y(n_5060)
);

CKINVDCx5p33_ASAP7_75t_R g5061 ( 
.A(n_1166),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_2087),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_2374),
.Y(n_5063)
);

CKINVDCx5p33_ASAP7_75t_R g5064 ( 
.A(n_1223),
.Y(n_5064)
);

CKINVDCx5p33_ASAP7_75t_R g5065 ( 
.A(n_1775),
.Y(n_5065)
);

CKINVDCx5p33_ASAP7_75t_R g5066 ( 
.A(n_2368),
.Y(n_5066)
);

CKINVDCx5p33_ASAP7_75t_R g5067 ( 
.A(n_3271),
.Y(n_5067)
);

BUFx10_ASAP7_75t_L g5068 ( 
.A(n_3128),
.Y(n_5068)
);

CKINVDCx5p33_ASAP7_75t_R g5069 ( 
.A(n_1258),
.Y(n_5069)
);

CKINVDCx5p33_ASAP7_75t_R g5070 ( 
.A(n_2644),
.Y(n_5070)
);

BUFx3_ASAP7_75t_L g5071 ( 
.A(n_3911),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_2284),
.Y(n_5072)
);

CKINVDCx16_ASAP7_75t_R g5073 ( 
.A(n_2670),
.Y(n_5073)
);

CKINVDCx5p33_ASAP7_75t_R g5074 ( 
.A(n_3905),
.Y(n_5074)
);

CKINVDCx16_ASAP7_75t_R g5075 ( 
.A(n_3557),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_1627),
.Y(n_5076)
);

CKINVDCx5p33_ASAP7_75t_R g5077 ( 
.A(n_2379),
.Y(n_5077)
);

CKINVDCx5p33_ASAP7_75t_R g5078 ( 
.A(n_3845),
.Y(n_5078)
);

CKINVDCx5p33_ASAP7_75t_R g5079 ( 
.A(n_381),
.Y(n_5079)
);

CKINVDCx5p33_ASAP7_75t_R g5080 ( 
.A(n_3032),
.Y(n_5080)
);

INVx2_ASAP7_75t_L g5081 ( 
.A(n_1249),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_304),
.Y(n_5082)
);

CKINVDCx5p33_ASAP7_75t_R g5083 ( 
.A(n_933),
.Y(n_5083)
);

CKINVDCx20_ASAP7_75t_R g5084 ( 
.A(n_4004),
.Y(n_5084)
);

CKINVDCx5p33_ASAP7_75t_R g5085 ( 
.A(n_3366),
.Y(n_5085)
);

INVx1_ASAP7_75t_SL g5086 ( 
.A(n_3425),
.Y(n_5086)
);

CKINVDCx5p33_ASAP7_75t_R g5087 ( 
.A(n_1850),
.Y(n_5087)
);

CKINVDCx20_ASAP7_75t_R g5088 ( 
.A(n_3810),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_1073),
.Y(n_5089)
);

CKINVDCx5p33_ASAP7_75t_R g5090 ( 
.A(n_3963),
.Y(n_5090)
);

CKINVDCx5p33_ASAP7_75t_R g5091 ( 
.A(n_4061),
.Y(n_5091)
);

CKINVDCx5p33_ASAP7_75t_R g5092 ( 
.A(n_1175),
.Y(n_5092)
);

INVx2_ASAP7_75t_SL g5093 ( 
.A(n_3222),
.Y(n_5093)
);

CKINVDCx5p33_ASAP7_75t_R g5094 ( 
.A(n_3396),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_745),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_741),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_3903),
.Y(n_5097)
);

CKINVDCx5p33_ASAP7_75t_R g5098 ( 
.A(n_3099),
.Y(n_5098)
);

BUFx2_ASAP7_75t_L g5099 ( 
.A(n_2955),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_3480),
.Y(n_5100)
);

CKINVDCx16_ASAP7_75t_R g5101 ( 
.A(n_39),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_1498),
.Y(n_5102)
);

INVx2_ASAP7_75t_L g5103 ( 
.A(n_3262),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_3708),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_1574),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_3146),
.Y(n_5106)
);

CKINVDCx5p33_ASAP7_75t_R g5107 ( 
.A(n_3347),
.Y(n_5107)
);

BUFx2_ASAP7_75t_L g5108 ( 
.A(n_3106),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_632),
.Y(n_5109)
);

CKINVDCx5p33_ASAP7_75t_R g5110 ( 
.A(n_3940),
.Y(n_5110)
);

CKINVDCx14_ASAP7_75t_R g5111 ( 
.A(n_4063),
.Y(n_5111)
);

CKINVDCx5p33_ASAP7_75t_R g5112 ( 
.A(n_2445),
.Y(n_5112)
);

CKINVDCx5p33_ASAP7_75t_R g5113 ( 
.A(n_2953),
.Y(n_5113)
);

CKINVDCx5p33_ASAP7_75t_R g5114 ( 
.A(n_1011),
.Y(n_5114)
);

CKINVDCx5p33_ASAP7_75t_R g5115 ( 
.A(n_3759),
.Y(n_5115)
);

INVx2_ASAP7_75t_SL g5116 ( 
.A(n_1740),
.Y(n_5116)
);

CKINVDCx5p33_ASAP7_75t_R g5117 ( 
.A(n_2802),
.Y(n_5117)
);

CKINVDCx5p33_ASAP7_75t_R g5118 ( 
.A(n_3475),
.Y(n_5118)
);

BUFx6f_ASAP7_75t_L g5119 ( 
.A(n_2224),
.Y(n_5119)
);

INVx1_ASAP7_75t_SL g5120 ( 
.A(n_2107),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_2394),
.Y(n_5121)
);

CKINVDCx5p33_ASAP7_75t_R g5122 ( 
.A(n_3247),
.Y(n_5122)
);

CKINVDCx5p33_ASAP7_75t_R g5123 ( 
.A(n_1876),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_1953),
.Y(n_5124)
);

CKINVDCx5p33_ASAP7_75t_R g5125 ( 
.A(n_2605),
.Y(n_5125)
);

CKINVDCx5p33_ASAP7_75t_R g5126 ( 
.A(n_3589),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_4044),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_1187),
.Y(n_5128)
);

INVx2_ASAP7_75t_L g5129 ( 
.A(n_2741),
.Y(n_5129)
);

CKINVDCx5p33_ASAP7_75t_R g5130 ( 
.A(n_220),
.Y(n_5130)
);

CKINVDCx5p33_ASAP7_75t_R g5131 ( 
.A(n_3933),
.Y(n_5131)
);

CKINVDCx5p33_ASAP7_75t_R g5132 ( 
.A(n_1286),
.Y(n_5132)
);

CKINVDCx5p33_ASAP7_75t_R g5133 ( 
.A(n_2679),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_1776),
.Y(n_5134)
);

CKINVDCx5p33_ASAP7_75t_R g5135 ( 
.A(n_1914),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_280),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_1013),
.Y(n_5137)
);

CKINVDCx5p33_ASAP7_75t_R g5138 ( 
.A(n_2597),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_3915),
.Y(n_5139)
);

INVx2_ASAP7_75t_L g5140 ( 
.A(n_3011),
.Y(n_5140)
);

CKINVDCx5p33_ASAP7_75t_R g5141 ( 
.A(n_1636),
.Y(n_5141)
);

CKINVDCx20_ASAP7_75t_R g5142 ( 
.A(n_84),
.Y(n_5142)
);

CKINVDCx20_ASAP7_75t_R g5143 ( 
.A(n_2378),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_1359),
.Y(n_5144)
);

CKINVDCx5p33_ASAP7_75t_R g5145 ( 
.A(n_3666),
.Y(n_5145)
);

INVx1_ASAP7_75t_SL g5146 ( 
.A(n_525),
.Y(n_5146)
);

BUFx10_ASAP7_75t_L g5147 ( 
.A(n_1752),
.Y(n_5147)
);

CKINVDCx5p33_ASAP7_75t_R g5148 ( 
.A(n_559),
.Y(n_5148)
);

CKINVDCx5p33_ASAP7_75t_R g5149 ( 
.A(n_2890),
.Y(n_5149)
);

CKINVDCx20_ASAP7_75t_R g5150 ( 
.A(n_757),
.Y(n_5150)
);

CKINVDCx5p33_ASAP7_75t_R g5151 ( 
.A(n_2733),
.Y(n_5151)
);

BUFx6f_ASAP7_75t_L g5152 ( 
.A(n_820),
.Y(n_5152)
);

CKINVDCx5p33_ASAP7_75t_R g5153 ( 
.A(n_1110),
.Y(n_5153)
);

CKINVDCx5p33_ASAP7_75t_R g5154 ( 
.A(n_649),
.Y(n_5154)
);

CKINVDCx5p33_ASAP7_75t_R g5155 ( 
.A(n_3697),
.Y(n_5155)
);

BUFx6f_ASAP7_75t_L g5156 ( 
.A(n_3214),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_3231),
.Y(n_5157)
);

CKINVDCx20_ASAP7_75t_R g5158 ( 
.A(n_3998),
.Y(n_5158)
);

CKINVDCx5p33_ASAP7_75t_R g5159 ( 
.A(n_406),
.Y(n_5159)
);

CKINVDCx5p33_ASAP7_75t_R g5160 ( 
.A(n_313),
.Y(n_5160)
);

CKINVDCx5p33_ASAP7_75t_R g5161 ( 
.A(n_2609),
.Y(n_5161)
);

CKINVDCx5p33_ASAP7_75t_R g5162 ( 
.A(n_4060),
.Y(n_5162)
);

INVx2_ASAP7_75t_L g5163 ( 
.A(n_2944),
.Y(n_5163)
);

CKINVDCx5p33_ASAP7_75t_R g5164 ( 
.A(n_209),
.Y(n_5164)
);

CKINVDCx20_ASAP7_75t_R g5165 ( 
.A(n_3562),
.Y(n_5165)
);

CKINVDCx5p33_ASAP7_75t_R g5166 ( 
.A(n_2452),
.Y(n_5166)
);

INVx2_ASAP7_75t_L g5167 ( 
.A(n_1947),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_2148),
.Y(n_5168)
);

CKINVDCx5p33_ASAP7_75t_R g5169 ( 
.A(n_2462),
.Y(n_5169)
);

CKINVDCx20_ASAP7_75t_R g5170 ( 
.A(n_3908),
.Y(n_5170)
);

CKINVDCx5p33_ASAP7_75t_R g5171 ( 
.A(n_3390),
.Y(n_5171)
);

BUFx3_ASAP7_75t_L g5172 ( 
.A(n_2319),
.Y(n_5172)
);

CKINVDCx5p33_ASAP7_75t_R g5173 ( 
.A(n_262),
.Y(n_5173)
);

INVx2_ASAP7_75t_L g5174 ( 
.A(n_431),
.Y(n_5174)
);

BUFx6f_ASAP7_75t_L g5175 ( 
.A(n_774),
.Y(n_5175)
);

CKINVDCx5p33_ASAP7_75t_R g5176 ( 
.A(n_1597),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4092),
.Y(n_5177)
);

INVx1_ASAP7_75t_SL g5178 ( 
.A(n_823),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_4070),
.Y(n_5179)
);

CKINVDCx5p33_ASAP7_75t_R g5180 ( 
.A(n_3902),
.Y(n_5180)
);

CKINVDCx5p33_ASAP7_75t_R g5181 ( 
.A(n_2021),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_4034),
.Y(n_5182)
);

CKINVDCx5p33_ASAP7_75t_R g5183 ( 
.A(n_1606),
.Y(n_5183)
);

INVxp67_ASAP7_75t_SL g5184 ( 
.A(n_666),
.Y(n_5184)
);

CKINVDCx5p33_ASAP7_75t_R g5185 ( 
.A(n_2407),
.Y(n_5185)
);

CKINVDCx5p33_ASAP7_75t_R g5186 ( 
.A(n_3453),
.Y(n_5186)
);

CKINVDCx5p33_ASAP7_75t_R g5187 ( 
.A(n_468),
.Y(n_5187)
);

CKINVDCx14_ASAP7_75t_R g5188 ( 
.A(n_538),
.Y(n_5188)
);

BUFx2_ASAP7_75t_L g5189 ( 
.A(n_3947),
.Y(n_5189)
);

CKINVDCx5p33_ASAP7_75t_R g5190 ( 
.A(n_3848),
.Y(n_5190)
);

CKINVDCx5p33_ASAP7_75t_R g5191 ( 
.A(n_3590),
.Y(n_5191)
);

INVx2_ASAP7_75t_L g5192 ( 
.A(n_1833),
.Y(n_5192)
);

CKINVDCx5p33_ASAP7_75t_R g5193 ( 
.A(n_3743),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_1219),
.Y(n_5194)
);

CKINVDCx5p33_ASAP7_75t_R g5195 ( 
.A(n_763),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_3125),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4078),
.Y(n_5197)
);

CKINVDCx16_ASAP7_75t_R g5198 ( 
.A(n_988),
.Y(n_5198)
);

CKINVDCx20_ASAP7_75t_R g5199 ( 
.A(n_4024),
.Y(n_5199)
);

CKINVDCx5p33_ASAP7_75t_R g5200 ( 
.A(n_917),
.Y(n_5200)
);

CKINVDCx5p33_ASAP7_75t_R g5201 ( 
.A(n_881),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_320),
.Y(n_5202)
);

BUFx10_ASAP7_75t_L g5203 ( 
.A(n_2434),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_2257),
.Y(n_5204)
);

CKINVDCx5p33_ASAP7_75t_R g5205 ( 
.A(n_3918),
.Y(n_5205)
);

CKINVDCx20_ASAP7_75t_R g5206 ( 
.A(n_2033),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_942),
.Y(n_5207)
);

CKINVDCx5p33_ASAP7_75t_R g5208 ( 
.A(n_325),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_4085),
.Y(n_5209)
);

CKINVDCx5p33_ASAP7_75t_R g5210 ( 
.A(n_2103),
.Y(n_5210)
);

CKINVDCx5p33_ASAP7_75t_R g5211 ( 
.A(n_970),
.Y(n_5211)
);

CKINVDCx5p33_ASAP7_75t_R g5212 ( 
.A(n_253),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_1757),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_479),
.Y(n_5214)
);

CKINVDCx5p33_ASAP7_75t_R g5215 ( 
.A(n_2262),
.Y(n_5215)
);

CKINVDCx5p33_ASAP7_75t_R g5216 ( 
.A(n_4062),
.Y(n_5216)
);

BUFx10_ASAP7_75t_L g5217 ( 
.A(n_3082),
.Y(n_5217)
);

BUFx2_ASAP7_75t_SL g5218 ( 
.A(n_640),
.Y(n_5218)
);

CKINVDCx5p33_ASAP7_75t_R g5219 ( 
.A(n_195),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_4055),
.Y(n_5220)
);

CKINVDCx5p33_ASAP7_75t_R g5221 ( 
.A(n_3679),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_72),
.Y(n_5222)
);

BUFx10_ASAP7_75t_L g5223 ( 
.A(n_4058),
.Y(n_5223)
);

CKINVDCx5p33_ASAP7_75t_R g5224 ( 
.A(n_958),
.Y(n_5224)
);

HB1xp67_ASAP7_75t_L g5225 ( 
.A(n_1596),
.Y(n_5225)
);

CKINVDCx5p33_ASAP7_75t_R g5226 ( 
.A(n_2403),
.Y(n_5226)
);

CKINVDCx5p33_ASAP7_75t_R g5227 ( 
.A(n_3569),
.Y(n_5227)
);

CKINVDCx5p33_ASAP7_75t_R g5228 ( 
.A(n_3416),
.Y(n_5228)
);

CKINVDCx5p33_ASAP7_75t_R g5229 ( 
.A(n_410),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_3505),
.Y(n_5230)
);

INVx1_ASAP7_75t_SL g5231 ( 
.A(n_2317),
.Y(n_5231)
);

INVx2_ASAP7_75t_SL g5232 ( 
.A(n_1221),
.Y(n_5232)
);

BUFx10_ASAP7_75t_L g5233 ( 
.A(n_2986),
.Y(n_5233)
);

CKINVDCx5p33_ASAP7_75t_R g5234 ( 
.A(n_261),
.Y(n_5234)
);

CKINVDCx5p33_ASAP7_75t_R g5235 ( 
.A(n_634),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_2223),
.Y(n_5236)
);

CKINVDCx5p33_ASAP7_75t_R g5237 ( 
.A(n_3205),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_1830),
.Y(n_5238)
);

CKINVDCx5p33_ASAP7_75t_R g5239 ( 
.A(n_819),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_2288),
.Y(n_5240)
);

CKINVDCx5p33_ASAP7_75t_R g5241 ( 
.A(n_2970),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_4028),
.Y(n_5242)
);

CKINVDCx5p33_ASAP7_75t_R g5243 ( 
.A(n_1010),
.Y(n_5243)
);

CKINVDCx5p33_ASAP7_75t_R g5244 ( 
.A(n_608),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_2332),
.Y(n_5245)
);

INVx2_ASAP7_75t_L g5246 ( 
.A(n_3321),
.Y(n_5246)
);

CKINVDCx5p33_ASAP7_75t_R g5247 ( 
.A(n_3790),
.Y(n_5247)
);

CKINVDCx14_ASAP7_75t_R g5248 ( 
.A(n_19),
.Y(n_5248)
);

CKINVDCx5p33_ASAP7_75t_R g5249 ( 
.A(n_721),
.Y(n_5249)
);

BUFx3_ASAP7_75t_L g5250 ( 
.A(n_1216),
.Y(n_5250)
);

CKINVDCx5p33_ASAP7_75t_R g5251 ( 
.A(n_2666),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_2488),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_4013),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_3572),
.Y(n_5254)
);

CKINVDCx5p33_ASAP7_75t_R g5255 ( 
.A(n_2849),
.Y(n_5255)
);

INVx1_ASAP7_75t_SL g5256 ( 
.A(n_4021),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_739),
.Y(n_5257)
);

CKINVDCx5p33_ASAP7_75t_R g5258 ( 
.A(n_2822),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_1337),
.Y(n_5259)
);

CKINVDCx20_ASAP7_75t_R g5260 ( 
.A(n_1667),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_480),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_2167),
.Y(n_5262)
);

CKINVDCx14_ASAP7_75t_R g5263 ( 
.A(n_1082),
.Y(n_5263)
);

INVx1_ASAP7_75t_SL g5264 ( 
.A(n_3593),
.Y(n_5264)
);

CKINVDCx5p33_ASAP7_75t_R g5265 ( 
.A(n_3957),
.Y(n_5265)
);

CKINVDCx5p33_ASAP7_75t_R g5266 ( 
.A(n_86),
.Y(n_5266)
);

INVx1_ASAP7_75t_SL g5267 ( 
.A(n_1729),
.Y(n_5267)
);

CKINVDCx5p33_ASAP7_75t_R g5268 ( 
.A(n_106),
.Y(n_5268)
);

CKINVDCx5p33_ASAP7_75t_R g5269 ( 
.A(n_2408),
.Y(n_5269)
);

CKINVDCx5p33_ASAP7_75t_R g5270 ( 
.A(n_258),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_2832),
.Y(n_5271)
);

BUFx10_ASAP7_75t_L g5272 ( 
.A(n_1839),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_2623),
.Y(n_5273)
);

CKINVDCx16_ASAP7_75t_R g5274 ( 
.A(n_3994),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_106),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_2725),
.Y(n_5276)
);

CKINVDCx5p33_ASAP7_75t_R g5277 ( 
.A(n_2534),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_2094),
.Y(n_5278)
);

CKINVDCx5p33_ASAP7_75t_R g5279 ( 
.A(n_2777),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_2880),
.Y(n_5280)
);

BUFx3_ASAP7_75t_L g5281 ( 
.A(n_3188),
.Y(n_5281)
);

CKINVDCx5p33_ASAP7_75t_R g5282 ( 
.A(n_1828),
.Y(n_5282)
);

CKINVDCx20_ASAP7_75t_R g5283 ( 
.A(n_1843),
.Y(n_5283)
);

CKINVDCx5p33_ASAP7_75t_R g5284 ( 
.A(n_3088),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_3910),
.Y(n_5285)
);

BUFx2_ASAP7_75t_L g5286 ( 
.A(n_3576),
.Y(n_5286)
);

CKINVDCx5p33_ASAP7_75t_R g5287 ( 
.A(n_1795),
.Y(n_5287)
);

CKINVDCx20_ASAP7_75t_R g5288 ( 
.A(n_3911),
.Y(n_5288)
);

BUFx2_ASAP7_75t_L g5289 ( 
.A(n_1542),
.Y(n_5289)
);

CKINVDCx5p33_ASAP7_75t_R g5290 ( 
.A(n_873),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_3948),
.Y(n_5291)
);

CKINVDCx5p33_ASAP7_75t_R g5292 ( 
.A(n_1874),
.Y(n_5292)
);

CKINVDCx20_ASAP7_75t_R g5293 ( 
.A(n_1553),
.Y(n_5293)
);

CKINVDCx5p33_ASAP7_75t_R g5294 ( 
.A(n_5),
.Y(n_5294)
);

CKINVDCx5p33_ASAP7_75t_R g5295 ( 
.A(n_1777),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_2476),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_1195),
.Y(n_5297)
);

CKINVDCx16_ASAP7_75t_R g5298 ( 
.A(n_1507),
.Y(n_5298)
);

BUFx3_ASAP7_75t_L g5299 ( 
.A(n_2861),
.Y(n_5299)
);

CKINVDCx5p33_ASAP7_75t_R g5300 ( 
.A(n_1822),
.Y(n_5300)
);

CKINVDCx5p33_ASAP7_75t_R g5301 ( 
.A(n_1364),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_4047),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_3057),
.Y(n_5303)
);

CKINVDCx5p33_ASAP7_75t_R g5304 ( 
.A(n_1333),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_3343),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_3976),
.Y(n_5306)
);

INVx1_ASAP7_75t_SL g5307 ( 
.A(n_2310),
.Y(n_5307)
);

CKINVDCx5p33_ASAP7_75t_R g5308 ( 
.A(n_2990),
.Y(n_5308)
);

CKINVDCx20_ASAP7_75t_R g5309 ( 
.A(n_2287),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_3129),
.Y(n_5310)
);

CKINVDCx5p33_ASAP7_75t_R g5311 ( 
.A(n_882),
.Y(n_5311)
);

BUFx2_ASAP7_75t_L g5312 ( 
.A(n_2804),
.Y(n_5312)
);

BUFx10_ASAP7_75t_L g5313 ( 
.A(n_2983),
.Y(n_5313)
);

CKINVDCx5p33_ASAP7_75t_R g5314 ( 
.A(n_767),
.Y(n_5314)
);

CKINVDCx5p33_ASAP7_75t_R g5315 ( 
.A(n_1056),
.Y(n_5315)
);

CKINVDCx5p33_ASAP7_75t_R g5316 ( 
.A(n_4086),
.Y(n_5316)
);

CKINVDCx5p33_ASAP7_75t_R g5317 ( 
.A(n_2346),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_919),
.Y(n_5318)
);

CKINVDCx5p33_ASAP7_75t_R g5319 ( 
.A(n_4051),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_2734),
.Y(n_5320)
);

CKINVDCx5p33_ASAP7_75t_R g5321 ( 
.A(n_3892),
.Y(n_5321)
);

CKINVDCx20_ASAP7_75t_R g5322 ( 
.A(n_3983),
.Y(n_5322)
);

CKINVDCx5p33_ASAP7_75t_R g5323 ( 
.A(n_3914),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_560),
.Y(n_5324)
);

CKINVDCx5p33_ASAP7_75t_R g5325 ( 
.A(n_254),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_3161),
.Y(n_5326)
);

CKINVDCx5p33_ASAP7_75t_R g5327 ( 
.A(n_955),
.Y(n_5327)
);

BUFx6f_ASAP7_75t_L g5328 ( 
.A(n_3536),
.Y(n_5328)
);

INVx1_ASAP7_75t_L g5329 ( 
.A(n_3699),
.Y(n_5329)
);

CKINVDCx5p33_ASAP7_75t_R g5330 ( 
.A(n_2012),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_1464),
.Y(n_5331)
);

CKINVDCx5p33_ASAP7_75t_R g5332 ( 
.A(n_2739),
.Y(n_5332)
);

BUFx10_ASAP7_75t_L g5333 ( 
.A(n_2194),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_1031),
.Y(n_5334)
);

CKINVDCx5p33_ASAP7_75t_R g5335 ( 
.A(n_2752),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_1691),
.Y(n_5336)
);

CKINVDCx20_ASAP7_75t_R g5337 ( 
.A(n_3405),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_1379),
.Y(n_5338)
);

CKINVDCx5p33_ASAP7_75t_R g5339 ( 
.A(n_4082),
.Y(n_5339)
);

CKINVDCx5p33_ASAP7_75t_R g5340 ( 
.A(n_1900),
.Y(n_5340)
);

CKINVDCx5p33_ASAP7_75t_R g5341 ( 
.A(n_2791),
.Y(n_5341)
);

CKINVDCx5p33_ASAP7_75t_R g5342 ( 
.A(n_2373),
.Y(n_5342)
);

CKINVDCx5p33_ASAP7_75t_R g5343 ( 
.A(n_2724),
.Y(n_5343)
);

CKINVDCx5p33_ASAP7_75t_R g5344 ( 
.A(n_3633),
.Y(n_5344)
);

BUFx6f_ASAP7_75t_L g5345 ( 
.A(n_3751),
.Y(n_5345)
);

CKINVDCx5p33_ASAP7_75t_R g5346 ( 
.A(n_71),
.Y(n_5346)
);

CKINVDCx5p33_ASAP7_75t_R g5347 ( 
.A(n_3935),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_4075),
.Y(n_5348)
);

CKINVDCx5p33_ASAP7_75t_R g5349 ( 
.A(n_218),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_1882),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_715),
.Y(n_5351)
);

CKINVDCx5p33_ASAP7_75t_R g5352 ( 
.A(n_1370),
.Y(n_5352)
);

CKINVDCx5p33_ASAP7_75t_R g5353 ( 
.A(n_1102),
.Y(n_5353)
);

CKINVDCx5p33_ASAP7_75t_R g5354 ( 
.A(n_1147),
.Y(n_5354)
);

INVx1_ASAP7_75t_SL g5355 ( 
.A(n_1728),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_3997),
.Y(n_5356)
);

CKINVDCx5p33_ASAP7_75t_R g5357 ( 
.A(n_1188),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_3999),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_2118),
.Y(n_5359)
);

CKINVDCx5p33_ASAP7_75t_R g5360 ( 
.A(n_1774),
.Y(n_5360)
);

CKINVDCx5p33_ASAP7_75t_R g5361 ( 
.A(n_3299),
.Y(n_5361)
);

CKINVDCx5p33_ASAP7_75t_R g5362 ( 
.A(n_2814),
.Y(n_5362)
);

BUFx6f_ASAP7_75t_L g5363 ( 
.A(n_1262),
.Y(n_5363)
);

CKINVDCx5p33_ASAP7_75t_R g5364 ( 
.A(n_4091),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_1221),
.Y(n_5365)
);

CKINVDCx5p33_ASAP7_75t_R g5366 ( 
.A(n_1629),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_1563),
.Y(n_5367)
);

BUFx3_ASAP7_75t_L g5368 ( 
.A(n_1940),
.Y(n_5368)
);

CKINVDCx5p33_ASAP7_75t_R g5369 ( 
.A(n_3436),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_309),
.Y(n_5370)
);

CKINVDCx5p33_ASAP7_75t_R g5371 ( 
.A(n_2533),
.Y(n_5371)
);

CKINVDCx5p33_ASAP7_75t_R g5372 ( 
.A(n_1299),
.Y(n_5372)
);

CKINVDCx5p33_ASAP7_75t_R g5373 ( 
.A(n_834),
.Y(n_5373)
);

CKINVDCx5p33_ASAP7_75t_R g5374 ( 
.A(n_3223),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_3995),
.Y(n_5375)
);

CKINVDCx5p33_ASAP7_75t_R g5376 ( 
.A(n_3215),
.Y(n_5376)
);

CKINVDCx5p33_ASAP7_75t_R g5377 ( 
.A(n_1474),
.Y(n_5377)
);

CKINVDCx5p33_ASAP7_75t_R g5378 ( 
.A(n_2151),
.Y(n_5378)
);

CKINVDCx5p33_ASAP7_75t_R g5379 ( 
.A(n_3530),
.Y(n_5379)
);

HB1xp67_ASAP7_75t_L g5380 ( 
.A(n_2650),
.Y(n_5380)
);

CKINVDCx5p33_ASAP7_75t_R g5381 ( 
.A(n_4012),
.Y(n_5381)
);

CKINVDCx5p33_ASAP7_75t_R g5382 ( 
.A(n_3108),
.Y(n_5382)
);

BUFx10_ASAP7_75t_L g5383 ( 
.A(n_3730),
.Y(n_5383)
);

CKINVDCx5p33_ASAP7_75t_R g5384 ( 
.A(n_731),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_1362),
.Y(n_5385)
);

INVx1_ASAP7_75t_SL g5386 ( 
.A(n_58),
.Y(n_5386)
);

CKINVDCx5p33_ASAP7_75t_R g5387 ( 
.A(n_4033),
.Y(n_5387)
);

INVxp67_ASAP7_75t_L g5388 ( 
.A(n_2604),
.Y(n_5388)
);

CKINVDCx20_ASAP7_75t_R g5389 ( 
.A(n_1560),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_2436),
.Y(n_5390)
);

CKINVDCx5p33_ASAP7_75t_R g5391 ( 
.A(n_1401),
.Y(n_5391)
);

CKINVDCx20_ASAP7_75t_R g5392 ( 
.A(n_3929),
.Y(n_5392)
);

CKINVDCx5p33_ASAP7_75t_R g5393 ( 
.A(n_1564),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_2859),
.Y(n_5394)
);

INVx2_ASAP7_75t_L g5395 ( 
.A(n_3712),
.Y(n_5395)
);

CKINVDCx5p33_ASAP7_75t_R g5396 ( 
.A(n_4086),
.Y(n_5396)
);

CKINVDCx5p33_ASAP7_75t_R g5397 ( 
.A(n_3582),
.Y(n_5397)
);

CKINVDCx5p33_ASAP7_75t_R g5398 ( 
.A(n_397),
.Y(n_5398)
);

CKINVDCx5p33_ASAP7_75t_R g5399 ( 
.A(n_1760),
.Y(n_5399)
);

CKINVDCx5p33_ASAP7_75t_R g5400 ( 
.A(n_2375),
.Y(n_5400)
);

CKINVDCx5p33_ASAP7_75t_R g5401 ( 
.A(n_2210),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_3318),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_499),
.Y(n_5403)
);

CKINVDCx5p33_ASAP7_75t_R g5404 ( 
.A(n_3240),
.Y(n_5404)
);

CKINVDCx5p33_ASAP7_75t_R g5405 ( 
.A(n_4041),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_259),
.Y(n_5406)
);

INVx1_ASAP7_75t_L g5407 ( 
.A(n_4004),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_3909),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_1372),
.Y(n_5409)
);

CKINVDCx5p33_ASAP7_75t_R g5410 ( 
.A(n_1999),
.Y(n_5410)
);

CKINVDCx5p33_ASAP7_75t_R g5411 ( 
.A(n_4045),
.Y(n_5411)
);

CKINVDCx5p33_ASAP7_75t_R g5412 ( 
.A(n_4110),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_3960),
.Y(n_5413)
);

CKINVDCx5p33_ASAP7_75t_R g5414 ( 
.A(n_2998),
.Y(n_5414)
);

CKINVDCx5p33_ASAP7_75t_R g5415 ( 
.A(n_953),
.Y(n_5415)
);

CKINVDCx5p33_ASAP7_75t_R g5416 ( 
.A(n_277),
.Y(n_5416)
);

CKINVDCx5p33_ASAP7_75t_R g5417 ( 
.A(n_3848),
.Y(n_5417)
);

CKINVDCx5p33_ASAP7_75t_R g5418 ( 
.A(n_3150),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_3953),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_701),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_45),
.Y(n_5421)
);

BUFx8_ASAP7_75t_SL g5422 ( 
.A(n_3978),
.Y(n_5422)
);

CKINVDCx5p33_ASAP7_75t_R g5423 ( 
.A(n_3209),
.Y(n_5423)
);

CKINVDCx5p33_ASAP7_75t_R g5424 ( 
.A(n_1338),
.Y(n_5424)
);

CKINVDCx5p33_ASAP7_75t_R g5425 ( 
.A(n_697),
.Y(n_5425)
);

CKINVDCx5p33_ASAP7_75t_R g5426 ( 
.A(n_1285),
.Y(n_5426)
);

INVx1_ASAP7_75t_SL g5427 ( 
.A(n_1613),
.Y(n_5427)
);

INVx2_ASAP7_75t_L g5428 ( 
.A(n_2267),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_2294),
.Y(n_5429)
);

CKINVDCx5p33_ASAP7_75t_R g5430 ( 
.A(n_3846),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_2986),
.Y(n_5431)
);

CKINVDCx5p33_ASAP7_75t_R g5432 ( 
.A(n_925),
.Y(n_5432)
);

CKINVDCx5p33_ASAP7_75t_R g5433 ( 
.A(n_3692),
.Y(n_5433)
);

CKINVDCx5p33_ASAP7_75t_R g5434 ( 
.A(n_820),
.Y(n_5434)
);

CKINVDCx5p33_ASAP7_75t_R g5435 ( 
.A(n_685),
.Y(n_5435)
);

CKINVDCx5p33_ASAP7_75t_R g5436 ( 
.A(n_3700),
.Y(n_5436)
);

CKINVDCx5p33_ASAP7_75t_R g5437 ( 
.A(n_2876),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_1081),
.Y(n_5438)
);

CKINVDCx5p33_ASAP7_75t_R g5439 ( 
.A(n_806),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_3005),
.Y(n_5440)
);

INVx2_ASAP7_75t_L g5441 ( 
.A(n_3748),
.Y(n_5441)
);

CKINVDCx5p33_ASAP7_75t_R g5442 ( 
.A(n_3898),
.Y(n_5442)
);

CKINVDCx5p33_ASAP7_75t_R g5443 ( 
.A(n_1490),
.Y(n_5443)
);

CKINVDCx20_ASAP7_75t_R g5444 ( 
.A(n_3920),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_1119),
.Y(n_5445)
);

CKINVDCx5p33_ASAP7_75t_R g5446 ( 
.A(n_3856),
.Y(n_5446)
);

CKINVDCx5p33_ASAP7_75t_R g5447 ( 
.A(n_835),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_3119),
.Y(n_5448)
);

CKINVDCx5p33_ASAP7_75t_R g5449 ( 
.A(n_2243),
.Y(n_5449)
);

CKINVDCx5p33_ASAP7_75t_R g5450 ( 
.A(n_4008),
.Y(n_5450)
);

CKINVDCx5p33_ASAP7_75t_R g5451 ( 
.A(n_398),
.Y(n_5451)
);

CKINVDCx5p33_ASAP7_75t_R g5452 ( 
.A(n_1805),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_3899),
.Y(n_5453)
);

CKINVDCx5p33_ASAP7_75t_R g5454 ( 
.A(n_2017),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_227),
.Y(n_5455)
);

CKINVDCx5p33_ASAP7_75t_R g5456 ( 
.A(n_2541),
.Y(n_5456)
);

BUFx3_ASAP7_75t_L g5457 ( 
.A(n_1736),
.Y(n_5457)
);

CKINVDCx5p33_ASAP7_75t_R g5458 ( 
.A(n_1942),
.Y(n_5458)
);

CKINVDCx5p33_ASAP7_75t_R g5459 ( 
.A(n_1625),
.Y(n_5459)
);

INVx2_ASAP7_75t_SL g5460 ( 
.A(n_2718),
.Y(n_5460)
);

CKINVDCx5p33_ASAP7_75t_R g5461 ( 
.A(n_1274),
.Y(n_5461)
);

INVx2_ASAP7_75t_SL g5462 ( 
.A(n_3544),
.Y(n_5462)
);

CKINVDCx5p33_ASAP7_75t_R g5463 ( 
.A(n_3938),
.Y(n_5463)
);

BUFx3_ASAP7_75t_L g5464 ( 
.A(n_913),
.Y(n_5464)
);

CKINVDCx5p33_ASAP7_75t_R g5465 ( 
.A(n_3190),
.Y(n_5465)
);

CKINVDCx5p33_ASAP7_75t_R g5466 ( 
.A(n_4084),
.Y(n_5466)
);

CKINVDCx16_ASAP7_75t_R g5467 ( 
.A(n_1675),
.Y(n_5467)
);

BUFx10_ASAP7_75t_L g5468 ( 
.A(n_3688),
.Y(n_5468)
);

CKINVDCx5p33_ASAP7_75t_R g5469 ( 
.A(n_3982),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_3700),
.Y(n_5470)
);

CKINVDCx5p33_ASAP7_75t_R g5471 ( 
.A(n_4038),
.Y(n_5471)
);

BUFx10_ASAP7_75t_L g5472 ( 
.A(n_239),
.Y(n_5472)
);

CKINVDCx5p33_ASAP7_75t_R g5473 ( 
.A(n_4025),
.Y(n_5473)
);

CKINVDCx5p33_ASAP7_75t_R g5474 ( 
.A(n_394),
.Y(n_5474)
);

CKINVDCx5p33_ASAP7_75t_R g5475 ( 
.A(n_4015),
.Y(n_5475)
);

CKINVDCx5p33_ASAP7_75t_R g5476 ( 
.A(n_240),
.Y(n_5476)
);

CKINVDCx5p33_ASAP7_75t_R g5477 ( 
.A(n_1738),
.Y(n_5477)
);

INVx2_ASAP7_75t_L g5478 ( 
.A(n_1120),
.Y(n_5478)
);

CKINVDCx5p33_ASAP7_75t_R g5479 ( 
.A(n_3943),
.Y(n_5479)
);

CKINVDCx5p33_ASAP7_75t_R g5480 ( 
.A(n_3640),
.Y(n_5480)
);

INVx2_ASAP7_75t_SL g5481 ( 
.A(n_2903),
.Y(n_5481)
);

CKINVDCx20_ASAP7_75t_R g5482 ( 
.A(n_4001),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_3901),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_3984),
.Y(n_5484)
);

BUFx2_ASAP7_75t_SL g5485 ( 
.A(n_741),
.Y(n_5485)
);

CKINVDCx5p33_ASAP7_75t_R g5486 ( 
.A(n_1382),
.Y(n_5486)
);

CKINVDCx5p33_ASAP7_75t_R g5487 ( 
.A(n_1314),
.Y(n_5487)
);

CKINVDCx5p33_ASAP7_75t_R g5488 ( 
.A(n_3906),
.Y(n_5488)
);

CKINVDCx5p33_ASAP7_75t_R g5489 ( 
.A(n_1996),
.Y(n_5489)
);

INVxp67_ASAP7_75t_L g5490 ( 
.A(n_1782),
.Y(n_5490)
);

CKINVDCx5p33_ASAP7_75t_R g5491 ( 
.A(n_3384),
.Y(n_5491)
);

INVx1_ASAP7_75t_L g5492 ( 
.A(n_1338),
.Y(n_5492)
);

CKINVDCx5p33_ASAP7_75t_R g5493 ( 
.A(n_3959),
.Y(n_5493)
);

CKINVDCx20_ASAP7_75t_R g5494 ( 
.A(n_4016),
.Y(n_5494)
);

CKINVDCx5p33_ASAP7_75t_R g5495 ( 
.A(n_2859),
.Y(n_5495)
);

CKINVDCx20_ASAP7_75t_R g5496 ( 
.A(n_395),
.Y(n_5496)
);

BUFx6f_ASAP7_75t_L g5497 ( 
.A(n_3574),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_98),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_3993),
.Y(n_5499)
);

CKINVDCx20_ASAP7_75t_R g5500 ( 
.A(n_2750),
.Y(n_5500)
);

CKINVDCx20_ASAP7_75t_R g5501 ( 
.A(n_4089),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_3136),
.Y(n_5502)
);

INVx1_ASAP7_75t_SL g5503 ( 
.A(n_1177),
.Y(n_5503)
);

CKINVDCx20_ASAP7_75t_R g5504 ( 
.A(n_582),
.Y(n_5504)
);

CKINVDCx5p33_ASAP7_75t_R g5505 ( 
.A(n_632),
.Y(n_5505)
);

INVx2_ASAP7_75t_L g5506 ( 
.A(n_1705),
.Y(n_5506)
);

CKINVDCx5p33_ASAP7_75t_R g5507 ( 
.A(n_2549),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_266),
.Y(n_5508)
);

CKINVDCx5p33_ASAP7_75t_R g5509 ( 
.A(n_1668),
.Y(n_5509)
);

CKINVDCx5p33_ASAP7_75t_R g5510 ( 
.A(n_2023),
.Y(n_5510)
);

CKINVDCx5p33_ASAP7_75t_R g5511 ( 
.A(n_3552),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_3937),
.Y(n_5512)
);

CKINVDCx5p33_ASAP7_75t_R g5513 ( 
.A(n_4079),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_327),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_3449),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_3847),
.Y(n_5516)
);

INVx2_ASAP7_75t_L g5517 ( 
.A(n_3927),
.Y(n_5517)
);

CKINVDCx16_ASAP7_75t_R g5518 ( 
.A(n_1863),
.Y(n_5518)
);

CKINVDCx5p33_ASAP7_75t_R g5519 ( 
.A(n_1288),
.Y(n_5519)
);

CKINVDCx5p33_ASAP7_75t_R g5520 ( 
.A(n_3557),
.Y(n_5520)
);

CKINVDCx5p33_ASAP7_75t_R g5521 ( 
.A(n_2537),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_3975),
.Y(n_5522)
);

INVx2_ASAP7_75t_L g5523 ( 
.A(n_3577),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_3103),
.Y(n_5524)
);

CKINVDCx5p33_ASAP7_75t_R g5525 ( 
.A(n_812),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_2448),
.Y(n_5526)
);

CKINVDCx20_ASAP7_75t_R g5527 ( 
.A(n_2232),
.Y(n_5527)
);

BUFx6f_ASAP7_75t_L g5528 ( 
.A(n_1860),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_4048),
.Y(n_5529)
);

CKINVDCx5p33_ASAP7_75t_R g5530 ( 
.A(n_3676),
.Y(n_5530)
);

CKINVDCx20_ASAP7_75t_R g5531 ( 
.A(n_3918),
.Y(n_5531)
);

CKINVDCx5p33_ASAP7_75t_R g5532 ( 
.A(n_1452),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_3189),
.Y(n_5533)
);

CKINVDCx5p33_ASAP7_75t_R g5534 ( 
.A(n_202),
.Y(n_5534)
);

BUFx5_ASAP7_75t_L g5535 ( 
.A(n_4022),
.Y(n_5535)
);

BUFx3_ASAP7_75t_L g5536 ( 
.A(n_3309),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_988),
.Y(n_5537)
);

CKINVDCx5p33_ASAP7_75t_R g5538 ( 
.A(n_2685),
.Y(n_5538)
);

CKINVDCx5p33_ASAP7_75t_R g5539 ( 
.A(n_2399),
.Y(n_5539)
);

CKINVDCx5p33_ASAP7_75t_R g5540 ( 
.A(n_2187),
.Y(n_5540)
);

CKINVDCx5p33_ASAP7_75t_R g5541 ( 
.A(n_3441),
.Y(n_5541)
);

CKINVDCx5p33_ASAP7_75t_R g5542 ( 
.A(n_3974),
.Y(n_5542)
);

CKINVDCx5p33_ASAP7_75t_R g5543 ( 
.A(n_3288),
.Y(n_5543)
);

CKINVDCx5p33_ASAP7_75t_R g5544 ( 
.A(n_3055),
.Y(n_5544)
);

INVx2_ASAP7_75t_L g5545 ( 
.A(n_3407),
.Y(n_5545)
);

CKINVDCx5p33_ASAP7_75t_R g5546 ( 
.A(n_1999),
.Y(n_5546)
);

INVx2_ASAP7_75t_SL g5547 ( 
.A(n_3949),
.Y(n_5547)
);

CKINVDCx20_ASAP7_75t_R g5548 ( 
.A(n_1370),
.Y(n_5548)
);

CKINVDCx5p33_ASAP7_75t_R g5549 ( 
.A(n_1025),
.Y(n_5549)
);

CKINVDCx20_ASAP7_75t_R g5550 ( 
.A(n_264),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_4993),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_4993),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4976),
.Y(n_5553)
);

CKINVDCx16_ASAP7_75t_R g5554 ( 
.A(n_5248),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_4194),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_4194),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4194),
.Y(n_5557)
);

CKINVDCx5p33_ASAP7_75t_R g5558 ( 
.A(n_4152),
.Y(n_5558)
);

CKINVDCx5p33_ASAP7_75t_R g5559 ( 
.A(n_4366),
.Y(n_5559)
);

BUFx6f_ASAP7_75t_L g5560 ( 
.A(n_4277),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_4194),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_4194),
.Y(n_5562)
);

INVx2_ASAP7_75t_L g5563 ( 
.A(n_4214),
.Y(n_5563)
);

CKINVDCx5p33_ASAP7_75t_R g5564 ( 
.A(n_4577),
.Y(n_5564)
);

NOR2xp67_ASAP7_75t_L g5565 ( 
.A(n_4514),
.B(n_0),
.Y(n_5565)
);

CKINVDCx20_ASAP7_75t_R g5566 ( 
.A(n_4233),
.Y(n_5566)
);

BUFx3_ASAP7_75t_L g5567 ( 
.A(n_4158),
.Y(n_5567)
);

CKINVDCx5p33_ASAP7_75t_R g5568 ( 
.A(n_4710),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_4214),
.Y(n_5569)
);

BUFx6f_ASAP7_75t_L g5570 ( 
.A(n_4277),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_4214),
.Y(n_5571)
);

CKINVDCx5p33_ASAP7_75t_R g5572 ( 
.A(n_5422),
.Y(n_5572)
);

BUFx2_ASAP7_75t_L g5573 ( 
.A(n_4406),
.Y(n_5573)
);

CKINVDCx5p33_ASAP7_75t_R g5574 ( 
.A(n_4186),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_4214),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_4214),
.Y(n_5576)
);

INVx2_ASAP7_75t_L g5577 ( 
.A(n_4443),
.Y(n_5577)
);

CKINVDCx5p33_ASAP7_75t_R g5578 ( 
.A(n_4204),
.Y(n_5578)
);

INVx2_ASAP7_75t_L g5579 ( 
.A(n_4443),
.Y(n_5579)
);

INVx2_ASAP7_75t_L g5580 ( 
.A(n_4443),
.Y(n_5580)
);

CKINVDCx5p33_ASAP7_75t_R g5581 ( 
.A(n_4206),
.Y(n_5581)
);

INVx2_ASAP7_75t_SL g5582 ( 
.A(n_4734),
.Y(n_5582)
);

INVx2_ASAP7_75t_L g5583 ( 
.A(n_4443),
.Y(n_5583)
);

CKINVDCx5p33_ASAP7_75t_R g5584 ( 
.A(n_4227),
.Y(n_5584)
);

HB1xp67_ASAP7_75t_L g5585 ( 
.A(n_5101),
.Y(n_5585)
);

INVx2_ASAP7_75t_L g5586 ( 
.A(n_4443),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_4569),
.Y(n_5587)
);

BUFx10_ASAP7_75t_L g5588 ( 
.A(n_4765),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_4569),
.Y(n_5589)
);

BUFx2_ASAP7_75t_SL g5590 ( 
.A(n_4569),
.Y(n_5590)
);

CKINVDCx5p33_ASAP7_75t_R g5591 ( 
.A(n_4247),
.Y(n_5591)
);

BUFx5_ASAP7_75t_L g5592 ( 
.A(n_4131),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_4569),
.Y(n_5593)
);

CKINVDCx5p33_ASAP7_75t_R g5594 ( 
.A(n_4312),
.Y(n_5594)
);

CKINVDCx16_ASAP7_75t_R g5595 ( 
.A(n_4504),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_4569),
.Y(n_5596)
);

CKINVDCx5p33_ASAP7_75t_R g5597 ( 
.A(n_4743),
.Y(n_5597)
);

CKINVDCx5p33_ASAP7_75t_R g5598 ( 
.A(n_4781),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_4752),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_4752),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_4752),
.Y(n_5601)
);

CKINVDCx5p33_ASAP7_75t_R g5602 ( 
.A(n_4822),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_4752),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_4752),
.Y(n_5604)
);

CKINVDCx20_ASAP7_75t_R g5605 ( 
.A(n_4834),
.Y(n_5605)
);

BUFx3_ASAP7_75t_L g5606 ( 
.A(n_4164),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_5044),
.Y(n_5607)
);

CKINVDCx5p33_ASAP7_75t_R g5608 ( 
.A(n_4849),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_5044),
.Y(n_5609)
);

CKINVDCx5p33_ASAP7_75t_R g5610 ( 
.A(n_4876),
.Y(n_5610)
);

CKINVDCx5p33_ASAP7_75t_R g5611 ( 
.A(n_4977),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5044),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5044),
.Y(n_5613)
);

INVx2_ASAP7_75t_L g5614 ( 
.A(n_5044),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5535),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5535),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5535),
.Y(n_5617)
);

CKINVDCx20_ASAP7_75t_R g5618 ( 
.A(n_4969),
.Y(n_5618)
);

CKINVDCx5p33_ASAP7_75t_R g5619 ( 
.A(n_5014),
.Y(n_5619)
);

CKINVDCx5p33_ASAP7_75t_R g5620 ( 
.A(n_5073),
.Y(n_5620)
);

CKINVDCx5p33_ASAP7_75t_R g5621 ( 
.A(n_5075),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5535),
.Y(n_5622)
);

BUFx3_ASAP7_75t_L g5623 ( 
.A(n_4166),
.Y(n_5623)
);

CKINVDCx5p33_ASAP7_75t_R g5624 ( 
.A(n_5198),
.Y(n_5624)
);

CKINVDCx5p33_ASAP7_75t_R g5625 ( 
.A(n_5274),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5535),
.Y(n_5626)
);

BUFx10_ASAP7_75t_L g5627 ( 
.A(n_4828),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_4301),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_4468),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_4530),
.Y(n_5630)
);

INVx2_ASAP7_75t_L g5631 ( 
.A(n_4587),
.Y(n_5631)
);

CKINVDCx20_ASAP7_75t_R g5632 ( 
.A(n_4997),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_4643),
.Y(n_5633)
);

INVx2_ASAP7_75t_SL g5634 ( 
.A(n_4734),
.Y(n_5634)
);

INVx1_ASAP7_75t_SL g5635 ( 
.A(n_5016),
.Y(n_5635)
);

CKINVDCx5p33_ASAP7_75t_R g5636 ( 
.A(n_5298),
.Y(n_5636)
);

CKINVDCx5p33_ASAP7_75t_R g5637 ( 
.A(n_5467),
.Y(n_5637)
);

INVx2_ASAP7_75t_L g5638 ( 
.A(n_4811),
.Y(n_5638)
);

CKINVDCx5p33_ASAP7_75t_R g5639 ( 
.A(n_5518),
.Y(n_5639)
);

CKINVDCx5p33_ASAP7_75t_R g5640 ( 
.A(n_5111),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_4951),
.Y(n_5641)
);

OR2x2_ASAP7_75t_L g5642 ( 
.A(n_4127),
.B(n_0),
.Y(n_5642)
);

INVxp33_ASAP7_75t_L g5643 ( 
.A(n_4919),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5059),
.Y(n_5644)
);

CKINVDCx5p33_ASAP7_75t_R g5645 ( 
.A(n_5188),
.Y(n_5645)
);

CKINVDCx20_ASAP7_75t_R g5646 ( 
.A(n_5263),
.Y(n_5646)
);

CKINVDCx5p33_ASAP7_75t_R g5647 ( 
.A(n_5549),
.Y(n_5647)
);

CKINVDCx5p33_ASAP7_75t_R g5648 ( 
.A(n_4123),
.Y(n_5648)
);

BUFx3_ASAP7_75t_L g5649 ( 
.A(n_4243),
.Y(n_5649)
);

BUFx6f_ASAP7_75t_L g5650 ( 
.A(n_4277),
.Y(n_5650)
);

CKINVDCx5p33_ASAP7_75t_R g5651 ( 
.A(n_4124),
.Y(n_5651)
);

CKINVDCx16_ASAP7_75t_R g5652 ( 
.A(n_4205),
.Y(n_5652)
);

CKINVDCx5p33_ASAP7_75t_R g5653 ( 
.A(n_5534),
.Y(n_5653)
);

CKINVDCx5p33_ASAP7_75t_R g5654 ( 
.A(n_5538),
.Y(n_5654)
);

CKINVDCx5p33_ASAP7_75t_R g5655 ( 
.A(n_5539),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5222),
.Y(n_5656)
);

CKINVDCx5p33_ASAP7_75t_R g5657 ( 
.A(n_5540),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5275),
.Y(n_5658)
);

CKINVDCx5p33_ASAP7_75t_R g5659 ( 
.A(n_5541),
.Y(n_5659)
);

CKINVDCx5p33_ASAP7_75t_R g5660 ( 
.A(n_5542),
.Y(n_5660)
);

CKINVDCx5p33_ASAP7_75t_R g5661 ( 
.A(n_5543),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5421),
.Y(n_5662)
);

CKINVDCx20_ASAP7_75t_R g5663 ( 
.A(n_5548),
.Y(n_5663)
);

BUFx2_ASAP7_75t_L g5664 ( 
.A(n_4183),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5498),
.Y(n_5665)
);

BUFx6f_ASAP7_75t_L g5666 ( 
.A(n_4629),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_4517),
.Y(n_5667)
);

CKINVDCx5p33_ASAP7_75t_R g5668 ( 
.A(n_4125),
.Y(n_5668)
);

CKINVDCx5p33_ASAP7_75t_R g5669 ( 
.A(n_4130),
.Y(n_5669)
);

CKINVDCx20_ASAP7_75t_R g5670 ( 
.A(n_5527),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_4126),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_4128),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_4132),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_4140),
.Y(n_5674)
);

CKINVDCx5p33_ASAP7_75t_R g5675 ( 
.A(n_5532),
.Y(n_5675)
);

CKINVDCx20_ASAP7_75t_R g5676 ( 
.A(n_5531),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_4141),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_4144),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_4148),
.Y(n_5679)
);

CKINVDCx5p33_ASAP7_75t_R g5680 ( 
.A(n_5544),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_4161),
.Y(n_5681)
);

INVx1_ASAP7_75t_L g5682 ( 
.A(n_4165),
.Y(n_5682)
);

CKINVDCx5p33_ASAP7_75t_R g5683 ( 
.A(n_4133),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_4168),
.Y(n_5684)
);

CKINVDCx5p33_ASAP7_75t_R g5685 ( 
.A(n_4134),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_4171),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_4175),
.Y(n_5687)
);

CKINVDCx5p33_ASAP7_75t_R g5688 ( 
.A(n_5525),
.Y(n_5688)
);

CKINVDCx5p33_ASAP7_75t_R g5689 ( 
.A(n_5530),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_4176),
.Y(n_5690)
);

HB1xp67_ASAP7_75t_L g5691 ( 
.A(n_5038),
.Y(n_5691)
);

CKINVDCx5p33_ASAP7_75t_R g5692 ( 
.A(n_5546),
.Y(n_5692)
);

CKINVDCx5p33_ASAP7_75t_R g5693 ( 
.A(n_4135),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_4177),
.Y(n_5694)
);

CKINVDCx20_ASAP7_75t_R g5695 ( 
.A(n_5550),
.Y(n_5695)
);

INVx1_ASAP7_75t_SL g5696 ( 
.A(n_4129),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_4181),
.Y(n_5697)
);

CKINVDCx5p33_ASAP7_75t_R g5698 ( 
.A(n_4137),
.Y(n_5698)
);

CKINVDCx5p33_ASAP7_75t_R g5699 ( 
.A(n_4138),
.Y(n_5699)
);

BUFx10_ASAP7_75t_L g5700 ( 
.A(n_5225),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_4187),
.Y(n_5701)
);

BUFx10_ASAP7_75t_L g5702 ( 
.A(n_5380),
.Y(n_5702)
);

INVx1_ASAP7_75t_SL g5703 ( 
.A(n_4173),
.Y(n_5703)
);

BUFx2_ASAP7_75t_SL g5704 ( 
.A(n_5528),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_4191),
.Y(n_5705)
);

CKINVDCx16_ASAP7_75t_R g5706 ( 
.A(n_4205),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_4629),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_4193),
.Y(n_5708)
);

BUFx5_ASAP7_75t_L g5709 ( 
.A(n_4195),
.Y(n_5709)
);

CKINVDCx5p33_ASAP7_75t_R g5710 ( 
.A(n_4139),
.Y(n_5710)
);

NOR2xp67_ASAP7_75t_L g5711 ( 
.A(n_4276),
.B(n_0),
.Y(n_5711)
);

CKINVDCx5p33_ASAP7_75t_R g5712 ( 
.A(n_4142),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_4196),
.Y(n_5713)
);

BUFx10_ASAP7_75t_L g5714 ( 
.A(n_4162),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_4198),
.Y(n_5715)
);

CKINVDCx5p33_ASAP7_75t_R g5716 ( 
.A(n_4143),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_4208),
.Y(n_5717)
);

CKINVDCx20_ASAP7_75t_R g5718 ( 
.A(n_4221),
.Y(n_5718)
);

INVx2_ASAP7_75t_L g5719 ( 
.A(n_4629),
.Y(n_5719)
);

CKINVDCx16_ASAP7_75t_R g5720 ( 
.A(n_4241),
.Y(n_5720)
);

CKINVDCx5p33_ASAP7_75t_R g5721 ( 
.A(n_5519),
.Y(n_5721)
);

CKINVDCx5p33_ASAP7_75t_R g5722 ( 
.A(n_5520),
.Y(n_5722)
);

INVx1_ASAP7_75t_L g5723 ( 
.A(n_4209),
.Y(n_5723)
);

CKINVDCx5p33_ASAP7_75t_R g5724 ( 
.A(n_5521),
.Y(n_5724)
);

CKINVDCx5p33_ASAP7_75t_R g5725 ( 
.A(n_4145),
.Y(n_5725)
);

CKINVDCx5p33_ASAP7_75t_R g5726 ( 
.A(n_4146),
.Y(n_5726)
);

NOR2xp67_ASAP7_75t_L g5727 ( 
.A(n_4816),
.B(n_1),
.Y(n_5727)
);

CKINVDCx5p33_ASAP7_75t_R g5728 ( 
.A(n_4147),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_4211),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_4213),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_4655),
.Y(n_5731)
);

INVxp67_ASAP7_75t_SL g5732 ( 
.A(n_4655),
.Y(n_5732)
);

CKINVDCx20_ASAP7_75t_R g5733 ( 
.A(n_4242),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_4219),
.Y(n_5734)
);

CKINVDCx14_ASAP7_75t_R g5735 ( 
.A(n_4241),
.Y(n_5735)
);

CKINVDCx5p33_ASAP7_75t_R g5736 ( 
.A(n_4149),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_4220),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_4229),
.Y(n_5738)
);

CKINVDCx5p33_ASAP7_75t_R g5739 ( 
.A(n_4150),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_4232),
.Y(n_5740)
);

CKINVDCx5p33_ASAP7_75t_R g5741 ( 
.A(n_4151),
.Y(n_5741)
);

INVxp67_ASAP7_75t_SL g5742 ( 
.A(n_4655),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_4235),
.Y(n_5743)
);

CKINVDCx5p33_ASAP7_75t_R g5744 ( 
.A(n_4153),
.Y(n_5744)
);

CKINVDCx14_ASAP7_75t_R g5745 ( 
.A(n_4309),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_4237),
.Y(n_5746)
);

CKINVDCx5p33_ASAP7_75t_R g5747 ( 
.A(n_4154),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_4238),
.Y(n_5748)
);

CKINVDCx5p33_ASAP7_75t_R g5749 ( 
.A(n_4155),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_4239),
.Y(n_5750)
);

CKINVDCx5p33_ASAP7_75t_R g5751 ( 
.A(n_4156),
.Y(n_5751)
);

INVx1_ASAP7_75t_SL g5752 ( 
.A(n_4266),
.Y(n_5752)
);

INVx2_ASAP7_75t_L g5753 ( 
.A(n_4708),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_4244),
.Y(n_5754)
);

CKINVDCx14_ASAP7_75t_R g5755 ( 
.A(n_4309),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_4246),
.Y(n_5756)
);

CKINVDCx5p33_ASAP7_75t_R g5757 ( 
.A(n_4157),
.Y(n_5757)
);

CKINVDCx5p33_ASAP7_75t_R g5758 ( 
.A(n_4159),
.Y(n_5758)
);

CKINVDCx5p33_ASAP7_75t_R g5759 ( 
.A(n_4160),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_4253),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_4260),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_4267),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_4270),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_4272),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_4273),
.Y(n_5765)
);

CKINVDCx5p33_ASAP7_75t_R g5766 ( 
.A(n_4163),
.Y(n_5766)
);

CKINVDCx5p33_ASAP7_75t_R g5767 ( 
.A(n_4167),
.Y(n_5767)
);

NOR2xp33_ASAP7_75t_L g5768 ( 
.A(n_4304),
.B(n_1),
.Y(n_5768)
);

INVx1_ASAP7_75t_L g5769 ( 
.A(n_4274),
.Y(n_5769)
);

CKINVDCx5p33_ASAP7_75t_R g5770 ( 
.A(n_4169),
.Y(n_5770)
);

CKINVDCx5p33_ASAP7_75t_R g5771 ( 
.A(n_4170),
.Y(n_5771)
);

INVx1_ASAP7_75t_SL g5772 ( 
.A(n_4290),
.Y(n_5772)
);

CKINVDCx5p33_ASAP7_75t_R g5773 ( 
.A(n_4174),
.Y(n_5773)
);

CKINVDCx16_ASAP7_75t_R g5774 ( 
.A(n_4669),
.Y(n_5774)
);

CKINVDCx5p33_ASAP7_75t_R g5775 ( 
.A(n_4179),
.Y(n_5775)
);

CKINVDCx5p33_ASAP7_75t_R g5776 ( 
.A(n_4180),
.Y(n_5776)
);

CKINVDCx5p33_ASAP7_75t_R g5777 ( 
.A(n_4182),
.Y(n_5777)
);

CKINVDCx5p33_ASAP7_75t_R g5778 ( 
.A(n_4184),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_4708),
.Y(n_5779)
);

CKINVDCx5p33_ASAP7_75t_R g5780 ( 
.A(n_4185),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_4280),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_4282),
.Y(n_5782)
);

CKINVDCx5p33_ASAP7_75t_R g5783 ( 
.A(n_4188),
.Y(n_5783)
);

CKINVDCx5p33_ASAP7_75t_R g5784 ( 
.A(n_4189),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_4283),
.Y(n_5785)
);

CKINVDCx5p33_ASAP7_75t_R g5786 ( 
.A(n_4190),
.Y(n_5786)
);

BUFx3_ASAP7_75t_L g5787 ( 
.A(n_4297),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_4286),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_4293),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_4313),
.Y(n_5790)
);

CKINVDCx5p33_ASAP7_75t_R g5791 ( 
.A(n_4192),
.Y(n_5791)
);

BUFx6f_ASAP7_75t_L g5792 ( 
.A(n_5528),
.Y(n_5792)
);

CKINVDCx5p33_ASAP7_75t_R g5793 ( 
.A(n_4197),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_4319),
.Y(n_5794)
);

BUFx6f_ASAP7_75t_L g5795 ( 
.A(n_5528),
.Y(n_5795)
);

CKINVDCx5p33_ASAP7_75t_R g5796 ( 
.A(n_4199),
.Y(n_5796)
);

CKINVDCx5p33_ASAP7_75t_R g5797 ( 
.A(n_4200),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_4321),
.Y(n_5798)
);

INVx2_ASAP7_75t_SL g5799 ( 
.A(n_4669),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_4322),
.Y(n_5800)
);

INVx1_ASAP7_75t_L g5801 ( 
.A(n_4323),
.Y(n_5801)
);

BUFx3_ASAP7_75t_L g5802 ( 
.A(n_5536),
.Y(n_5802)
);

BUFx6f_ASAP7_75t_L g5803 ( 
.A(n_4708),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_4325),
.Y(n_5804)
);

INVx1_ASAP7_75t_SL g5805 ( 
.A(n_4292),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_4327),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_4329),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_4330),
.Y(n_5808)
);

CKINVDCx5p33_ASAP7_75t_R g5809 ( 
.A(n_5513),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_4331),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_4339),
.Y(n_5811)
);

CKINVDCx5p33_ASAP7_75t_R g5812 ( 
.A(n_4202),
.Y(n_5812)
);

CKINVDCx5p33_ASAP7_75t_R g5813 ( 
.A(n_4207),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_4344),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_4347),
.Y(n_5815)
);

CKINVDCx5p33_ASAP7_75t_R g5816 ( 
.A(n_4210),
.Y(n_5816)
);

CKINVDCx5p33_ASAP7_75t_R g5817 ( 
.A(n_4215),
.Y(n_5817)
);

CKINVDCx5p33_ASAP7_75t_R g5818 ( 
.A(n_4216),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_4350),
.Y(n_5819)
);

INVx2_ASAP7_75t_L g5820 ( 
.A(n_4756),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_4356),
.Y(n_5821)
);

BUFx6f_ASAP7_75t_L g5822 ( 
.A(n_4756),
.Y(n_5822)
);

CKINVDCx5p33_ASAP7_75t_R g5823 ( 
.A(n_4217),
.Y(n_5823)
);

BUFx6f_ASAP7_75t_L g5824 ( 
.A(n_4756),
.Y(n_5824)
);

CKINVDCx5p33_ASAP7_75t_R g5825 ( 
.A(n_4218),
.Y(n_5825)
);

BUFx10_ASAP7_75t_L g5826 ( 
.A(n_4245),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_4359),
.Y(n_5827)
);

CKINVDCx5p33_ASAP7_75t_R g5828 ( 
.A(n_4222),
.Y(n_5828)
);

OR2x2_ASAP7_75t_L g5829 ( 
.A(n_4360),
.B(n_1),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_4361),
.Y(n_5830)
);

CKINVDCx5p33_ASAP7_75t_R g5831 ( 
.A(n_4223),
.Y(n_5831)
);

CKINVDCx20_ASAP7_75t_R g5832 ( 
.A(n_4314),
.Y(n_5832)
);

CKINVDCx5p33_ASAP7_75t_R g5833 ( 
.A(n_4225),
.Y(n_5833)
);

CKINVDCx5p33_ASAP7_75t_R g5834 ( 
.A(n_4226),
.Y(n_5834)
);

CKINVDCx5p33_ASAP7_75t_R g5835 ( 
.A(n_4228),
.Y(n_5835)
);

CKINVDCx16_ASAP7_75t_R g5836 ( 
.A(n_4694),
.Y(n_5836)
);

INVxp67_ASAP7_75t_SL g5837 ( 
.A(n_4944),
.Y(n_5837)
);

INVx2_ASAP7_75t_SL g5838 ( 
.A(n_4694),
.Y(n_5838)
);

CKINVDCx5p33_ASAP7_75t_R g5839 ( 
.A(n_4230),
.Y(n_5839)
);

XNOR2x1_ASAP7_75t_L g5840 ( 
.A(n_4343),
.B(n_2),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_4363),
.Y(n_5841)
);

CKINVDCx5p33_ASAP7_75t_R g5842 ( 
.A(n_4231),
.Y(n_5842)
);

CKINVDCx5p33_ASAP7_75t_R g5843 ( 
.A(n_4234),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_4370),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_4372),
.Y(n_5845)
);

CKINVDCx5p33_ASAP7_75t_R g5846 ( 
.A(n_4236),
.Y(n_5846)
);

CKINVDCx5p33_ASAP7_75t_R g5847 ( 
.A(n_4240),
.Y(n_5847)
);

INVxp67_ASAP7_75t_SL g5848 ( 
.A(n_4944),
.Y(n_5848)
);

BUFx10_ASAP7_75t_L g5849 ( 
.A(n_4349),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_4374),
.Y(n_5850)
);

BUFx6f_ASAP7_75t_L g5851 ( 
.A(n_4944),
.Y(n_5851)
);

CKINVDCx5p33_ASAP7_75t_R g5852 ( 
.A(n_4248),
.Y(n_5852)
);

BUFx3_ASAP7_75t_L g5853 ( 
.A(n_4317),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_4379),
.Y(n_5854)
);

INVx2_ASAP7_75t_L g5855 ( 
.A(n_4971),
.Y(n_5855)
);

CKINVDCx5p33_ASAP7_75t_R g5856 ( 
.A(n_4249),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_4383),
.Y(n_5857)
);

CKINVDCx5p33_ASAP7_75t_R g5858 ( 
.A(n_4250),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_4398),
.Y(n_5859)
);

CKINVDCx20_ASAP7_75t_R g5860 ( 
.A(n_4328),
.Y(n_5860)
);

INVx1_ASAP7_75t_L g5861 ( 
.A(n_4399),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_4407),
.Y(n_5862)
);

CKINVDCx5p33_ASAP7_75t_R g5863 ( 
.A(n_4251),
.Y(n_5863)
);

CKINVDCx5p33_ASAP7_75t_R g5864 ( 
.A(n_4252),
.Y(n_5864)
);

CKINVDCx5p33_ASAP7_75t_R g5865 ( 
.A(n_4254),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_4408),
.Y(n_5866)
);

CKINVDCx5p33_ASAP7_75t_R g5867 ( 
.A(n_4255),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_4413),
.Y(n_5868)
);

CKINVDCx16_ASAP7_75t_R g5869 ( 
.A(n_4696),
.Y(n_5869)
);

CKINVDCx5p33_ASAP7_75t_R g5870 ( 
.A(n_4256),
.Y(n_5870)
);

CKINVDCx20_ASAP7_75t_R g5871 ( 
.A(n_4335),
.Y(n_5871)
);

CKINVDCx5p33_ASAP7_75t_R g5872 ( 
.A(n_4257),
.Y(n_5872)
);

CKINVDCx5p33_ASAP7_75t_R g5873 ( 
.A(n_4258),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_4414),
.Y(n_5874)
);

CKINVDCx5p33_ASAP7_75t_R g5875 ( 
.A(n_4259),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_4419),
.Y(n_5876)
);

CKINVDCx5p33_ASAP7_75t_R g5877 ( 
.A(n_4261),
.Y(n_5877)
);

INVx1_ASAP7_75t_SL g5878 ( 
.A(n_4336),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_4420),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_4422),
.Y(n_5880)
);

CKINVDCx5p33_ASAP7_75t_R g5881 ( 
.A(n_4262),
.Y(n_5881)
);

CKINVDCx5p33_ASAP7_75t_R g5882 ( 
.A(n_4263),
.Y(n_5882)
);

CKINVDCx5p33_ASAP7_75t_R g5883 ( 
.A(n_4264),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_4429),
.Y(n_5884)
);

BUFx6f_ASAP7_75t_L g5885 ( 
.A(n_4971),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_4430),
.Y(n_5886)
);

NOR2xp67_ASAP7_75t_L g5887 ( 
.A(n_4824),
.B(n_2),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_4434),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_4445),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_4447),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_4453),
.Y(n_5891)
);

BUFx6f_ASAP7_75t_L g5892 ( 
.A(n_4971),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_4471),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_4477),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_4483),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_4493),
.Y(n_5896)
);

INVxp67_ASAP7_75t_L g5897 ( 
.A(n_4369),
.Y(n_5897)
);

CKINVDCx20_ASAP7_75t_R g5898 ( 
.A(n_4338),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_4507),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_4509),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_4521),
.Y(n_5901)
);

CKINVDCx5p33_ASAP7_75t_R g5902 ( 
.A(n_4265),
.Y(n_5902)
);

INVx1_ASAP7_75t_SL g5903 ( 
.A(n_4341),
.Y(n_5903)
);

CKINVDCx5p33_ASAP7_75t_R g5904 ( 
.A(n_4268),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_4539),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_4543),
.Y(n_5906)
);

CKINVDCx5p33_ASAP7_75t_R g5907 ( 
.A(n_4269),
.Y(n_5907)
);

CKINVDCx20_ASAP7_75t_R g5908 ( 
.A(n_4367),
.Y(n_5908)
);

CKINVDCx20_ASAP7_75t_R g5909 ( 
.A(n_4389),
.Y(n_5909)
);

CKINVDCx5p33_ASAP7_75t_R g5910 ( 
.A(n_4275),
.Y(n_5910)
);

INVx1_ASAP7_75t_L g5911 ( 
.A(n_4549),
.Y(n_5911)
);

INVx2_ASAP7_75t_L g5912 ( 
.A(n_5054),
.Y(n_5912)
);

CKINVDCx20_ASAP7_75t_R g5913 ( 
.A(n_4418),
.Y(n_5913)
);

CKINVDCx5p33_ASAP7_75t_R g5914 ( 
.A(n_4278),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_4550),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_4552),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_4553),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_4556),
.Y(n_5918)
);

CKINVDCx5p33_ASAP7_75t_R g5919 ( 
.A(n_4279),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_4557),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_4562),
.Y(n_5921)
);

CKINVDCx5p33_ASAP7_75t_R g5922 ( 
.A(n_4281),
.Y(n_5922)
);

CKINVDCx5p33_ASAP7_75t_R g5923 ( 
.A(n_4284),
.Y(n_5923)
);

BUFx6f_ASAP7_75t_L g5924 ( 
.A(n_5054),
.Y(n_5924)
);

INVxp67_ASAP7_75t_SL g5925 ( 
.A(n_5054),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_4564),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_4567),
.Y(n_5927)
);

BUFx10_ASAP7_75t_L g5928 ( 
.A(n_4364),
.Y(n_5928)
);

CKINVDCx5p33_ASAP7_75t_R g5929 ( 
.A(n_4285),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5119),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_4568),
.Y(n_5931)
);

CKINVDCx5p33_ASAP7_75t_R g5932 ( 
.A(n_4288),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_4571),
.Y(n_5933)
);

CKINVDCx5p33_ASAP7_75t_R g5934 ( 
.A(n_4289),
.Y(n_5934)
);

CKINVDCx5p33_ASAP7_75t_R g5935 ( 
.A(n_4291),
.Y(n_5935)
);

CKINVDCx5p33_ASAP7_75t_R g5936 ( 
.A(n_4294),
.Y(n_5936)
);

INVxp67_ASAP7_75t_L g5937 ( 
.A(n_4459),
.Y(n_5937)
);

INVx2_ASAP7_75t_L g5938 ( 
.A(n_5119),
.Y(n_5938)
);

INVx1_ASAP7_75t_L g5939 ( 
.A(n_4573),
.Y(n_5939)
);

BUFx3_ASAP7_75t_L g5940 ( 
.A(n_4326),
.Y(n_5940)
);

XNOR2xp5_ASAP7_75t_L g5941 ( 
.A(n_4920),
.B(n_5142),
.Y(n_5941)
);

HB1xp67_ASAP7_75t_L g5942 ( 
.A(n_4376),
.Y(n_5942)
);

BUFx2_ASAP7_75t_L g5943 ( 
.A(n_4510),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_4578),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_4579),
.Y(n_5945)
);

BUFx6f_ASAP7_75t_L g5946 ( 
.A(n_5119),
.Y(n_5946)
);

CKINVDCx5p33_ASAP7_75t_R g5947 ( 
.A(n_5511),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_4580),
.Y(n_5948)
);

CKINVDCx5p33_ASAP7_75t_R g5949 ( 
.A(n_4295),
.Y(n_5949)
);

CKINVDCx5p33_ASAP7_75t_R g5950 ( 
.A(n_4296),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_4585),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_4590),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_4602),
.Y(n_5953)
);

CKINVDCx5p33_ASAP7_75t_R g5954 ( 
.A(n_4298),
.Y(n_5954)
);

CKINVDCx5p33_ASAP7_75t_R g5955 ( 
.A(n_4300),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_4603),
.Y(n_5956)
);

CKINVDCx5p33_ASAP7_75t_R g5957 ( 
.A(n_4302),
.Y(n_5957)
);

HB1xp67_ASAP7_75t_L g5958 ( 
.A(n_4512),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_4611),
.Y(n_5959)
);

CKINVDCx5p33_ASAP7_75t_R g5960 ( 
.A(n_4303),
.Y(n_5960)
);

BUFx6f_ASAP7_75t_L g5961 ( 
.A(n_5152),
.Y(n_5961)
);

INVx1_ASAP7_75t_SL g5962 ( 
.A(n_4427),
.Y(n_5962)
);

NOR2xp33_ASAP7_75t_L g5963 ( 
.A(n_4548),
.B(n_3),
.Y(n_5963)
);

CKINVDCx5p33_ASAP7_75t_R g5964 ( 
.A(n_5510),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_4615),
.Y(n_5965)
);

INVx1_ASAP7_75t_SL g5966 ( 
.A(n_4433),
.Y(n_5966)
);

BUFx6f_ASAP7_75t_L g5967 ( 
.A(n_5152),
.Y(n_5967)
);

CKINVDCx20_ASAP7_75t_R g5968 ( 
.A(n_4446),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_4622),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_4624),
.Y(n_5970)
);

CKINVDCx5p33_ASAP7_75t_R g5971 ( 
.A(n_4305),
.Y(n_5971)
);

CKINVDCx5p33_ASAP7_75t_R g5972 ( 
.A(n_4306),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_4645),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_4658),
.Y(n_5974)
);

CKINVDCx5p33_ASAP7_75t_R g5975 ( 
.A(n_4307),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_4670),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_4679),
.Y(n_5977)
);

CKINVDCx5p33_ASAP7_75t_R g5978 ( 
.A(n_4308),
.Y(n_5978)
);

BUFx8_ASAP7_75t_SL g5979 ( 
.A(n_4746),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_4688),
.Y(n_5980)
);

INVx2_ASAP7_75t_L g5981 ( 
.A(n_5152),
.Y(n_5981)
);

HB1xp67_ASAP7_75t_L g5982 ( 
.A(n_4551),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_4692),
.Y(n_5983)
);

CKINVDCx5p33_ASAP7_75t_R g5984 ( 
.A(n_4311),
.Y(n_5984)
);

CKINVDCx5p33_ASAP7_75t_R g5985 ( 
.A(n_4315),
.Y(n_5985)
);

INVxp33_ASAP7_75t_L g5986 ( 
.A(n_4770),
.Y(n_5986)
);

INVx2_ASAP7_75t_SL g5987 ( 
.A(n_4696),
.Y(n_5987)
);

BUFx2_ASAP7_75t_L g5988 ( 
.A(n_4884),
.Y(n_5988)
);

CKINVDCx5p33_ASAP7_75t_R g5989 ( 
.A(n_4316),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_4693),
.Y(n_5990)
);

CKINVDCx5p33_ASAP7_75t_R g5991 ( 
.A(n_4318),
.Y(n_5991)
);

INVx1_ASAP7_75t_L g5992 ( 
.A(n_4703),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_4704),
.Y(n_5993)
);

CKINVDCx5p33_ASAP7_75t_R g5994 ( 
.A(n_4320),
.Y(n_5994)
);

BUFx10_ASAP7_75t_L g5995 ( 
.A(n_4591),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5732),
.Y(n_5996)
);

INVx2_ASAP7_75t_L g5997 ( 
.A(n_5560),
.Y(n_5997)
);

INVx2_ASAP7_75t_L g5998 ( 
.A(n_5560),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5742),
.Y(n_5999)
);

INVxp67_ASAP7_75t_L g6000 ( 
.A(n_5585),
.Y(n_6000)
);

INVxp33_ASAP7_75t_SL g6001 ( 
.A(n_5558),
.Y(n_6001)
);

INVx1_ASAP7_75t_L g6002 ( 
.A(n_5837),
.Y(n_6002)
);

INVxp67_ASAP7_75t_L g6003 ( 
.A(n_5942),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5848),
.Y(n_6004)
);

CKINVDCx5p33_ASAP7_75t_R g6005 ( 
.A(n_5559),
.Y(n_6005)
);

CKINVDCx5p33_ASAP7_75t_R g6006 ( 
.A(n_5564),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5925),
.Y(n_6007)
);

CKINVDCx20_ASAP7_75t_R g6008 ( 
.A(n_5663),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5551),
.Y(n_6009)
);

CKINVDCx20_ASAP7_75t_R g6010 ( 
.A(n_5670),
.Y(n_6010)
);

HB1xp67_ASAP7_75t_L g6011 ( 
.A(n_5573),
.Y(n_6011)
);

INVxp67_ASAP7_75t_SL g6012 ( 
.A(n_5567),
.Y(n_6012)
);

CKINVDCx20_ASAP7_75t_R g6013 ( 
.A(n_5676),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5552),
.Y(n_6014)
);

BUFx2_ASAP7_75t_SL g6015 ( 
.A(n_5566),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5555),
.Y(n_6016)
);

CKINVDCx5p33_ASAP7_75t_R g6017 ( 
.A(n_5568),
.Y(n_6017)
);

INVxp67_ASAP7_75t_SL g6018 ( 
.A(n_5606),
.Y(n_6018)
);

CKINVDCx5p33_ASAP7_75t_R g6019 ( 
.A(n_5572),
.Y(n_6019)
);

INVxp67_ASAP7_75t_SL g6020 ( 
.A(n_5623),
.Y(n_6020)
);

INVxp67_ASAP7_75t_L g6021 ( 
.A(n_5958),
.Y(n_6021)
);

BUFx3_ASAP7_75t_L g6022 ( 
.A(n_5649),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5556),
.Y(n_6023)
);

CKINVDCx20_ASAP7_75t_R g6024 ( 
.A(n_5695),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5557),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_5561),
.Y(n_6026)
);

CKINVDCx16_ASAP7_75t_R g6027 ( 
.A(n_5554),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5569),
.Y(n_6028)
);

INVx1_ASAP7_75t_L g6029 ( 
.A(n_5571),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5575),
.Y(n_6030)
);

INVx2_ASAP7_75t_L g6031 ( 
.A(n_5570),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_5587),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5589),
.Y(n_6033)
);

INVxp33_ASAP7_75t_L g6034 ( 
.A(n_5941),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5593),
.Y(n_6035)
);

CKINVDCx5p33_ASAP7_75t_R g6036 ( 
.A(n_5696),
.Y(n_6036)
);

CKINVDCx20_ASAP7_75t_R g6037 ( 
.A(n_5718),
.Y(n_6037)
);

INVx4_ASAP7_75t_R g6038 ( 
.A(n_5703),
.Y(n_6038)
);

CKINVDCx20_ASAP7_75t_R g6039 ( 
.A(n_5733),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5596),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5599),
.Y(n_6041)
);

BUFx2_ASAP7_75t_L g6042 ( 
.A(n_5574),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_5600),
.Y(n_6043)
);

CKINVDCx5p33_ASAP7_75t_R g6044 ( 
.A(n_5752),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5601),
.Y(n_6045)
);

CKINVDCx14_ASAP7_75t_R g6046 ( 
.A(n_5735),
.Y(n_6046)
);

INVxp67_ASAP7_75t_SL g6047 ( 
.A(n_5787),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_5570),
.Y(n_6048)
);

BUFx2_ASAP7_75t_L g6049 ( 
.A(n_5578),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5603),
.Y(n_6050)
);

CKINVDCx5p33_ASAP7_75t_R g6051 ( 
.A(n_5772),
.Y(n_6051)
);

HB1xp67_ASAP7_75t_L g6052 ( 
.A(n_5581),
.Y(n_6052)
);

CKINVDCx16_ASAP7_75t_R g6053 ( 
.A(n_5595),
.Y(n_6053)
);

CKINVDCx5p33_ASAP7_75t_R g6054 ( 
.A(n_5805),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5604),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5607),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5609),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5612),
.Y(n_6058)
);

INVxp67_ASAP7_75t_SL g6059 ( 
.A(n_5802),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5613),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_5615),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5616),
.Y(n_6062)
);

CKINVDCx20_ASAP7_75t_R g6063 ( 
.A(n_5832),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_5617),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5622),
.Y(n_6065)
);

INVxp67_ASAP7_75t_L g6066 ( 
.A(n_5982),
.Y(n_6066)
);

INVxp33_ASAP7_75t_SL g6067 ( 
.A(n_5584),
.Y(n_6067)
);

CKINVDCx20_ASAP7_75t_R g6068 ( 
.A(n_5860),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_5626),
.Y(n_6069)
);

CKINVDCx5p33_ASAP7_75t_R g6070 ( 
.A(n_5878),
.Y(n_6070)
);

INVx1_ASAP7_75t_L g6071 ( 
.A(n_5562),
.Y(n_6071)
);

CKINVDCx5p33_ASAP7_75t_R g6072 ( 
.A(n_5903),
.Y(n_6072)
);

HB1xp67_ASAP7_75t_L g6073 ( 
.A(n_5591),
.Y(n_6073)
);

CKINVDCx5p33_ASAP7_75t_R g6074 ( 
.A(n_5962),
.Y(n_6074)
);

INVxp67_ASAP7_75t_SL g6075 ( 
.A(n_5853),
.Y(n_6075)
);

CKINVDCx20_ASAP7_75t_R g6076 ( 
.A(n_5871),
.Y(n_6076)
);

INVxp67_ASAP7_75t_L g6077 ( 
.A(n_5966),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_5563),
.Y(n_6078)
);

CKINVDCx5p33_ASAP7_75t_R g6079 ( 
.A(n_5647),
.Y(n_6079)
);

INVxp67_ASAP7_75t_SL g6080 ( 
.A(n_5940),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5576),
.Y(n_6081)
);

INVx2_ASAP7_75t_L g6082 ( 
.A(n_5650),
.Y(n_6082)
);

INVxp33_ASAP7_75t_L g6083 ( 
.A(n_5979),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_5577),
.Y(n_6084)
);

CKINVDCx5p33_ASAP7_75t_R g6085 ( 
.A(n_5648),
.Y(n_6085)
);

BUFx3_ASAP7_75t_L g6086 ( 
.A(n_5553),
.Y(n_6086)
);

INVx1_ASAP7_75t_L g6087 ( 
.A(n_5579),
.Y(n_6087)
);

CKINVDCx20_ASAP7_75t_R g6088 ( 
.A(n_5898),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5580),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5583),
.Y(n_6090)
);

CKINVDCx5p33_ASAP7_75t_R g6091 ( 
.A(n_5651),
.Y(n_6091)
);

INVxp67_ASAP7_75t_L g6092 ( 
.A(n_5664),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_5586),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_5614),
.Y(n_6094)
);

CKINVDCx16_ASAP7_75t_R g6095 ( 
.A(n_5652),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_5704),
.Y(n_6096)
);

CKINVDCx20_ASAP7_75t_R g6097 ( 
.A(n_5908),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5671),
.Y(n_6098)
);

CKINVDCx20_ASAP7_75t_R g6099 ( 
.A(n_5909),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_5672),
.Y(n_6100)
);

INVxp67_ASAP7_75t_SL g6101 ( 
.A(n_5650),
.Y(n_6101)
);

HB1xp67_ASAP7_75t_L g6102 ( 
.A(n_5594),
.Y(n_6102)
);

INVxp67_ASAP7_75t_L g6103 ( 
.A(n_5943),
.Y(n_6103)
);

CKINVDCx16_ASAP7_75t_R g6104 ( 
.A(n_5706),
.Y(n_6104)
);

INVx1_ASAP7_75t_L g6105 ( 
.A(n_5673),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_5674),
.Y(n_6106)
);

INVx2_ASAP7_75t_L g6107 ( 
.A(n_5666),
.Y(n_6107)
);

CKINVDCx20_ASAP7_75t_R g6108 ( 
.A(n_5913),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_5677),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_5678),
.Y(n_6110)
);

INVxp67_ASAP7_75t_SL g6111 ( 
.A(n_5666),
.Y(n_6111)
);

INVx1_ASAP7_75t_L g6112 ( 
.A(n_5679),
.Y(n_6112)
);

INVxp67_ASAP7_75t_SL g6113 ( 
.A(n_5792),
.Y(n_6113)
);

CKINVDCx5p33_ASAP7_75t_R g6114 ( 
.A(n_5653),
.Y(n_6114)
);

CKINVDCx5p33_ASAP7_75t_R g6115 ( 
.A(n_5654),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_5681),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5682),
.Y(n_6117)
);

CKINVDCx5p33_ASAP7_75t_R g6118 ( 
.A(n_5655),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5684),
.Y(n_6119)
);

INVxp33_ASAP7_75t_L g6120 ( 
.A(n_5986),
.Y(n_6120)
);

INVx2_ASAP7_75t_L g6121 ( 
.A(n_5792),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5686),
.Y(n_6122)
);

INVx1_ASAP7_75t_SL g6123 ( 
.A(n_5605),
.Y(n_6123)
);

CKINVDCx5p33_ASAP7_75t_R g6124 ( 
.A(n_5657),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_5687),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5690),
.Y(n_6126)
);

CKINVDCx5p33_ASAP7_75t_R g6127 ( 
.A(n_5659),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5694),
.Y(n_6128)
);

CKINVDCx20_ASAP7_75t_R g6129 ( 
.A(n_5968),
.Y(n_6129)
);

BUFx3_ASAP7_75t_L g6130 ( 
.A(n_5795),
.Y(n_6130)
);

CKINVDCx5p33_ASAP7_75t_R g6131 ( 
.A(n_5660),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_5697),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_5701),
.Y(n_6133)
);

BUFx3_ASAP7_75t_L g6134 ( 
.A(n_5795),
.Y(n_6134)
);

CKINVDCx5p33_ASAP7_75t_R g6135 ( 
.A(n_5661),
.Y(n_6135)
);

CKINVDCx5p33_ASAP7_75t_R g6136 ( 
.A(n_5668),
.Y(n_6136)
);

CKINVDCx20_ASAP7_75t_R g6137 ( 
.A(n_5618),
.Y(n_6137)
);

CKINVDCx16_ASAP7_75t_R g6138 ( 
.A(n_5720),
.Y(n_6138)
);

CKINVDCx5p33_ASAP7_75t_R g6139 ( 
.A(n_5669),
.Y(n_6139)
);

INVxp33_ASAP7_75t_L g6140 ( 
.A(n_5643),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5705),
.Y(n_6141)
);

INVxp33_ASAP7_75t_SL g6142 ( 
.A(n_5597),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5708),
.Y(n_6143)
);

CKINVDCx5p33_ASAP7_75t_R g6144 ( 
.A(n_5675),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_5713),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_5715),
.Y(n_6146)
);

INVxp67_ASAP7_75t_SL g6147 ( 
.A(n_5803),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_5717),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_5723),
.Y(n_6149)
);

INVxp67_ASAP7_75t_SL g6150 ( 
.A(n_5803),
.Y(n_6150)
);

INVxp67_ASAP7_75t_SL g6151 ( 
.A(n_5822),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5729),
.Y(n_6152)
);

CKINVDCx5p33_ASAP7_75t_R g6153 ( 
.A(n_5680),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_5730),
.Y(n_6154)
);

INVx1_ASAP7_75t_L g6155 ( 
.A(n_5734),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5737),
.Y(n_6156)
);

CKINVDCx5p33_ASAP7_75t_R g6157 ( 
.A(n_5683),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_5822),
.Y(n_6158)
);

INVxp33_ASAP7_75t_SL g6159 ( 
.A(n_5598),
.Y(n_6159)
);

INVxp67_ASAP7_75t_L g6160 ( 
.A(n_5988),
.Y(n_6160)
);

INVxp67_ASAP7_75t_SL g6161 ( 
.A(n_5824),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5738),
.Y(n_6162)
);

CKINVDCx20_ASAP7_75t_R g6163 ( 
.A(n_5632),
.Y(n_6163)
);

CKINVDCx20_ASAP7_75t_R g6164 ( 
.A(n_5646),
.Y(n_6164)
);

CKINVDCx5p33_ASAP7_75t_R g6165 ( 
.A(n_5685),
.Y(n_6165)
);

CKINVDCx5p33_ASAP7_75t_R g6166 ( 
.A(n_5688),
.Y(n_6166)
);

CKINVDCx20_ASAP7_75t_R g6167 ( 
.A(n_5774),
.Y(n_6167)
);

CKINVDCx20_ASAP7_75t_R g6168 ( 
.A(n_5836),
.Y(n_6168)
);

CKINVDCx5p33_ASAP7_75t_R g6169 ( 
.A(n_5689),
.Y(n_6169)
);

CKINVDCx16_ASAP7_75t_R g6170 ( 
.A(n_5869),
.Y(n_6170)
);

CKINVDCx20_ASAP7_75t_R g6171 ( 
.A(n_5745),
.Y(n_6171)
);

CKINVDCx5p33_ASAP7_75t_R g6172 ( 
.A(n_5692),
.Y(n_6172)
);

INVxp67_ASAP7_75t_SL g6173 ( 
.A(n_5824),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_5740),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5743),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_5746),
.Y(n_6176)
);

CKINVDCx5p33_ASAP7_75t_R g6177 ( 
.A(n_5693),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_5748),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_5750),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_5754),
.Y(n_6180)
);

INVx1_ASAP7_75t_L g6181 ( 
.A(n_5756),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_5760),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_5761),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_5762),
.Y(n_6184)
);

HB1xp67_ASAP7_75t_L g6185 ( 
.A(n_5602),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5763),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_5764),
.Y(n_6187)
);

HB1xp67_ASAP7_75t_L g6188 ( 
.A(n_5608),
.Y(n_6188)
);

CKINVDCx14_ASAP7_75t_R g6189 ( 
.A(n_5755),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5765),
.Y(n_6190)
);

CKINVDCx5p33_ASAP7_75t_R g6191 ( 
.A(n_5698),
.Y(n_6191)
);

INVx2_ASAP7_75t_L g6192 ( 
.A(n_5851),
.Y(n_6192)
);

CKINVDCx5p33_ASAP7_75t_R g6193 ( 
.A(n_5699),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_5769),
.Y(n_6194)
);

CKINVDCx5p33_ASAP7_75t_R g6195 ( 
.A(n_5710),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5781),
.Y(n_6196)
);

INVxp67_ASAP7_75t_SL g6197 ( 
.A(n_5851),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_5782),
.Y(n_6198)
);

INVxp67_ASAP7_75t_L g6199 ( 
.A(n_5691),
.Y(n_6199)
);

CKINVDCx20_ASAP7_75t_R g6200 ( 
.A(n_5610),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_5785),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_5788),
.Y(n_6202)
);

CKINVDCx14_ASAP7_75t_R g6203 ( 
.A(n_5640),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_5789),
.Y(n_6204)
);

INVx3_ASAP7_75t_L g6205 ( 
.A(n_5885),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5790),
.Y(n_6206)
);

INVxp33_ASAP7_75t_SL g6207 ( 
.A(n_5611),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_5794),
.Y(n_6208)
);

INVxp67_ASAP7_75t_L g6209 ( 
.A(n_5582),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_5798),
.Y(n_6210)
);

CKINVDCx20_ASAP7_75t_R g6211 ( 
.A(n_5619),
.Y(n_6211)
);

CKINVDCx16_ASAP7_75t_R g6212 ( 
.A(n_5714),
.Y(n_6212)
);

CKINVDCx5p33_ASAP7_75t_R g6213 ( 
.A(n_5712),
.Y(n_6213)
);

CKINVDCx20_ASAP7_75t_R g6214 ( 
.A(n_5620),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_5800),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_5801),
.Y(n_6216)
);

INVxp67_ASAP7_75t_L g6217 ( 
.A(n_5634),
.Y(n_6217)
);

CKINVDCx5p33_ASAP7_75t_R g6218 ( 
.A(n_5716),
.Y(n_6218)
);

INVxp67_ASAP7_75t_SL g6219 ( 
.A(n_5885),
.Y(n_6219)
);

CKINVDCx5p33_ASAP7_75t_R g6220 ( 
.A(n_5721),
.Y(n_6220)
);

CKINVDCx5p33_ASAP7_75t_R g6221 ( 
.A(n_5722),
.Y(n_6221)
);

INVxp67_ASAP7_75t_L g6222 ( 
.A(n_5621),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5804),
.Y(n_6223)
);

CKINVDCx5p33_ASAP7_75t_R g6224 ( 
.A(n_5724),
.Y(n_6224)
);

CKINVDCx20_ASAP7_75t_R g6225 ( 
.A(n_5624),
.Y(n_6225)
);

INVx1_ASAP7_75t_L g6226 ( 
.A(n_5806),
.Y(n_6226)
);

INVx1_ASAP7_75t_L g6227 ( 
.A(n_5807),
.Y(n_6227)
);

INVx1_ASAP7_75t_L g6228 ( 
.A(n_5808),
.Y(n_6228)
);

CKINVDCx20_ASAP7_75t_R g6229 ( 
.A(n_5625),
.Y(n_6229)
);

INVxp33_ASAP7_75t_SL g6230 ( 
.A(n_5636),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5810),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_5811),
.Y(n_6232)
);

INVx1_ASAP7_75t_L g6233 ( 
.A(n_5814),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_5815),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_5819),
.Y(n_6235)
);

INVxp67_ASAP7_75t_SL g6236 ( 
.A(n_5892),
.Y(n_6236)
);

CKINVDCx5p33_ASAP7_75t_R g6237 ( 
.A(n_5725),
.Y(n_6237)
);

INVx2_ASAP7_75t_L g6238 ( 
.A(n_5892),
.Y(n_6238)
);

BUFx10_ASAP7_75t_L g6239 ( 
.A(n_5637),
.Y(n_6239)
);

INVx1_ASAP7_75t_L g6240 ( 
.A(n_5821),
.Y(n_6240)
);

CKINVDCx20_ASAP7_75t_R g6241 ( 
.A(n_5639),
.Y(n_6241)
);

INVxp33_ASAP7_75t_L g6242 ( 
.A(n_5840),
.Y(n_6242)
);

BUFx3_ASAP7_75t_L g6243 ( 
.A(n_5924),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_5827),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_5830),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_5841),
.Y(n_6246)
);

CKINVDCx16_ASAP7_75t_R g6247 ( 
.A(n_5826),
.Y(n_6247)
);

CKINVDCx5p33_ASAP7_75t_R g6248 ( 
.A(n_5726),
.Y(n_6248)
);

INVx2_ASAP7_75t_L g6249 ( 
.A(n_5924),
.Y(n_6249)
);

CKINVDCx20_ASAP7_75t_R g6250 ( 
.A(n_5728),
.Y(n_6250)
);

CKINVDCx5p33_ASAP7_75t_R g6251 ( 
.A(n_5736),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_5844),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_5845),
.Y(n_6253)
);

INVx2_ASAP7_75t_L g6254 ( 
.A(n_5946),
.Y(n_6254)
);

INVxp67_ASAP7_75t_SL g6255 ( 
.A(n_5946),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5850),
.Y(n_6256)
);

INVx1_ASAP7_75t_L g6257 ( 
.A(n_5854),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5857),
.Y(n_6258)
);

INVxp33_ASAP7_75t_SL g6259 ( 
.A(n_5739),
.Y(n_6259)
);

INVxp33_ASAP7_75t_SL g6260 ( 
.A(n_5741),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_5961),
.Y(n_6261)
);

INVxp67_ASAP7_75t_SL g6262 ( 
.A(n_5961),
.Y(n_6262)
);

CKINVDCx5p33_ASAP7_75t_R g6263 ( 
.A(n_5744),
.Y(n_6263)
);

CKINVDCx5p33_ASAP7_75t_R g6264 ( 
.A(n_5747),
.Y(n_6264)
);

CKINVDCx5p33_ASAP7_75t_R g6265 ( 
.A(n_5749),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_5859),
.Y(n_6266)
);

CKINVDCx5p33_ASAP7_75t_R g6267 ( 
.A(n_5751),
.Y(n_6267)
);

INVxp67_ASAP7_75t_SL g6268 ( 
.A(n_5967),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_5861),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_5862),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_5866),
.Y(n_6271)
);

CKINVDCx5p33_ASAP7_75t_R g6272 ( 
.A(n_5757),
.Y(n_6272)
);

INVx1_ASAP7_75t_L g6273 ( 
.A(n_5868),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5874),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_5876),
.Y(n_6275)
);

CKINVDCx5p33_ASAP7_75t_R g6276 ( 
.A(n_5758),
.Y(n_6276)
);

INVxp67_ASAP7_75t_SL g6277 ( 
.A(n_5967),
.Y(n_6277)
);

INVxp67_ASAP7_75t_SL g6278 ( 
.A(n_5768),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_5879),
.Y(n_6279)
);

CKINVDCx5p33_ASAP7_75t_R g6280 ( 
.A(n_5759),
.Y(n_6280)
);

CKINVDCx20_ASAP7_75t_R g6281 ( 
.A(n_5766),
.Y(n_6281)
);

CKINVDCx20_ASAP7_75t_R g6282 ( 
.A(n_5767),
.Y(n_6282)
);

INVxp67_ASAP7_75t_L g6283 ( 
.A(n_5770),
.Y(n_6283)
);

INVxp67_ASAP7_75t_L g6284 ( 
.A(n_5771),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_5880),
.Y(n_6285)
);

CKINVDCx16_ASAP7_75t_R g6286 ( 
.A(n_5849),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_5884),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_5886),
.Y(n_6288)
);

INVxp33_ASAP7_75t_SL g6289 ( 
.A(n_5773),
.Y(n_6289)
);

INVx1_ASAP7_75t_L g6290 ( 
.A(n_5888),
.Y(n_6290)
);

INVxp67_ASAP7_75t_SL g6291 ( 
.A(n_5963),
.Y(n_6291)
);

CKINVDCx5p33_ASAP7_75t_R g6292 ( 
.A(n_5775),
.Y(n_6292)
);

INVxp67_ASAP7_75t_L g6293 ( 
.A(n_5776),
.Y(n_6293)
);

INVxp67_ASAP7_75t_SL g6294 ( 
.A(n_5667),
.Y(n_6294)
);

INVxp67_ASAP7_75t_SL g6295 ( 
.A(n_5642),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_5889),
.Y(n_6296)
);

CKINVDCx5p33_ASAP7_75t_R g6297 ( 
.A(n_5777),
.Y(n_6297)
);

CKINVDCx5p33_ASAP7_75t_R g6298 ( 
.A(n_5778),
.Y(n_6298)
);

CKINVDCx20_ASAP7_75t_R g6299 ( 
.A(n_5780),
.Y(n_6299)
);

INVxp67_ASAP7_75t_L g6300 ( 
.A(n_5783),
.Y(n_6300)
);

BUFx6f_ASAP7_75t_L g6301 ( 
.A(n_5707),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_5890),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_5891),
.Y(n_6303)
);

INVx1_ASAP7_75t_SL g6304 ( 
.A(n_5645),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_5893),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_5894),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_5895),
.Y(n_6307)
);

INVx1_ASAP7_75t_L g6308 ( 
.A(n_5896),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_5899),
.Y(n_6309)
);

CKINVDCx5p33_ASAP7_75t_R g6310 ( 
.A(n_5784),
.Y(n_6310)
);

INVx2_ASAP7_75t_L g6311 ( 
.A(n_5592),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_5900),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_5901),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_5905),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_5906),
.Y(n_6315)
);

INVx2_ASAP7_75t_L g6316 ( 
.A(n_5592),
.Y(n_6316)
);

INVxp67_ASAP7_75t_SL g6317 ( 
.A(n_5829),
.Y(n_6317)
);

CKINVDCx5p33_ASAP7_75t_R g6318 ( 
.A(n_5786),
.Y(n_6318)
);

CKINVDCx5p33_ASAP7_75t_R g6319 ( 
.A(n_5791),
.Y(n_6319)
);

INVx1_ASAP7_75t_L g6320 ( 
.A(n_5911),
.Y(n_6320)
);

CKINVDCx5p33_ASAP7_75t_R g6321 ( 
.A(n_5793),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_5915),
.Y(n_6322)
);

HB1xp67_ASAP7_75t_L g6323 ( 
.A(n_5796),
.Y(n_6323)
);

CKINVDCx20_ASAP7_75t_R g6324 ( 
.A(n_5797),
.Y(n_6324)
);

CKINVDCx20_ASAP7_75t_R g6325 ( 
.A(n_5809),
.Y(n_6325)
);

CKINVDCx5p33_ASAP7_75t_R g6326 ( 
.A(n_5812),
.Y(n_6326)
);

CKINVDCx20_ASAP7_75t_R g6327 ( 
.A(n_5813),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_5916),
.Y(n_6328)
);

CKINVDCx5p33_ASAP7_75t_R g6329 ( 
.A(n_5816),
.Y(n_6329)
);

CKINVDCx20_ASAP7_75t_R g6330 ( 
.A(n_5817),
.Y(n_6330)
);

CKINVDCx20_ASAP7_75t_R g6331 ( 
.A(n_5818),
.Y(n_6331)
);

CKINVDCx5p33_ASAP7_75t_R g6332 ( 
.A(n_5823),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_5917),
.Y(n_6333)
);

CKINVDCx5p33_ASAP7_75t_R g6334 ( 
.A(n_5825),
.Y(n_6334)
);

CKINVDCx20_ASAP7_75t_R g6335 ( 
.A(n_5828),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_5918),
.Y(n_6336)
);

CKINVDCx5p33_ASAP7_75t_R g6337 ( 
.A(n_5831),
.Y(n_6337)
);

INVx1_ASAP7_75t_L g6338 ( 
.A(n_5920),
.Y(n_6338)
);

CKINVDCx5p33_ASAP7_75t_R g6339 ( 
.A(n_5833),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_5921),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_5926),
.Y(n_6341)
);

CKINVDCx5p33_ASAP7_75t_R g6342 ( 
.A(n_5834),
.Y(n_6342)
);

INVxp33_ASAP7_75t_SL g6343 ( 
.A(n_5835),
.Y(n_6343)
);

CKINVDCx20_ASAP7_75t_R g6344 ( 
.A(n_5839),
.Y(n_6344)
);

INVxp67_ASAP7_75t_SL g6345 ( 
.A(n_5565),
.Y(n_6345)
);

INVx2_ASAP7_75t_L g6346 ( 
.A(n_5592),
.Y(n_6346)
);

INVx1_ASAP7_75t_L g6347 ( 
.A(n_5927),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_5931),
.Y(n_6348)
);

INVxp33_ASAP7_75t_SL g6349 ( 
.A(n_5842),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_5933),
.Y(n_6350)
);

CKINVDCx16_ASAP7_75t_R g6351 ( 
.A(n_5928),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_5939),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_5944),
.Y(n_6353)
);

CKINVDCx5p33_ASAP7_75t_R g6354 ( 
.A(n_5843),
.Y(n_6354)
);

INVxp67_ASAP7_75t_SL g6355 ( 
.A(n_5719),
.Y(n_6355)
);

INVx1_ASAP7_75t_L g6356 ( 
.A(n_5945),
.Y(n_6356)
);

CKINVDCx16_ASAP7_75t_R g6357 ( 
.A(n_5995),
.Y(n_6357)
);

CKINVDCx5p33_ASAP7_75t_R g6358 ( 
.A(n_5846),
.Y(n_6358)
);

INVx1_ASAP7_75t_L g6359 ( 
.A(n_5948),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_5951),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_5952),
.Y(n_6361)
);

CKINVDCx20_ASAP7_75t_R g6362 ( 
.A(n_5847),
.Y(n_6362)
);

CKINVDCx20_ASAP7_75t_R g6363 ( 
.A(n_5852),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_5953),
.Y(n_6364)
);

CKINVDCx5p33_ASAP7_75t_R g6365 ( 
.A(n_5856),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_5956),
.Y(n_6366)
);

CKINVDCx5p33_ASAP7_75t_R g6367 ( 
.A(n_5858),
.Y(n_6367)
);

INVx1_ASAP7_75t_L g6368 ( 
.A(n_5959),
.Y(n_6368)
);

CKINVDCx5p33_ASAP7_75t_R g6369 ( 
.A(n_5863),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_5965),
.Y(n_6370)
);

CKINVDCx14_ASAP7_75t_R g6371 ( 
.A(n_5864),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_5969),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_5970),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_5973),
.Y(n_6374)
);

INVxp67_ASAP7_75t_SL g6375 ( 
.A(n_5731),
.Y(n_6375)
);

HB1xp67_ASAP7_75t_L g6376 ( 
.A(n_5865),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_5974),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_5976),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_5977),
.Y(n_6379)
);

CKINVDCx20_ASAP7_75t_R g6380 ( 
.A(n_5867),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_5980),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_5983),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_5990),
.Y(n_6383)
);

INVxp67_ASAP7_75t_L g6384 ( 
.A(n_5870),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_5992),
.Y(n_6385)
);

CKINVDCx5p33_ASAP7_75t_R g6386 ( 
.A(n_5872),
.Y(n_6386)
);

CKINVDCx20_ASAP7_75t_R g6387 ( 
.A(n_5873),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_5993),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_5628),
.Y(n_6389)
);

BUFx2_ASAP7_75t_L g6390 ( 
.A(n_5875),
.Y(n_6390)
);

CKINVDCx20_ASAP7_75t_R g6391 ( 
.A(n_5877),
.Y(n_6391)
);

INVx1_ASAP7_75t_SL g6392 ( 
.A(n_5881),
.Y(n_6392)
);

CKINVDCx20_ASAP7_75t_R g6393 ( 
.A(n_5882),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_5629),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_5630),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_5641),
.Y(n_6396)
);

CKINVDCx16_ASAP7_75t_R g6397 ( 
.A(n_5588),
.Y(n_6397)
);

CKINVDCx5p33_ASAP7_75t_R g6398 ( 
.A(n_5883),
.Y(n_6398)
);

BUFx3_ASAP7_75t_L g6399 ( 
.A(n_5592),
.Y(n_6399)
);

BUFx2_ASAP7_75t_L g6400 ( 
.A(n_5902),
.Y(n_6400)
);

INVx2_ASAP7_75t_L g6401 ( 
.A(n_5753),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_5644),
.Y(n_6402)
);

INVx1_ASAP7_75t_L g6403 ( 
.A(n_5656),
.Y(n_6403)
);

CKINVDCx20_ASAP7_75t_R g6404 ( 
.A(n_5904),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_5658),
.Y(n_6405)
);

HB1xp67_ASAP7_75t_L g6406 ( 
.A(n_5907),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_5662),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_5665),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_5590),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5709),
.Y(n_6410)
);

CKINVDCx16_ASAP7_75t_R g6411 ( 
.A(n_5627),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_5709),
.Y(n_6412)
);

INVx1_ASAP7_75t_L g6413 ( 
.A(n_5709),
.Y(n_6413)
);

INVxp67_ASAP7_75t_L g6414 ( 
.A(n_5910),
.Y(n_6414)
);

CKINVDCx5p33_ASAP7_75t_R g6415 ( 
.A(n_5914),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_5709),
.Y(n_6416)
);

CKINVDCx16_ASAP7_75t_R g6417 ( 
.A(n_5700),
.Y(n_6417)
);

CKINVDCx20_ASAP7_75t_R g6418 ( 
.A(n_5919),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_5631),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_5633),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5638),
.Y(n_6421)
);

INVx3_ASAP7_75t_L g6422 ( 
.A(n_5779),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_5820),
.Y(n_6423)
);

CKINVDCx5p33_ASAP7_75t_R g6424 ( 
.A(n_5922),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_5855),
.Y(n_6425)
);

INVxp67_ASAP7_75t_SL g6426 ( 
.A(n_5912),
.Y(n_6426)
);

INVx2_ASAP7_75t_L g6427 ( 
.A(n_5930),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_5938),
.Y(n_6428)
);

CKINVDCx20_ASAP7_75t_R g6429 ( 
.A(n_5923),
.Y(n_6429)
);

CKINVDCx5p33_ASAP7_75t_R g6430 ( 
.A(n_5929),
.Y(n_6430)
);

CKINVDCx5p33_ASAP7_75t_R g6431 ( 
.A(n_5932),
.Y(n_6431)
);

CKINVDCx20_ASAP7_75t_R g6432 ( 
.A(n_5934),
.Y(n_6432)
);

CKINVDCx5p33_ASAP7_75t_R g6433 ( 
.A(n_5935),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_5981),
.Y(n_6434)
);

CKINVDCx5p33_ASAP7_75t_R g6435 ( 
.A(n_5936),
.Y(n_6435)
);

CKINVDCx20_ASAP7_75t_R g6436 ( 
.A(n_5947),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_5711),
.Y(n_6437)
);

CKINVDCx20_ASAP7_75t_R g6438 ( 
.A(n_5949),
.Y(n_6438)
);

CKINVDCx5p33_ASAP7_75t_R g6439 ( 
.A(n_5950),
.Y(n_6439)
);

CKINVDCx20_ASAP7_75t_R g6440 ( 
.A(n_5954),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_5727),
.Y(n_6441)
);

CKINVDCx5p33_ASAP7_75t_R g6442 ( 
.A(n_5955),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_5887),
.Y(n_6443)
);

HB1xp67_ASAP7_75t_L g6444 ( 
.A(n_5957),
.Y(n_6444)
);

INVxp33_ASAP7_75t_SL g6445 ( 
.A(n_5960),
.Y(n_6445)
);

INVxp67_ASAP7_75t_L g6446 ( 
.A(n_5964),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_5971),
.Y(n_6447)
);

INVx2_ASAP7_75t_L g6448 ( 
.A(n_5972),
.Y(n_6448)
);

CKINVDCx5p33_ASAP7_75t_R g6449 ( 
.A(n_5975),
.Y(n_6449)
);

CKINVDCx20_ASAP7_75t_R g6450 ( 
.A(n_5978),
.Y(n_6450)
);

INVx1_ASAP7_75t_L g6451 ( 
.A(n_5984),
.Y(n_6451)
);

INVxp67_ASAP7_75t_SL g6452 ( 
.A(n_5897),
.Y(n_6452)
);

BUFx2_ASAP7_75t_L g6453 ( 
.A(n_5985),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_5989),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_5991),
.Y(n_6455)
);

CKINVDCx16_ASAP7_75t_R g6456 ( 
.A(n_5702),
.Y(n_6456)
);

CKINVDCx5p33_ASAP7_75t_R g6457 ( 
.A(n_5994),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_5799),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_5838),
.Y(n_6459)
);

BUFx3_ASAP7_75t_L g6460 ( 
.A(n_5987),
.Y(n_6460)
);

CKINVDCx5p33_ASAP7_75t_R g6461 ( 
.A(n_5635),
.Y(n_6461)
);

CKINVDCx5p33_ASAP7_75t_R g6462 ( 
.A(n_5937),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_5732),
.Y(n_6463)
);

CKINVDCx5p33_ASAP7_75t_R g6464 ( 
.A(n_5558),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_5732),
.Y(n_6465)
);

INVx1_ASAP7_75t_SL g6466 ( 
.A(n_5696),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_5732),
.Y(n_6467)
);

CKINVDCx20_ASAP7_75t_R g6468 ( 
.A(n_5663),
.Y(n_6468)
);

CKINVDCx20_ASAP7_75t_R g6469 ( 
.A(n_5663),
.Y(n_6469)
);

CKINVDCx5p33_ASAP7_75t_R g6470 ( 
.A(n_5558),
.Y(n_6470)
);

CKINVDCx5p33_ASAP7_75t_R g6471 ( 
.A(n_5558),
.Y(n_6471)
);

CKINVDCx5p33_ASAP7_75t_R g6472 ( 
.A(n_5558),
.Y(n_6472)
);

CKINVDCx5p33_ASAP7_75t_R g6473 ( 
.A(n_5558),
.Y(n_6473)
);

CKINVDCx5p33_ASAP7_75t_R g6474 ( 
.A(n_5558),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_5732),
.Y(n_6475)
);

HB1xp67_ASAP7_75t_L g6476 ( 
.A(n_5585),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_5732),
.Y(n_6477)
);

CKINVDCx14_ASAP7_75t_R g6478 ( 
.A(n_5735),
.Y(n_6478)
);

CKINVDCx5p33_ASAP7_75t_R g6479 ( 
.A(n_5558),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_5732),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_5732),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_5732),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_5732),
.Y(n_6483)
);

INVx2_ASAP7_75t_L g6484 ( 
.A(n_5560),
.Y(n_6484)
);

CKINVDCx20_ASAP7_75t_R g6485 ( 
.A(n_5663),
.Y(n_6485)
);

CKINVDCx20_ASAP7_75t_R g6486 ( 
.A(n_5663),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_5732),
.Y(n_6487)
);

CKINVDCx20_ASAP7_75t_R g6488 ( 
.A(n_5663),
.Y(n_6488)
);

CKINVDCx5p33_ASAP7_75t_R g6489 ( 
.A(n_5558),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_5732),
.Y(n_6490)
);

CKINVDCx20_ASAP7_75t_R g6491 ( 
.A(n_5663),
.Y(n_6491)
);

INVx1_ASAP7_75t_L g6492 ( 
.A(n_5732),
.Y(n_6492)
);

CKINVDCx5p33_ASAP7_75t_R g6493 ( 
.A(n_5558),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_5732),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_5732),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_5732),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_5732),
.Y(n_6497)
);

CKINVDCx20_ASAP7_75t_R g6498 ( 
.A(n_5663),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_5732),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_5732),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_5732),
.Y(n_6501)
);

CKINVDCx20_ASAP7_75t_R g6502 ( 
.A(n_5663),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_5732),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_5732),
.Y(n_6504)
);

INVxp67_ASAP7_75t_SL g6505 ( 
.A(n_5732),
.Y(n_6505)
);

CKINVDCx5p33_ASAP7_75t_R g6506 ( 
.A(n_5558),
.Y(n_6506)
);

BUFx3_ASAP7_75t_L g6507 ( 
.A(n_5567),
.Y(n_6507)
);

INVx1_ASAP7_75t_L g6508 ( 
.A(n_5732),
.Y(n_6508)
);

CKINVDCx5p33_ASAP7_75t_R g6509 ( 
.A(n_5558),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_5732),
.Y(n_6510)
);

CKINVDCx20_ASAP7_75t_R g6511 ( 
.A(n_5663),
.Y(n_6511)
);

INVx3_ASAP7_75t_L g6512 ( 
.A(n_6022),
.Y(n_6512)
);

AND2x2_ASAP7_75t_L g6513 ( 
.A(n_6140),
.B(n_4954),
.Y(n_6513)
);

INVx2_ASAP7_75t_L g6514 ( 
.A(n_6301),
.Y(n_6514)
);

BUFx6f_ASAP7_75t_L g6515 ( 
.A(n_6507),
.Y(n_6515)
);

CKINVDCx5p33_ASAP7_75t_R g6516 ( 
.A(n_6079),
.Y(n_6516)
);

HB1xp67_ASAP7_75t_L g6517 ( 
.A(n_6011),
.Y(n_6517)
);

INVx2_ASAP7_75t_L g6518 ( 
.A(n_6301),
.Y(n_6518)
);

AND2x4_ASAP7_75t_L g6519 ( 
.A(n_6460),
.B(n_5006),
.Y(n_6519)
);

INVx2_ASAP7_75t_L g6520 ( 
.A(n_6301),
.Y(n_6520)
);

BUFx6f_ASAP7_75t_L g6521 ( 
.A(n_6130),
.Y(n_6521)
);

INVx2_ASAP7_75t_L g6522 ( 
.A(n_6419),
.Y(n_6522)
);

INVx1_ASAP7_75t_L g6523 ( 
.A(n_6009),
.Y(n_6523)
);

AND2x2_ASAP7_75t_L g6524 ( 
.A(n_6120),
.B(n_5027),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6014),
.Y(n_6525)
);

BUFx6f_ASAP7_75t_L g6526 ( 
.A(n_6134),
.Y(n_6526)
);

INVx1_ASAP7_75t_L g6527 ( 
.A(n_6098),
.Y(n_6527)
);

INVx2_ASAP7_75t_L g6528 ( 
.A(n_6420),
.Y(n_6528)
);

BUFx6f_ASAP7_75t_L g6529 ( 
.A(n_6243),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_6100),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6105),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_6106),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_6421),
.Y(n_6533)
);

OAI22xp5_ASAP7_75t_SL g6534 ( 
.A1(n_6242),
.A2(n_4450),
.B1(n_4454),
.B2(n_4449),
.Y(n_6534)
);

BUFx6f_ASAP7_75t_L g6535 ( 
.A(n_6036),
.Y(n_6535)
);

INVx2_ASAP7_75t_L g6536 ( 
.A(n_6401),
.Y(n_6536)
);

INVx2_ASAP7_75t_L g6537 ( 
.A(n_6427),
.Y(n_6537)
);

INVx3_ASAP7_75t_L g6538 ( 
.A(n_6086),
.Y(n_6538)
);

INVx2_ASAP7_75t_L g6539 ( 
.A(n_6071),
.Y(n_6539)
);

INVx1_ASAP7_75t_L g6540 ( 
.A(n_6109),
.Y(n_6540)
);

AND2x6_ASAP7_75t_L g6541 ( 
.A(n_6392),
.B(n_4848),
.Y(n_6541)
);

INVx3_ASAP7_75t_L g6542 ( 
.A(n_6466),
.Y(n_6542)
);

AOI22xp5_ASAP7_75t_L g6543 ( 
.A1(n_6278),
.A2(n_4667),
.B1(n_4699),
.B2(n_4639),
.Y(n_6543)
);

INVx4_ASAP7_75t_L g6544 ( 
.A(n_6085),
.Y(n_6544)
);

BUFx6f_ASAP7_75t_L g6545 ( 
.A(n_6044),
.Y(n_6545)
);

INVx3_ASAP7_75t_L g6546 ( 
.A(n_6205),
.Y(n_6546)
);

BUFx2_ASAP7_75t_L g6547 ( 
.A(n_6462),
.Y(n_6547)
);

CKINVDCx5p33_ASAP7_75t_R g6548 ( 
.A(n_6091),
.Y(n_6548)
);

NAND2xp5_ASAP7_75t_L g6549 ( 
.A(n_6409),
.B(n_5156),
.Y(n_6549)
);

NAND2xp5_ASAP7_75t_L g6550 ( 
.A(n_6291),
.B(n_6016),
.Y(n_6550)
);

NAND2xp5_ASAP7_75t_SL g6551 ( 
.A(n_6259),
.B(n_4333),
.Y(n_6551)
);

INVx2_ASAP7_75t_L g6552 ( 
.A(n_6078),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_6110),
.Y(n_6553)
);

INVx2_ASAP7_75t_L g6554 ( 
.A(n_6081),
.Y(n_6554)
);

AND2x4_ASAP7_75t_L g6555 ( 
.A(n_6077),
.B(n_5099),
.Y(n_6555)
);

BUFx3_ASAP7_75t_L g6556 ( 
.A(n_6250),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6112),
.Y(n_6557)
);

BUFx6f_ASAP7_75t_L g6558 ( 
.A(n_6051),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_6084),
.Y(n_6559)
);

INVx2_ASAP7_75t_L g6560 ( 
.A(n_6087),
.Y(n_6560)
);

NAND2xp5_ASAP7_75t_L g6561 ( 
.A(n_6023),
.B(n_5156),
.Y(n_6561)
);

BUFx6f_ASAP7_75t_L g6562 ( 
.A(n_6054),
.Y(n_6562)
);

BUFx6f_ASAP7_75t_L g6563 ( 
.A(n_6070),
.Y(n_6563)
);

INVx2_ASAP7_75t_L g6564 ( 
.A(n_6089),
.Y(n_6564)
);

NAND2xp33_ASAP7_75t_L g6565 ( 
.A(n_6114),
.B(n_6115),
.Y(n_6565)
);

INVx4_ASAP7_75t_L g6566 ( 
.A(n_6118),
.Y(n_6566)
);

INVx3_ASAP7_75t_L g6567 ( 
.A(n_6205),
.Y(n_6567)
);

AND2x4_ASAP7_75t_L g6568 ( 
.A(n_6012),
.B(n_5108),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6116),
.Y(n_6569)
);

OAI22xp5_ASAP7_75t_SL g6570 ( 
.A1(n_6008),
.A2(n_4488),
.B1(n_4526),
.B2(n_4487),
.Y(n_6570)
);

INVx2_ASAP7_75t_L g6571 ( 
.A(n_6090),
.Y(n_6571)
);

AOI22xp5_ASAP7_75t_L g6572 ( 
.A1(n_6295),
.A2(n_4845),
.B1(n_4856),
.B2(n_4735),
.Y(n_6572)
);

XNOR2x2_ASAP7_75t_L g6573 ( 
.A(n_6123),
.B(n_5386),
.Y(n_6573)
);

INVx1_ASAP7_75t_L g6574 ( 
.A(n_6117),
.Y(n_6574)
);

AND2x2_ASAP7_75t_L g6575 ( 
.A(n_6452),
.B(n_5189),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6119),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6122),
.Y(n_6577)
);

INVx2_ASAP7_75t_L g6578 ( 
.A(n_6093),
.Y(n_6578)
);

NAND2xp5_ASAP7_75t_L g6579 ( 
.A(n_6025),
.B(n_5156),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_6125),
.Y(n_6580)
);

HB1xp67_ASAP7_75t_L g6581 ( 
.A(n_6476),
.Y(n_6581)
);

BUFx6f_ASAP7_75t_L g6582 ( 
.A(n_6072),
.Y(n_6582)
);

HB1xp67_ASAP7_75t_L g6583 ( 
.A(n_6000),
.Y(n_6583)
);

AND2x4_ASAP7_75t_L g6584 ( 
.A(n_6018),
.B(n_5286),
.Y(n_6584)
);

INVx2_ASAP7_75t_L g6585 ( 
.A(n_6094),
.Y(n_6585)
);

CKINVDCx5p33_ASAP7_75t_R g6586 ( 
.A(n_6124),
.Y(n_6586)
);

AND2x4_ASAP7_75t_L g6587 ( 
.A(n_6020),
.B(n_6047),
.Y(n_6587)
);

HB1xp67_ASAP7_75t_L g6588 ( 
.A(n_6092),
.Y(n_6588)
);

BUFx2_ASAP7_75t_L g6589 ( 
.A(n_6281),
.Y(n_6589)
);

OAI22xp5_ASAP7_75t_SL g6590 ( 
.A1(n_6010),
.A2(n_4559),
.B1(n_4581),
.B2(n_4534),
.Y(n_6590)
);

INVx2_ASAP7_75t_L g6591 ( 
.A(n_6311),
.Y(n_6591)
);

INVx3_ASAP7_75t_L g6592 ( 
.A(n_6096),
.Y(n_6592)
);

AND2x4_ASAP7_75t_L g6593 ( 
.A(n_6059),
.B(n_6075),
.Y(n_6593)
);

AND2x2_ASAP7_75t_L g6594 ( 
.A(n_6371),
.B(n_5289),
.Y(n_6594)
);

INVx2_ASAP7_75t_L g6595 ( 
.A(n_6316),
.Y(n_6595)
);

INVx3_ASAP7_75t_L g6596 ( 
.A(n_6074),
.Y(n_6596)
);

INVx3_ASAP7_75t_L g6597 ( 
.A(n_6422),
.Y(n_6597)
);

BUFx3_ASAP7_75t_L g6598 ( 
.A(n_6282),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6126),
.Y(n_6599)
);

INVx2_ASAP7_75t_L g6600 ( 
.A(n_6346),
.Y(n_6600)
);

INVx1_ASAP7_75t_L g6601 ( 
.A(n_6128),
.Y(n_6601)
);

AND2x4_ASAP7_75t_L g6602 ( 
.A(n_6080),
.B(n_5312),
.Y(n_6602)
);

AND2x4_ASAP7_75t_L g6603 ( 
.A(n_6304),
.B(n_4332),
.Y(n_6603)
);

NAND2xp5_ASAP7_75t_L g6604 ( 
.A(n_6026),
.B(n_6028),
.Y(n_6604)
);

OAI22x1_ASAP7_75t_R g6605 ( 
.A1(n_6299),
.A2(n_6325),
.B1(n_6327),
.B2(n_6324),
.Y(n_6605)
);

NOR2x1_ASAP7_75t_L g6606 ( 
.A(n_6447),
.B(n_4474),
.Y(n_6606)
);

OA21x2_ASAP7_75t_L g6607 ( 
.A1(n_6410),
.A2(n_4719),
.B(n_4712),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6132),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6133),
.Y(n_6609)
);

INVx1_ASAP7_75t_L g6610 ( 
.A(n_6141),
.Y(n_6610)
);

INVx2_ASAP7_75t_L g6611 ( 
.A(n_6422),
.Y(n_6611)
);

INVx2_ASAP7_75t_L g6612 ( 
.A(n_6423),
.Y(n_6612)
);

OAI21x1_ASAP7_75t_L g6613 ( 
.A1(n_6412),
.A2(n_4224),
.B(n_4212),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6143),
.Y(n_6614)
);

NAND2xp5_ASAP7_75t_L g6615 ( 
.A(n_6029),
.B(n_5175),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_6030),
.B(n_5175),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_6145),
.Y(n_6617)
);

INVx1_ASAP7_75t_L g6618 ( 
.A(n_6146),
.Y(n_6618)
);

AND2x2_ASAP7_75t_L g6619 ( 
.A(n_6003),
.B(n_6021),
.Y(n_6619)
);

INVx2_ASAP7_75t_L g6620 ( 
.A(n_6425),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6148),
.Y(n_6621)
);

INVx2_ASAP7_75t_L g6622 ( 
.A(n_6428),
.Y(n_6622)
);

NAND2xp5_ASAP7_75t_L g6623 ( 
.A(n_6032),
.B(n_6033),
.Y(n_6623)
);

AND2x4_ASAP7_75t_L g6624 ( 
.A(n_6390),
.B(n_4485),
.Y(n_6624)
);

INVx5_ASAP7_75t_L g6625 ( 
.A(n_6095),
.Y(n_6625)
);

INVx2_ASAP7_75t_L g6626 ( 
.A(n_6434),
.Y(n_6626)
);

OA21x2_ASAP7_75t_L g6627 ( 
.A1(n_6413),
.A2(n_4731),
.B(n_4720),
.Y(n_6627)
);

INVx2_ASAP7_75t_L g6628 ( 
.A(n_6035),
.Y(n_6628)
);

BUFx3_ASAP7_75t_L g6629 ( 
.A(n_6330),
.Y(n_6629)
);

AND2x4_ASAP7_75t_L g6630 ( 
.A(n_6400),
.B(n_6453),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6066),
.B(n_4721),
.Y(n_6631)
);

NOR2xp33_ASAP7_75t_L g6632 ( 
.A(n_6448),
.B(n_4136),
.Y(n_6632)
);

BUFx6f_ASAP7_75t_L g6633 ( 
.A(n_6239),
.Y(n_6633)
);

BUFx6f_ASAP7_75t_L g6634 ( 
.A(n_6239),
.Y(n_6634)
);

NOR2xp33_ASAP7_75t_L g6635 ( 
.A(n_6451),
.B(n_4172),
.Y(n_6635)
);

BUFx6f_ASAP7_75t_L g6636 ( 
.A(n_5997),
.Y(n_6636)
);

BUFx6f_ASAP7_75t_L g6637 ( 
.A(n_5998),
.Y(n_6637)
);

INVx3_ASAP7_75t_L g6638 ( 
.A(n_6389),
.Y(n_6638)
);

AND2x4_ASAP7_75t_L g6639 ( 
.A(n_6042),
.B(n_4496),
.Y(n_6639)
);

OAI22xp5_ASAP7_75t_L g6640 ( 
.A1(n_6317),
.A2(n_4921),
.B1(n_4983),
.B2(n_4865),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_6149),
.Y(n_6641)
);

NOR2xp33_ASAP7_75t_L g6642 ( 
.A(n_6454),
.B(n_4203),
.Y(n_6642)
);

INVx3_ASAP7_75t_L g6643 ( 
.A(n_6394),
.Y(n_6643)
);

OAI22xp5_ASAP7_75t_L g6644 ( 
.A1(n_6455),
.A2(n_6283),
.B1(n_6293),
.B2(n_6284),
.Y(n_6644)
);

INVx2_ASAP7_75t_L g6645 ( 
.A(n_6040),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6152),
.Y(n_6646)
);

BUFx6f_ASAP7_75t_L g6647 ( 
.A(n_6031),
.Y(n_6647)
);

OAI22x1_ASAP7_75t_L g6648 ( 
.A1(n_6103),
.A2(n_4713),
.B1(n_4995),
.B2(n_4991),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6154),
.Y(n_6649)
);

INVx2_ASAP7_75t_L g6650 ( 
.A(n_6041),
.Y(n_6650)
);

BUFx6f_ASAP7_75t_L g6651 ( 
.A(n_6048),
.Y(n_6651)
);

INVx3_ASAP7_75t_L g6652 ( 
.A(n_6395),
.Y(n_6652)
);

AND2x4_ASAP7_75t_L g6653 ( 
.A(n_6049),
.B(n_4599),
.Y(n_6653)
);

INVx6_ASAP7_75t_L g6654 ( 
.A(n_6397),
.Y(n_6654)
);

BUFx12f_ASAP7_75t_L g6655 ( 
.A(n_6005),
.Y(n_6655)
);

BUFx2_ASAP7_75t_L g6656 ( 
.A(n_6331),
.Y(n_6656)
);

INVx2_ASAP7_75t_L g6657 ( 
.A(n_6043),
.Y(n_6657)
);

INVx2_ASAP7_75t_L g6658 ( 
.A(n_6045),
.Y(n_6658)
);

AND2x2_ASAP7_75t_SL g6659 ( 
.A(n_6027),
.B(n_4310),
.Y(n_6659)
);

BUFx6f_ASAP7_75t_L g6660 ( 
.A(n_6082),
.Y(n_6660)
);

BUFx6f_ASAP7_75t_L g6661 ( 
.A(n_6107),
.Y(n_6661)
);

BUFx6f_ASAP7_75t_L g6662 ( 
.A(n_6121),
.Y(n_6662)
);

INVx3_ASAP7_75t_L g6663 ( 
.A(n_6396),
.Y(n_6663)
);

INVx5_ASAP7_75t_L g6664 ( 
.A(n_6104),
.Y(n_6664)
);

HB1xp67_ASAP7_75t_L g6665 ( 
.A(n_6160),
.Y(n_6665)
);

INVx4_ASAP7_75t_L g6666 ( 
.A(n_6127),
.Y(n_6666)
);

AND2x2_ASAP7_75t_L g6667 ( 
.A(n_6199),
.B(n_4721),
.Y(n_6667)
);

INVx6_ASAP7_75t_L g6668 ( 
.A(n_6411),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6050),
.Y(n_6669)
);

BUFx2_ASAP7_75t_L g6670 ( 
.A(n_6335),
.Y(n_6670)
);

INVxp67_ASAP7_75t_L g6671 ( 
.A(n_6015),
.Y(n_6671)
);

NAND2xp5_ASAP7_75t_L g6672 ( 
.A(n_6055),
.B(n_5175),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6056),
.Y(n_6673)
);

INVxp67_ASAP7_75t_L g6674 ( 
.A(n_6052),
.Y(n_6674)
);

BUFx6f_ASAP7_75t_L g6675 ( 
.A(n_6158),
.Y(n_6675)
);

AND2x4_ASAP7_75t_L g6676 ( 
.A(n_6209),
.B(n_4625),
.Y(n_6676)
);

NOR2x1_ASAP7_75t_L g6677 ( 
.A(n_6458),
.B(n_4727),
.Y(n_6677)
);

INVx3_ASAP7_75t_L g6678 ( 
.A(n_6402),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_6155),
.Y(n_6679)
);

BUFx6f_ASAP7_75t_L g6680 ( 
.A(n_6192),
.Y(n_6680)
);

OAI21x1_ASAP7_75t_L g6681 ( 
.A1(n_6416),
.A2(n_4353),
.B(n_4324),
.Y(n_6681)
);

BUFx6f_ASAP7_75t_L g6682 ( 
.A(n_6238),
.Y(n_6682)
);

CKINVDCx6p67_ASAP7_75t_R g6683 ( 
.A(n_6344),
.Y(n_6683)
);

INVx4_ASAP7_75t_L g6684 ( 
.A(n_6131),
.Y(n_6684)
);

CKINVDCx5p33_ASAP7_75t_R g6685 ( 
.A(n_6135),
.Y(n_6685)
);

CKINVDCx5p33_ASAP7_75t_R g6686 ( 
.A(n_6136),
.Y(n_6686)
);

BUFx6f_ASAP7_75t_L g6687 ( 
.A(n_6249),
.Y(n_6687)
);

INVx5_ASAP7_75t_L g6688 ( 
.A(n_6138),
.Y(n_6688)
);

BUFx2_ASAP7_75t_L g6689 ( 
.A(n_6362),
.Y(n_6689)
);

INVx6_ASAP7_75t_L g6690 ( 
.A(n_6417),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6156),
.Y(n_6691)
);

BUFx6f_ASAP7_75t_L g6692 ( 
.A(n_6254),
.Y(n_6692)
);

INVx6_ASAP7_75t_L g6693 ( 
.A(n_6456),
.Y(n_6693)
);

INVx1_ASAP7_75t_L g6694 ( 
.A(n_6162),
.Y(n_6694)
);

BUFx6f_ASAP7_75t_L g6695 ( 
.A(n_6261),
.Y(n_6695)
);

OA21x2_ASAP7_75t_L g6696 ( 
.A1(n_6057),
.A2(n_4740),
.B(n_4736),
.Y(n_6696)
);

NAND2xp5_ASAP7_75t_L g6697 ( 
.A(n_6058),
.B(n_5328),
.Y(n_6697)
);

INVx2_ASAP7_75t_L g6698 ( 
.A(n_6060),
.Y(n_6698)
);

HB1xp67_ASAP7_75t_L g6699 ( 
.A(n_6139),
.Y(n_6699)
);

INVx2_ASAP7_75t_L g6700 ( 
.A(n_6061),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_6062),
.Y(n_6701)
);

BUFx2_ASAP7_75t_L g6702 ( 
.A(n_6363),
.Y(n_6702)
);

CKINVDCx8_ASAP7_75t_R g6703 ( 
.A(n_6170),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_L g6704 ( 
.A(n_6064),
.B(n_5328),
.Y(n_6704)
);

NAND2xp5_ASAP7_75t_L g6705 ( 
.A(n_6065),
.B(n_5328),
.Y(n_6705)
);

OAI22xp5_ASAP7_75t_SL g6706 ( 
.A1(n_6013),
.A2(n_4601),
.B1(n_4619),
.B2(n_4583),
.Y(n_6706)
);

OA21x2_ASAP7_75t_L g6707 ( 
.A1(n_6069),
.A2(n_4747),
.B(n_4741),
.Y(n_6707)
);

INVx2_ASAP7_75t_L g6708 ( 
.A(n_5996),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6174),
.Y(n_6709)
);

INVx3_ASAP7_75t_L g6710 ( 
.A(n_6403),
.Y(n_6710)
);

AND2x4_ASAP7_75t_L g6711 ( 
.A(n_6217),
.B(n_4755),
.Y(n_6711)
);

INVx2_ASAP7_75t_L g6712 ( 
.A(n_5999),
.Y(n_6712)
);

BUFx6f_ASAP7_75t_L g6713 ( 
.A(n_6484),
.Y(n_6713)
);

BUFx6f_ASAP7_75t_L g6714 ( 
.A(n_6006),
.Y(n_6714)
);

AND2x2_ASAP7_75t_L g6715 ( 
.A(n_6203),
.B(n_4757),
.Y(n_6715)
);

BUFx12f_ASAP7_75t_L g6716 ( 
.A(n_6017),
.Y(n_6716)
);

BUFx2_ASAP7_75t_L g6717 ( 
.A(n_6380),
.Y(n_6717)
);

INVx5_ASAP7_75t_L g6718 ( 
.A(n_6212),
.Y(n_6718)
);

INVx5_ASAP7_75t_L g6719 ( 
.A(n_6247),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6175),
.Y(n_6720)
);

INVx3_ASAP7_75t_L g6721 ( 
.A(n_6405),
.Y(n_6721)
);

BUFx6f_ASAP7_75t_L g6722 ( 
.A(n_6019),
.Y(n_6722)
);

HB1xp67_ASAP7_75t_L g6723 ( 
.A(n_6144),
.Y(n_6723)
);

INVx2_ASAP7_75t_SL g6724 ( 
.A(n_6153),
.Y(n_6724)
);

AND2x4_ASAP7_75t_L g6725 ( 
.A(n_6222),
.B(n_4772),
.Y(n_6725)
);

BUFx6f_ASAP7_75t_L g6726 ( 
.A(n_6464),
.Y(n_6726)
);

BUFx12f_ASAP7_75t_L g6727 ( 
.A(n_6470),
.Y(n_6727)
);

INVxp33_ASAP7_75t_SL g6728 ( 
.A(n_6471),
.Y(n_6728)
);

INVx2_ASAP7_75t_L g6729 ( 
.A(n_6002),
.Y(n_6729)
);

BUFx12f_ASAP7_75t_L g6730 ( 
.A(n_6472),
.Y(n_6730)
);

BUFx2_ASAP7_75t_L g6731 ( 
.A(n_6387),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6176),
.Y(n_6732)
);

INVx2_ASAP7_75t_L g6733 ( 
.A(n_6004),
.Y(n_6733)
);

AND2x2_ASAP7_75t_L g6734 ( 
.A(n_6046),
.B(n_4757),
.Y(n_6734)
);

NAND2xp5_ASAP7_75t_L g6735 ( 
.A(n_6505),
.B(n_5345),
.Y(n_6735)
);

BUFx6f_ASAP7_75t_L g6736 ( 
.A(n_6473),
.Y(n_6736)
);

BUFx6f_ASAP7_75t_L g6737 ( 
.A(n_6474),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6178),
.Y(n_6738)
);

BUFx8_ASAP7_75t_L g6739 ( 
.A(n_6459),
.Y(n_6739)
);

AOI22xp5_ASAP7_75t_L g6740 ( 
.A1(n_6345),
.A2(n_5266),
.B1(n_5268),
.B2(n_5033),
.Y(n_6740)
);

INVx3_ASAP7_75t_L g6741 ( 
.A(n_6407),
.Y(n_6741)
);

INVx2_ASAP7_75t_L g6742 ( 
.A(n_6007),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_SL g6743 ( 
.A(n_6260),
.B(n_4334),
.Y(n_6743)
);

AND2x2_ASAP7_75t_L g6744 ( 
.A(n_6189),
.B(n_4761),
.Y(n_6744)
);

NAND2xp5_ASAP7_75t_L g6745 ( 
.A(n_6399),
.B(n_6463),
.Y(n_6745)
);

INVx2_ASAP7_75t_L g6746 ( 
.A(n_6465),
.Y(n_6746)
);

CKINVDCx20_ASAP7_75t_R g6747 ( 
.A(n_6024),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6467),
.Y(n_6748)
);

CKINVDCx20_ASAP7_75t_R g6749 ( 
.A(n_6037),
.Y(n_6749)
);

INVx2_ASAP7_75t_L g6750 ( 
.A(n_6475),
.Y(n_6750)
);

OAI22x1_ASAP7_75t_SL g6751 ( 
.A1(n_6391),
.A2(n_4631),
.B1(n_4635),
.B2(n_4628),
.Y(n_6751)
);

NAND2xp5_ASAP7_75t_L g6752 ( 
.A(n_6477),
.B(n_5345),
.Y(n_6752)
);

NAND2xp5_ASAP7_75t_L g6753 ( 
.A(n_6480),
.B(n_6481),
.Y(n_6753)
);

AND2x4_ASAP7_75t_L g6754 ( 
.A(n_6300),
.B(n_6384),
.Y(n_6754)
);

INVx1_ASAP7_75t_L g6755 ( 
.A(n_6179),
.Y(n_6755)
);

BUFx6f_ASAP7_75t_L g6756 ( 
.A(n_6479),
.Y(n_6756)
);

BUFx3_ASAP7_75t_L g6757 ( 
.A(n_6393),
.Y(n_6757)
);

BUFx12f_ASAP7_75t_L g6758 ( 
.A(n_6489),
.Y(n_6758)
);

INVx2_ASAP7_75t_L g6759 ( 
.A(n_6482),
.Y(n_6759)
);

OAI22xp5_ASAP7_75t_L g6760 ( 
.A1(n_6414),
.A2(n_5346),
.B1(n_5294),
.B2(n_4955),
.Y(n_6760)
);

INVx3_ASAP7_75t_L g6761 ( 
.A(n_6408),
.Y(n_6761)
);

NOR2xp33_ASAP7_75t_L g6762 ( 
.A(n_6483),
.B(n_4271),
.Y(n_6762)
);

INVxp67_ASAP7_75t_L g6763 ( 
.A(n_6073),
.Y(n_6763)
);

AND2x4_ASAP7_75t_L g6764 ( 
.A(n_6446),
.B(n_4869),
.Y(n_6764)
);

INVx2_ASAP7_75t_L g6765 ( 
.A(n_6487),
.Y(n_6765)
);

INVx2_ASAP7_75t_L g6766 ( 
.A(n_6490),
.Y(n_6766)
);

INVx1_ASAP7_75t_L g6767 ( 
.A(n_6180),
.Y(n_6767)
);

BUFx6f_ASAP7_75t_L g6768 ( 
.A(n_6493),
.Y(n_6768)
);

BUFx12f_ASAP7_75t_L g6769 ( 
.A(n_6506),
.Y(n_6769)
);

CKINVDCx5p33_ASAP7_75t_R g6770 ( 
.A(n_6157),
.Y(n_6770)
);

INVx1_ASAP7_75t_L g6771 ( 
.A(n_6181),
.Y(n_6771)
);

CKINVDCx8_ASAP7_75t_R g6772 ( 
.A(n_6053),
.Y(n_6772)
);

CKINVDCx5p33_ASAP7_75t_R g6773 ( 
.A(n_6165),
.Y(n_6773)
);

INVxp33_ASAP7_75t_SL g6774 ( 
.A(n_6509),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_6182),
.Y(n_6775)
);

BUFx6f_ASAP7_75t_L g6776 ( 
.A(n_6166),
.Y(n_6776)
);

AND2x2_ASAP7_75t_L g6777 ( 
.A(n_6478),
.B(n_6102),
.Y(n_6777)
);

OA21x2_ASAP7_75t_L g6778 ( 
.A1(n_6437),
.A2(n_4750),
.B(n_4749),
.Y(n_6778)
);

BUFx6f_ASAP7_75t_L g6779 ( 
.A(n_6169),
.Y(n_6779)
);

OA21x2_ASAP7_75t_L g6780 ( 
.A1(n_6441),
.A2(n_4773),
.B(n_4753),
.Y(n_6780)
);

INVx2_ASAP7_75t_L g6781 ( 
.A(n_6492),
.Y(n_6781)
);

CKINVDCx5p33_ASAP7_75t_R g6782 ( 
.A(n_6172),
.Y(n_6782)
);

INVx3_ASAP7_75t_L g6783 ( 
.A(n_6183),
.Y(n_6783)
);

BUFx6f_ASAP7_75t_L g6784 ( 
.A(n_6177),
.Y(n_6784)
);

AND2x4_ASAP7_75t_L g6785 ( 
.A(n_6323),
.B(n_4902),
.Y(n_6785)
);

BUFx6f_ASAP7_75t_L g6786 ( 
.A(n_6191),
.Y(n_6786)
);

NAND2xp5_ASAP7_75t_L g6787 ( 
.A(n_6494),
.B(n_5345),
.Y(n_6787)
);

CKINVDCx5p33_ASAP7_75t_R g6788 ( 
.A(n_6193),
.Y(n_6788)
);

AND2x6_ASAP7_75t_L g6789 ( 
.A(n_6443),
.B(n_4929),
.Y(n_6789)
);

INVx2_ASAP7_75t_L g6790 ( 
.A(n_6495),
.Y(n_6790)
);

CKINVDCx20_ASAP7_75t_R g6791 ( 
.A(n_6039),
.Y(n_6791)
);

OAI22x1_ASAP7_75t_SL g6792 ( 
.A1(n_6404),
.A2(n_4648),
.B1(n_4654),
.B2(n_4638),
.Y(n_6792)
);

INVx2_ASAP7_75t_L g6793 ( 
.A(n_6496),
.Y(n_6793)
);

OAI22xp5_ASAP7_75t_SL g6794 ( 
.A1(n_6063),
.A2(n_4668),
.B1(n_4672),
.B2(n_4659),
.Y(n_6794)
);

CKINVDCx5p33_ASAP7_75t_R g6795 ( 
.A(n_6195),
.Y(n_6795)
);

BUFx3_ASAP7_75t_L g6796 ( 
.A(n_6418),
.Y(n_6796)
);

AND2x4_ASAP7_75t_L g6797 ( 
.A(n_6376),
.B(n_5071),
.Y(n_6797)
);

INVx2_ASAP7_75t_L g6798 ( 
.A(n_6497),
.Y(n_6798)
);

HB1xp67_ASAP7_75t_L g6799 ( 
.A(n_6213),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6184),
.Y(n_6800)
);

AND2x2_ASAP7_75t_L g6801 ( 
.A(n_6185),
.B(n_4761),
.Y(n_6801)
);

CKINVDCx20_ASAP7_75t_R g6802 ( 
.A(n_6068),
.Y(n_6802)
);

AND2x4_ASAP7_75t_L g6803 ( 
.A(n_6406),
.B(n_5172),
.Y(n_6803)
);

HB1xp67_ASAP7_75t_L g6804 ( 
.A(n_6218),
.Y(n_6804)
);

NAND2xp5_ASAP7_75t_SL g6805 ( 
.A(n_6289),
.B(n_4337),
.Y(n_6805)
);

BUFx6f_ASAP7_75t_L g6806 ( 
.A(n_6220),
.Y(n_6806)
);

INVx5_ASAP7_75t_L g6807 ( 
.A(n_6286),
.Y(n_6807)
);

CKINVDCx5p33_ASAP7_75t_R g6808 ( 
.A(n_6221),
.Y(n_6808)
);

OAI21x1_ASAP7_75t_L g6809 ( 
.A1(n_6186),
.A2(n_4382),
.B(n_4377),
.Y(n_6809)
);

BUFx3_ASAP7_75t_L g6810 ( 
.A(n_6429),
.Y(n_6810)
);

NOR2xp33_ASAP7_75t_L g6811 ( 
.A(n_6499),
.B(n_4299),
.Y(n_6811)
);

AND2x2_ASAP7_75t_L g6812 ( 
.A(n_6188),
.B(n_4785),
.Y(n_6812)
);

INVx2_ASAP7_75t_L g6813 ( 
.A(n_6500),
.Y(n_6813)
);

INVx2_ASAP7_75t_L g6814 ( 
.A(n_6501),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6503),
.Y(n_6815)
);

HB1xp67_ASAP7_75t_L g6816 ( 
.A(n_6224),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_6187),
.Y(n_6817)
);

BUFx6f_ASAP7_75t_L g6818 ( 
.A(n_6237),
.Y(n_6818)
);

INVx3_ASAP7_75t_L g6819 ( 
.A(n_6190),
.Y(n_6819)
);

AND2x4_ASAP7_75t_L g6820 ( 
.A(n_6444),
.B(n_5250),
.Y(n_6820)
);

AND2x4_ASAP7_75t_L g6821 ( 
.A(n_6432),
.B(n_5281),
.Y(n_6821)
);

BUFx6f_ASAP7_75t_L g6822 ( 
.A(n_6248),
.Y(n_6822)
);

OAI22xp5_ASAP7_75t_L g6823 ( 
.A1(n_6343),
.A2(n_5007),
.B1(n_5388),
.B2(n_4898),
.Y(n_6823)
);

INVx2_ASAP7_75t_L g6824 ( 
.A(n_6504),
.Y(n_6824)
);

OAI22xp5_ASAP7_75t_L g6825 ( 
.A1(n_6349),
.A2(n_5490),
.B1(n_4634),
.B2(n_4768),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_6194),
.Y(n_6826)
);

INVx1_ASAP7_75t_L g6827 ( 
.A(n_6196),
.Y(n_6827)
);

INVx3_ASAP7_75t_L g6828 ( 
.A(n_6198),
.Y(n_6828)
);

AND2x4_ASAP7_75t_L g6829 ( 
.A(n_6436),
.B(n_5299),
.Y(n_6829)
);

BUFx2_ASAP7_75t_L g6830 ( 
.A(n_6438),
.Y(n_6830)
);

BUFx3_ASAP7_75t_L g6831 ( 
.A(n_6440),
.Y(n_6831)
);

OAI21x1_ASAP7_75t_L g6832 ( 
.A1(n_6201),
.A2(n_4451),
.B(n_4432),
.Y(n_6832)
);

OA21x2_ASAP7_75t_L g6833 ( 
.A1(n_6202),
.A2(n_4779),
.B(n_4774),
.Y(n_6833)
);

BUFx3_ASAP7_75t_L g6834 ( 
.A(n_6450),
.Y(n_6834)
);

AOI22xp5_ASAP7_75t_L g6835 ( 
.A1(n_6445),
.A2(n_4201),
.B1(n_4287),
.B2(n_4178),
.Y(n_6835)
);

BUFx6f_ASAP7_75t_L g6836 ( 
.A(n_6251),
.Y(n_6836)
);

AND2x4_ASAP7_75t_L g6837 ( 
.A(n_6171),
.B(n_5368),
.Y(n_6837)
);

BUFx8_ASAP7_75t_SL g6838 ( 
.A(n_6076),
.Y(n_6838)
);

INVx2_ASAP7_75t_L g6839 ( 
.A(n_6508),
.Y(n_6839)
);

BUFx6f_ASAP7_75t_L g6840 ( 
.A(n_6263),
.Y(n_6840)
);

INVx3_ASAP7_75t_L g6841 ( 
.A(n_6204),
.Y(n_6841)
);

INVx5_ASAP7_75t_L g6842 ( 
.A(n_6351),
.Y(n_6842)
);

BUFx3_ASAP7_75t_L g6843 ( 
.A(n_6264),
.Y(n_6843)
);

BUFx3_ASAP7_75t_L g6844 ( 
.A(n_6265),
.Y(n_6844)
);

AOI22xp5_ASAP7_75t_L g6845 ( 
.A1(n_6267),
.A2(n_4391),
.B1(n_4423),
.B2(n_4352),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_6206),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6208),
.Y(n_6847)
);

OA21x2_ASAP7_75t_L g6848 ( 
.A1(n_6210),
.A2(n_4788),
.B(n_4780),
.Y(n_6848)
);

NAND2xp5_ASAP7_75t_SL g6849 ( 
.A(n_6272),
.B(n_6276),
.Y(n_6849)
);

BUFx6f_ASAP7_75t_L g6850 ( 
.A(n_6280),
.Y(n_6850)
);

INVx2_ASAP7_75t_L g6851 ( 
.A(n_6510),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6215),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6216),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6223),
.Y(n_6854)
);

BUFx2_ASAP7_75t_L g6855 ( 
.A(n_6200),
.Y(n_6855)
);

AOI22x1_ASAP7_75t_SL g6856 ( 
.A1(n_6088),
.A2(n_4698),
.B1(n_4702),
.B2(n_4681),
.Y(n_6856)
);

OAI22x1_ASAP7_75t_SL g6857 ( 
.A1(n_6097),
.A2(n_4748),
.B1(n_4814),
.B2(n_4742),
.Y(n_6857)
);

INVx1_ASAP7_75t_L g6858 ( 
.A(n_6226),
.Y(n_6858)
);

INVx2_ASAP7_75t_L g6859 ( 
.A(n_6227),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_6228),
.Y(n_6860)
);

INVx6_ASAP7_75t_L g6861 ( 
.A(n_6357),
.Y(n_6861)
);

INVx1_ASAP7_75t_L g6862 ( 
.A(n_6231),
.Y(n_6862)
);

BUFx2_ASAP7_75t_L g6863 ( 
.A(n_6211),
.Y(n_6863)
);

INVx2_ASAP7_75t_L g6864 ( 
.A(n_6232),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6233),
.Y(n_6865)
);

CKINVDCx6p67_ASAP7_75t_R g6866 ( 
.A(n_6137),
.Y(n_6866)
);

AOI22xp5_ASAP7_75t_L g6867 ( 
.A1(n_6292),
.A2(n_4540),
.B1(n_4555),
.B2(n_4470),
.Y(n_6867)
);

AND2x2_ASAP7_75t_SL g6868 ( 
.A(n_6038),
.B(n_4469),
.Y(n_6868)
);

BUFx6f_ASAP7_75t_L g6869 ( 
.A(n_6297),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6234),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6235),
.Y(n_6871)
);

HB1xp67_ASAP7_75t_L g6872 ( 
.A(n_6298),
.Y(n_6872)
);

INVx5_ASAP7_75t_L g6873 ( 
.A(n_6001),
.Y(n_6873)
);

AOI22xp5_ASAP7_75t_SL g6874 ( 
.A1(n_6099),
.A2(n_4852),
.B1(n_4853),
.B2(n_4831),
.Y(n_6874)
);

BUFx6f_ASAP7_75t_L g6875 ( 
.A(n_6310),
.Y(n_6875)
);

NAND2xp5_ASAP7_75t_L g6876 ( 
.A(n_6294),
.B(n_5363),
.Y(n_6876)
);

AND2x4_ASAP7_75t_L g6877 ( 
.A(n_6214),
.B(n_5457),
.Y(n_6877)
);

NOR2x1_ASAP7_75t_L g6878 ( 
.A(n_6240),
.B(n_5464),
.Y(n_6878)
);

INVx6_ASAP7_75t_L g6879 ( 
.A(n_6083),
.Y(n_6879)
);

NAND2xp5_ASAP7_75t_L g6880 ( 
.A(n_6244),
.B(n_5363),
.Y(n_6880)
);

BUFx12f_ASAP7_75t_L g6881 ( 
.A(n_6318),
.Y(n_6881)
);

BUFx2_ASAP7_75t_L g6882 ( 
.A(n_6225),
.Y(n_6882)
);

NAND2xp5_ASAP7_75t_L g6883 ( 
.A(n_6245),
.B(n_5363),
.Y(n_6883)
);

OAI21x1_ASAP7_75t_L g6884 ( 
.A1(n_6246),
.A2(n_6253),
.B(n_6252),
.Y(n_6884)
);

INVx3_ASAP7_75t_L g6885 ( 
.A(n_6256),
.Y(n_6885)
);

INVx2_ASAP7_75t_SL g6886 ( 
.A(n_6319),
.Y(n_6886)
);

OAI22xp5_ASAP7_75t_L g6887 ( 
.A1(n_6321),
.A2(n_4956),
.B1(n_5056),
.B2(n_4613),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_6257),
.Y(n_6888)
);

BUFx6f_ASAP7_75t_L g6889 ( 
.A(n_6326),
.Y(n_6889)
);

INVx2_ASAP7_75t_L g6890 ( 
.A(n_6258),
.Y(n_6890)
);

AND2x2_ASAP7_75t_L g6891 ( 
.A(n_6329),
.B(n_4785),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6266),
.Y(n_6892)
);

INVxp33_ASAP7_75t_SL g6893 ( 
.A(n_6332),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6269),
.Y(n_6894)
);

HB1xp67_ASAP7_75t_L g6895 ( 
.A(n_6334),
.Y(n_6895)
);

INVx1_ASAP7_75t_L g6896 ( 
.A(n_6270),
.Y(n_6896)
);

INVx2_ASAP7_75t_SL g6897 ( 
.A(n_6337),
.Y(n_6897)
);

AND2x4_ASAP7_75t_L g6898 ( 
.A(n_6229),
.B(n_4392),
.Y(n_6898)
);

INVx2_ASAP7_75t_L g6899 ( 
.A(n_6271),
.Y(n_6899)
);

AND2x4_ASAP7_75t_L g6900 ( 
.A(n_6241),
.B(n_4424),
.Y(n_6900)
);

INVx3_ASAP7_75t_L g6901 ( 
.A(n_6273),
.Y(n_6901)
);

INVx3_ASAP7_75t_L g6902 ( 
.A(n_6274),
.Y(n_6902)
);

INVx3_ASAP7_75t_L g6903 ( 
.A(n_6275),
.Y(n_6903)
);

OAI21x1_ASAP7_75t_L g6904 ( 
.A1(n_6279),
.A2(n_4535),
.B(n_4478),
.Y(n_6904)
);

BUFx3_ASAP7_75t_L g6905 ( 
.A(n_6339),
.Y(n_6905)
);

HB1xp67_ASAP7_75t_L g6906 ( 
.A(n_6342),
.Y(n_6906)
);

OAI22xp5_ASAP7_75t_L g6907 ( 
.A1(n_6354),
.A2(n_5184),
.B1(n_4342),
.B2(n_4345),
.Y(n_6907)
);

INVx3_ASAP7_75t_L g6908 ( 
.A(n_6285),
.Y(n_6908)
);

AND2x4_ASAP7_75t_L g6909 ( 
.A(n_6108),
.B(n_4495),
.Y(n_6909)
);

BUFx12f_ASAP7_75t_L g6910 ( 
.A(n_6358),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6287),
.Y(n_6911)
);

BUFx12f_ASAP7_75t_L g6912 ( 
.A(n_6365),
.Y(n_6912)
);

CKINVDCx6p67_ASAP7_75t_R g6913 ( 
.A(n_6163),
.Y(n_6913)
);

INVx5_ASAP7_75t_L g6914 ( 
.A(n_6167),
.Y(n_6914)
);

INVx3_ASAP7_75t_L g6915 ( 
.A(n_6288),
.Y(n_6915)
);

BUFx6f_ASAP7_75t_L g6916 ( 
.A(n_6367),
.Y(n_6916)
);

AOI22xp5_ASAP7_75t_L g6917 ( 
.A1(n_6369),
.A2(n_4614),
.B1(n_4637),
.B2(n_4593),
.Y(n_6917)
);

INVx2_ASAP7_75t_L g6918 ( 
.A(n_6290),
.Y(n_6918)
);

HB1xp67_ASAP7_75t_L g6919 ( 
.A(n_6386),
.Y(n_6919)
);

INVx1_ASAP7_75t_L g6920 ( 
.A(n_6296),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6302),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6303),
.Y(n_6922)
);

BUFx6f_ASAP7_75t_L g6923 ( 
.A(n_6398),
.Y(n_6923)
);

HB1xp67_ASAP7_75t_L g6924 ( 
.A(n_6415),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_6305),
.Y(n_6925)
);

INVx1_ASAP7_75t_L g6926 ( 
.A(n_6306),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_6307),
.Y(n_6927)
);

INVx2_ASAP7_75t_L g6928 ( 
.A(n_6308),
.Y(n_6928)
);

CKINVDCx5p33_ASAP7_75t_R g6929 ( 
.A(n_6424),
.Y(n_6929)
);

INVx4_ASAP7_75t_L g6930 ( 
.A(n_6430),
.Y(n_6930)
);

NAND2xp5_ASAP7_75t_L g6931 ( 
.A(n_6309),
.B(n_5497),
.Y(n_6931)
);

OAI21x1_ASAP7_75t_L g6932 ( 
.A1(n_6312),
.A2(n_4570),
.B(n_4558),
.Y(n_6932)
);

INVx2_ASAP7_75t_L g6933 ( 
.A(n_6313),
.Y(n_6933)
);

HB1xp67_ASAP7_75t_L g6934 ( 
.A(n_6431),
.Y(n_6934)
);

INVx2_ASAP7_75t_L g6935 ( 
.A(n_6314),
.Y(n_6935)
);

INVx3_ASAP7_75t_L g6936 ( 
.A(n_6315),
.Y(n_6936)
);

OAI22x1_ASAP7_75t_R g6937 ( 
.A1(n_6129),
.A2(n_4877),
.B1(n_4881),
.B2(n_4870),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6320),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6322),
.Y(n_6939)
);

INVx2_ASAP7_75t_L g6940 ( 
.A(n_6328),
.Y(n_6940)
);

AND2x4_ASAP7_75t_SL g6941 ( 
.A(n_6168),
.B(n_4797),
.Y(n_6941)
);

BUFx6f_ASAP7_75t_L g6942 ( 
.A(n_6433),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6333),
.Y(n_6943)
);

BUFx6f_ASAP7_75t_L g6944 ( 
.A(n_6435),
.Y(n_6944)
);

INVx2_ASAP7_75t_L g6945 ( 
.A(n_6336),
.Y(n_6945)
);

BUFx8_ASAP7_75t_L g6946 ( 
.A(n_6468),
.Y(n_6946)
);

AND2x4_ASAP7_75t_L g6947 ( 
.A(n_6469),
.B(n_6485),
.Y(n_6947)
);

BUFx6f_ASAP7_75t_L g6948 ( 
.A(n_6439),
.Y(n_6948)
);

BUFx6f_ASAP7_75t_L g6949 ( 
.A(n_6442),
.Y(n_6949)
);

BUFx3_ASAP7_75t_L g6950 ( 
.A(n_6449),
.Y(n_6950)
);

INVx6_ASAP7_75t_L g6951 ( 
.A(n_6486),
.Y(n_6951)
);

INVx1_ASAP7_75t_L g6952 ( 
.A(n_6338),
.Y(n_6952)
);

INVx6_ASAP7_75t_L g6953 ( 
.A(n_6488),
.Y(n_6953)
);

AOI22xp5_ASAP7_75t_SL g6954 ( 
.A1(n_6491),
.A2(n_4931),
.B1(n_4933),
.B2(n_4911),
.Y(n_6954)
);

BUFx6f_ASAP7_75t_L g6955 ( 
.A(n_6457),
.Y(n_6955)
);

BUFx6f_ASAP7_75t_L g6956 ( 
.A(n_6340),
.Y(n_6956)
);

NAND2xp5_ASAP7_75t_L g6957 ( 
.A(n_6341),
.B(n_5497),
.Y(n_6957)
);

OA21x2_ASAP7_75t_L g6958 ( 
.A1(n_6347),
.A2(n_4793),
.B(n_4792),
.Y(n_6958)
);

INVx4_ASAP7_75t_L g6959 ( 
.A(n_6348),
.Y(n_6959)
);

AND2x6_ASAP7_75t_L g6960 ( 
.A(n_6350),
.B(n_4641),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6352),
.Y(n_6961)
);

OA21x2_ASAP7_75t_L g6962 ( 
.A1(n_6353),
.A2(n_4795),
.B(n_4794),
.Y(n_6962)
);

INVx3_ASAP7_75t_L g6963 ( 
.A(n_6356),
.Y(n_6963)
);

HB1xp67_ASAP7_75t_L g6964 ( 
.A(n_6498),
.Y(n_6964)
);

INVx2_ASAP7_75t_L g6965 ( 
.A(n_6359),
.Y(n_6965)
);

BUFx8_ASAP7_75t_L g6966 ( 
.A(n_6502),
.Y(n_6966)
);

BUFx6f_ASAP7_75t_L g6967 ( 
.A(n_6360),
.Y(n_6967)
);

INVx2_ASAP7_75t_L g6968 ( 
.A(n_6361),
.Y(n_6968)
);

INVxp67_ASAP7_75t_L g6969 ( 
.A(n_6101),
.Y(n_6969)
);

INVx2_ASAP7_75t_L g6970 ( 
.A(n_6364),
.Y(n_6970)
);

AND2x4_ASAP7_75t_L g6971 ( 
.A(n_6511),
.B(n_4525),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_6366),
.Y(n_6972)
);

BUFx6f_ASAP7_75t_L g6973 ( 
.A(n_6368),
.Y(n_6973)
);

OAI22xp5_ASAP7_75t_SL g6974 ( 
.A1(n_6164),
.A2(n_4941),
.B1(n_4966),
.B2(n_4937),
.Y(n_6974)
);

AND2x4_ASAP7_75t_L g6975 ( 
.A(n_6370),
.B(n_4588),
.Y(n_6975)
);

INVx1_ASAP7_75t_L g6976 ( 
.A(n_6372),
.Y(n_6976)
);

INVx3_ASAP7_75t_L g6977 ( 
.A(n_6373),
.Y(n_6977)
);

AND2x6_ASAP7_75t_L g6978 ( 
.A(n_6374),
.B(n_4663),
.Y(n_6978)
);

BUFx3_ASAP7_75t_L g6979 ( 
.A(n_6067),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_6377),
.Y(n_6980)
);

INVx1_ASAP7_75t_L g6981 ( 
.A(n_6378),
.Y(n_6981)
);

INVx2_ASAP7_75t_L g6982 ( 
.A(n_6379),
.Y(n_6982)
);

INVx2_ASAP7_75t_L g6983 ( 
.A(n_6381),
.Y(n_6983)
);

NOR2x1_ASAP7_75t_L g6984 ( 
.A(n_6382),
.B(n_4796),
.Y(n_6984)
);

OAI22xp5_ASAP7_75t_SL g6985 ( 
.A1(n_6034),
.A2(n_5020),
.B1(n_5037),
.B2(n_4985),
.Y(n_6985)
);

CKINVDCx16_ASAP7_75t_R g6986 ( 
.A(n_6142),
.Y(n_6986)
);

INVx2_ASAP7_75t_L g6987 ( 
.A(n_6383),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_6385),
.B(n_5497),
.Y(n_6988)
);

HB1xp67_ASAP7_75t_L g6989 ( 
.A(n_6159),
.Y(n_6989)
);

INVx5_ASAP7_75t_L g6990 ( 
.A(n_6207),
.Y(n_6990)
);

INVx2_ASAP7_75t_L g6991 ( 
.A(n_6388),
.Y(n_6991)
);

AND2x4_ASAP7_75t_L g6992 ( 
.A(n_6111),
.B(n_4612),
.Y(n_6992)
);

OA21x2_ASAP7_75t_L g6993 ( 
.A1(n_6355),
.A2(n_4803),
.B(n_4800),
.Y(n_6993)
);

NAND2xp5_ASAP7_75t_L g6994 ( 
.A(n_6375),
.B(n_4617),
.Y(n_6994)
);

INVx2_ASAP7_75t_L g6995 ( 
.A(n_6426),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6113),
.Y(n_6996)
);

CKINVDCx6p67_ASAP7_75t_R g6997 ( 
.A(n_6230),
.Y(n_6997)
);

INVx3_ASAP7_75t_L g6998 ( 
.A(n_6461),
.Y(n_6998)
);

BUFx6f_ASAP7_75t_L g6999 ( 
.A(n_6147),
.Y(n_6999)
);

NAND2xp5_ASAP7_75t_L g7000 ( 
.A(n_6150),
.B(n_4917),
.Y(n_7000)
);

INVx3_ASAP7_75t_L g7001 ( 
.A(n_6151),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6161),
.B(n_4797),
.Y(n_7002)
);

INVx2_ASAP7_75t_L g7003 ( 
.A(n_6173),
.Y(n_7003)
);

AOI22xp5_ASAP7_75t_L g7004 ( 
.A1(n_6197),
.A2(n_4723),
.B1(n_4799),
.B2(n_4674),
.Y(n_7004)
);

INVx2_ASAP7_75t_L g7005 ( 
.A(n_6219),
.Y(n_7005)
);

BUFx2_ASAP7_75t_L g7006 ( 
.A(n_6236),
.Y(n_7006)
);

BUFx6f_ASAP7_75t_L g7007 ( 
.A(n_6255),
.Y(n_7007)
);

OAI22xp5_ASAP7_75t_L g7008 ( 
.A1(n_6262),
.A2(n_4346),
.B1(n_4348),
.B2(n_4340),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6268),
.Y(n_7009)
);

AND2x2_ASAP7_75t_L g7010 ( 
.A(n_6277),
.B(n_4837),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6009),
.Y(n_7011)
);

BUFx3_ASAP7_75t_L g7012 ( 
.A(n_6022),
.Y(n_7012)
);

INVx2_ASAP7_75t_L g7013 ( 
.A(n_6301),
.Y(n_7013)
);

BUFx6f_ASAP7_75t_L g7014 ( 
.A(n_6022),
.Y(n_7014)
);

INVx2_ASAP7_75t_L g7015 ( 
.A(n_6301),
.Y(n_7015)
);

INVx2_ASAP7_75t_L g7016 ( 
.A(n_6301),
.Y(n_7016)
);

OA21x2_ASAP7_75t_L g7017 ( 
.A1(n_6410),
.A2(n_4808),
.B(n_4804),
.Y(n_7017)
);

BUFx6f_ASAP7_75t_L g7018 ( 
.A(n_6022),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6009),
.Y(n_7019)
);

INVx2_ASAP7_75t_L g7020 ( 
.A(n_6301),
.Y(n_7020)
);

AND2x2_ASAP7_75t_SL g7021 ( 
.A(n_6027),
.B(n_4575),
.Y(n_7021)
);

INVx2_ASAP7_75t_L g7022 ( 
.A(n_6301),
.Y(n_7022)
);

INVx2_ASAP7_75t_L g7023 ( 
.A(n_6301),
.Y(n_7023)
);

NAND2xp5_ASAP7_75t_L g7024 ( 
.A(n_6409),
.B(n_4924),
.Y(n_7024)
);

INVx2_ASAP7_75t_L g7025 ( 
.A(n_6301),
.Y(n_7025)
);

INVx3_ASAP7_75t_L g7026 ( 
.A(n_6022),
.Y(n_7026)
);

OAI22xp5_ASAP7_75t_L g7027 ( 
.A1(n_6295),
.A2(n_4354),
.B1(n_4355),
.B2(n_4351),
.Y(n_7027)
);

BUFx6f_ASAP7_75t_L g7028 ( 
.A(n_6022),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6009),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6009),
.Y(n_7030)
);

NAND2xp5_ASAP7_75t_L g7031 ( 
.A(n_6409),
.B(n_4936),
.Y(n_7031)
);

NAND2xp5_ASAP7_75t_L g7032 ( 
.A(n_6409),
.B(n_4990),
.Y(n_7032)
);

AND2x2_ASAP7_75t_SL g7033 ( 
.A(n_6027),
.B(n_4598),
.Y(n_7033)
);

INVx2_ASAP7_75t_L g7034 ( 
.A(n_6301),
.Y(n_7034)
);

INVx3_ASAP7_75t_L g7035 ( 
.A(n_6022),
.Y(n_7035)
);

AND2x4_ASAP7_75t_L g7036 ( 
.A(n_6460),
.B(n_5043),
.Y(n_7036)
);

AOI22x1_ASAP7_75t_SL g7037 ( 
.A1(n_6008),
.A2(n_5053),
.B1(n_5058),
.B2(n_5039),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6009),
.Y(n_7038)
);

AND2x4_ASAP7_75t_L g7039 ( 
.A(n_6460),
.B(n_5093),
.Y(n_7039)
);

BUFx6f_ASAP7_75t_L g7040 ( 
.A(n_6022),
.Y(n_7040)
);

BUFx8_ASAP7_75t_L g7041 ( 
.A(n_6042),
.Y(n_7041)
);

BUFx6f_ASAP7_75t_L g7042 ( 
.A(n_6022),
.Y(n_7042)
);

AND2x2_ASAP7_75t_L g7043 ( 
.A(n_6140),
.B(n_4837),
.Y(n_7043)
);

AND2x4_ASAP7_75t_L g7044 ( 
.A(n_6460),
.B(n_5116),
.Y(n_7044)
);

INVx1_ASAP7_75t_L g7045 ( 
.A(n_6009),
.Y(n_7045)
);

INVx5_ASAP7_75t_L g7046 ( 
.A(n_6095),
.Y(n_7046)
);

BUFx6f_ASAP7_75t_L g7047 ( 
.A(n_6022),
.Y(n_7047)
);

NAND2xp5_ASAP7_75t_L g7048 ( 
.A(n_6409),
.B(n_5232),
.Y(n_7048)
);

AOI22xp5_ASAP7_75t_L g7049 ( 
.A1(n_6278),
.A2(n_4857),
.B1(n_4872),
.B2(n_4843),
.Y(n_7049)
);

HB1xp67_ASAP7_75t_L g7050 ( 
.A(n_6011),
.Y(n_7050)
);

INVx4_ASAP7_75t_L g7051 ( 
.A(n_6079),
.Y(n_7051)
);

OAI22xp5_ASAP7_75t_L g7052 ( 
.A1(n_6295),
.A2(n_4358),
.B1(n_4362),
.B2(n_4357),
.Y(n_7052)
);

CKINVDCx20_ASAP7_75t_R g7053 ( 
.A(n_6008),
.Y(n_7053)
);

AND2x4_ASAP7_75t_L g7054 ( 
.A(n_6460),
.B(n_5460),
.Y(n_7054)
);

BUFx3_ASAP7_75t_L g7055 ( 
.A(n_6022),
.Y(n_7055)
);

BUFx2_ASAP7_75t_L g7056 ( 
.A(n_6462),
.Y(n_7056)
);

BUFx2_ASAP7_75t_L g7057 ( 
.A(n_6462),
.Y(n_7057)
);

AOI22x1_ASAP7_75t_SL g7058 ( 
.A1(n_6008),
.A2(n_5088),
.B1(n_5143),
.B2(n_5084),
.Y(n_7058)
);

NOR2xp33_ASAP7_75t_L g7059 ( 
.A(n_6409),
.B(n_5462),
.Y(n_7059)
);

AOI22xp5_ASAP7_75t_L g7060 ( 
.A1(n_6278),
.A2(n_4904),
.B1(n_4950),
.B2(n_4887),
.Y(n_7060)
);

INVx2_ASAP7_75t_L g7061 ( 
.A(n_6301),
.Y(n_7061)
);

AND2x2_ASAP7_75t_L g7062 ( 
.A(n_6140),
.B(n_4885),
.Y(n_7062)
);

AND2x4_ASAP7_75t_L g7063 ( 
.A(n_6460),
.B(n_5481),
.Y(n_7063)
);

INVx1_ASAP7_75t_SL g7064 ( 
.A(n_6466),
.Y(n_7064)
);

BUFx6f_ASAP7_75t_L g7065 ( 
.A(n_6022),
.Y(n_7065)
);

AND2x2_ASAP7_75t_L g7066 ( 
.A(n_6140),
.B(n_4885),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6009),
.Y(n_7067)
);

INVx2_ASAP7_75t_L g7068 ( 
.A(n_6301),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6301),
.Y(n_7069)
);

BUFx6f_ASAP7_75t_L g7070 ( 
.A(n_6022),
.Y(n_7070)
);

INVx2_ASAP7_75t_L g7071 ( 
.A(n_6301),
.Y(n_7071)
);

INVx1_ASAP7_75t_L g7072 ( 
.A(n_6009),
.Y(n_7072)
);

INVx2_ASAP7_75t_L g7073 ( 
.A(n_6301),
.Y(n_7073)
);

AND2x4_ASAP7_75t_L g7074 ( 
.A(n_6460),
.B(n_5547),
.Y(n_7074)
);

HB1xp67_ASAP7_75t_L g7075 ( 
.A(n_6011),
.Y(n_7075)
);

XNOR2xp5_ASAP7_75t_L g7076 ( 
.A(n_6008),
.B(n_5150),
.Y(n_7076)
);

AOI22xp5_ASAP7_75t_L g7077 ( 
.A1(n_6278),
.A2(n_5026),
.B1(n_5047),
.B2(n_5019),
.Y(n_7077)
);

BUFx6f_ASAP7_75t_L g7078 ( 
.A(n_6022),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6009),
.Y(n_7079)
);

BUFx6f_ASAP7_75t_L g7080 ( 
.A(n_6022),
.Y(n_7080)
);

NOR2xp33_ASAP7_75t_L g7081 ( 
.A(n_6409),
.B(n_4365),
.Y(n_7081)
);

OAI22x1_ASAP7_75t_R g7082 ( 
.A1(n_6250),
.A2(n_5165),
.B1(n_5170),
.B2(n_5158),
.Y(n_7082)
);

INVx3_ASAP7_75t_L g7083 ( 
.A(n_6022),
.Y(n_7083)
);

INVx2_ASAP7_75t_L g7084 ( 
.A(n_6301),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6009),
.Y(n_7085)
);

BUFx6f_ASAP7_75t_L g7086 ( 
.A(n_6022),
.Y(n_7086)
);

INVx4_ASAP7_75t_L g7087 ( 
.A(n_6079),
.Y(n_7087)
);

INVx2_ASAP7_75t_L g7088 ( 
.A(n_6301),
.Y(n_7088)
);

AND2x4_ASAP7_75t_L g7089 ( 
.A(n_6460),
.B(n_5199),
.Y(n_7089)
);

BUFx2_ASAP7_75t_L g7090 ( 
.A(n_6462),
.Y(n_7090)
);

AND2x6_ASAP7_75t_L g7091 ( 
.A(n_6392),
.B(n_5060),
.Y(n_7091)
);

NAND2xp5_ASAP7_75t_L g7092 ( 
.A(n_6550),
.B(n_4368),
.Y(n_7092)
);

HB1xp67_ASAP7_75t_L g7093 ( 
.A(n_6517),
.Y(n_7093)
);

CKINVDCx5p33_ASAP7_75t_R g7094 ( 
.A(n_6516),
.Y(n_7094)
);

INVx2_ASAP7_75t_L g7095 ( 
.A(n_6611),
.Y(n_7095)
);

BUFx2_ASAP7_75t_L g7096 ( 
.A(n_6747),
.Y(n_7096)
);

BUFx6f_ASAP7_75t_L g7097 ( 
.A(n_6633),
.Y(n_7097)
);

CKINVDCx20_ASAP7_75t_R g7098 ( 
.A(n_6749),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6884),
.Y(n_7099)
);

INVx1_ASAP7_75t_L g7100 ( 
.A(n_6708),
.Y(n_7100)
);

HB1xp67_ASAP7_75t_L g7101 ( 
.A(n_7050),
.Y(n_7101)
);

BUFx6f_ASAP7_75t_L g7102 ( 
.A(n_6634),
.Y(n_7102)
);

CKINVDCx5p33_ASAP7_75t_R g7103 ( 
.A(n_6548),
.Y(n_7103)
);

BUFx2_ASAP7_75t_L g7104 ( 
.A(n_6791),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6712),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6729),
.Y(n_7106)
);

INVx1_ASAP7_75t_L g7107 ( 
.A(n_6733),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6742),
.Y(n_7108)
);

OA21x2_ASAP7_75t_L g7109 ( 
.A1(n_6613),
.A2(n_4812),
.B(n_4810),
.Y(n_7109)
);

INVx2_ASAP7_75t_L g7110 ( 
.A(n_6536),
.Y(n_7110)
);

NOR2xp33_ASAP7_75t_R g7111 ( 
.A(n_6586),
.B(n_5206),
.Y(n_7111)
);

AND2x2_ASAP7_75t_L g7112 ( 
.A(n_7064),
.B(n_5260),
.Y(n_7112)
);

CKINVDCx5p33_ASAP7_75t_R g7113 ( 
.A(n_6685),
.Y(n_7113)
);

NOR2xp33_ASAP7_75t_L g7114 ( 
.A(n_6619),
.B(n_5086),
.Y(n_7114)
);

CKINVDCx5p33_ASAP7_75t_R g7115 ( 
.A(n_6686),
.Y(n_7115)
);

CKINVDCx20_ASAP7_75t_R g7116 ( 
.A(n_6802),
.Y(n_7116)
);

BUFx6f_ASAP7_75t_L g7117 ( 
.A(n_6515),
.Y(n_7117)
);

INVx1_ASAP7_75t_L g7118 ( 
.A(n_6746),
.Y(n_7118)
);

CKINVDCx5p33_ASAP7_75t_R g7119 ( 
.A(n_6770),
.Y(n_7119)
);

CKINVDCx5p33_ASAP7_75t_R g7120 ( 
.A(n_6773),
.Y(n_7120)
);

INVx1_ASAP7_75t_L g7121 ( 
.A(n_6748),
.Y(n_7121)
);

INVx2_ASAP7_75t_L g7122 ( 
.A(n_6537),
.Y(n_7122)
);

INVx3_ASAP7_75t_L g7123 ( 
.A(n_6542),
.Y(n_7123)
);

INVx3_ASAP7_75t_L g7124 ( 
.A(n_6535),
.Y(n_7124)
);

BUFx2_ASAP7_75t_L g7125 ( 
.A(n_7053),
.Y(n_7125)
);

CKINVDCx5p33_ASAP7_75t_R g7126 ( 
.A(n_6782),
.Y(n_7126)
);

CKINVDCx5p33_ASAP7_75t_R g7127 ( 
.A(n_6788),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_6750),
.Y(n_7128)
);

CKINVDCx5p33_ASAP7_75t_R g7129 ( 
.A(n_6795),
.Y(n_7129)
);

HB1xp67_ASAP7_75t_L g7130 ( 
.A(n_7075),
.Y(n_7130)
);

INVx2_ASAP7_75t_L g7131 ( 
.A(n_6522),
.Y(n_7131)
);

CKINVDCx5p33_ASAP7_75t_R g7132 ( 
.A(n_6808),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_6759),
.Y(n_7133)
);

INVx2_ASAP7_75t_L g7134 ( 
.A(n_6528),
.Y(n_7134)
);

NAND2xp5_ASAP7_75t_L g7135 ( 
.A(n_6592),
.B(n_4371),
.Y(n_7135)
);

BUFx6f_ASAP7_75t_L g7136 ( 
.A(n_7014),
.Y(n_7136)
);

BUFx2_ASAP7_75t_L g7137 ( 
.A(n_6547),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_6533),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_6765),
.Y(n_7139)
);

OAI21x1_ASAP7_75t_L g7140 ( 
.A1(n_6681),
.A2(n_4604),
.B(n_4600),
.Y(n_7140)
);

CKINVDCx5p33_ASAP7_75t_R g7141 ( 
.A(n_6929),
.Y(n_7141)
);

NAND2xp5_ASAP7_75t_SL g7142 ( 
.A(n_6754),
.B(n_4373),
.Y(n_7142)
);

NOR2xp33_ASAP7_75t_R g7143 ( 
.A(n_6986),
.B(n_5283),
.Y(n_7143)
);

INVx1_ASAP7_75t_L g7144 ( 
.A(n_6766),
.Y(n_7144)
);

INVx2_ASAP7_75t_L g7145 ( 
.A(n_6539),
.Y(n_7145)
);

INVx2_ASAP7_75t_L g7146 ( 
.A(n_6552),
.Y(n_7146)
);

HB1xp67_ASAP7_75t_L g7147 ( 
.A(n_6581),
.Y(n_7147)
);

INVx2_ASAP7_75t_L g7148 ( 
.A(n_6554),
.Y(n_7148)
);

NAND2xp5_ASAP7_75t_SL g7149 ( 
.A(n_6544),
.B(n_4375),
.Y(n_7149)
);

INVx1_ASAP7_75t_L g7150 ( 
.A(n_6781),
.Y(n_7150)
);

INVx3_ASAP7_75t_L g7151 ( 
.A(n_6545),
.Y(n_7151)
);

NOR2xp33_ASAP7_75t_L g7152 ( 
.A(n_6893),
.B(n_5120),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6790),
.Y(n_7153)
);

INVx1_ASAP7_75t_L g7154 ( 
.A(n_6793),
.Y(n_7154)
);

INVx3_ASAP7_75t_L g7155 ( 
.A(n_6558),
.Y(n_7155)
);

CKINVDCx5p33_ASAP7_75t_R g7156 ( 
.A(n_6728),
.Y(n_7156)
);

AND2x2_ASAP7_75t_L g7157 ( 
.A(n_6596),
.B(n_5288),
.Y(n_7157)
);

CKINVDCx5p33_ASAP7_75t_R g7158 ( 
.A(n_6774),
.Y(n_7158)
);

CKINVDCx11_ASAP7_75t_R g7159 ( 
.A(n_6655),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_6798),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_6813),
.Y(n_7161)
);

CKINVDCx5p33_ASAP7_75t_R g7162 ( 
.A(n_6838),
.Y(n_7162)
);

HB1xp67_ASAP7_75t_L g7163 ( 
.A(n_6947),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_6814),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_6815),
.Y(n_7165)
);

CKINVDCx5p33_ASAP7_75t_R g7166 ( 
.A(n_6881),
.Y(n_7166)
);

NOR2xp33_ASAP7_75t_L g7167 ( 
.A(n_6588),
.B(n_5146),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6824),
.Y(n_7168)
);

CKINVDCx20_ASAP7_75t_R g7169 ( 
.A(n_6997),
.Y(n_7169)
);

CKINVDCx5p33_ASAP7_75t_R g7170 ( 
.A(n_6910),
.Y(n_7170)
);

CKINVDCx5p33_ASAP7_75t_R g7171 ( 
.A(n_6912),
.Y(n_7171)
);

CKINVDCx5p33_ASAP7_75t_R g7172 ( 
.A(n_6716),
.Y(n_7172)
);

BUFx2_ASAP7_75t_L g7173 ( 
.A(n_7056),
.Y(n_7173)
);

INVx2_ASAP7_75t_L g7174 ( 
.A(n_6559),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6839),
.Y(n_7175)
);

CKINVDCx20_ASAP7_75t_R g7176 ( 
.A(n_6683),
.Y(n_7176)
);

CKINVDCx20_ASAP7_75t_R g7177 ( 
.A(n_6946),
.Y(n_7177)
);

INVx1_ASAP7_75t_SL g7178 ( 
.A(n_6951),
.Y(n_7178)
);

CKINVDCx5p33_ASAP7_75t_R g7179 ( 
.A(n_6727),
.Y(n_7179)
);

HB1xp67_ASAP7_75t_L g7180 ( 
.A(n_6964),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6851),
.Y(n_7181)
);

INVx1_ASAP7_75t_L g7182 ( 
.A(n_6527),
.Y(n_7182)
);

NOR2xp33_ASAP7_75t_R g7183 ( 
.A(n_6772),
.B(n_5293),
.Y(n_7183)
);

CKINVDCx20_ASAP7_75t_R g7184 ( 
.A(n_6966),
.Y(n_7184)
);

CKINVDCx5p33_ASAP7_75t_R g7185 ( 
.A(n_6730),
.Y(n_7185)
);

AND2x2_ASAP7_75t_L g7186 ( 
.A(n_7057),
.B(n_5309),
.Y(n_7186)
);

INVx2_ASAP7_75t_L g7187 ( 
.A(n_6560),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_SL g7188 ( 
.A(n_6566),
.B(n_4378),
.Y(n_7188)
);

CKINVDCx20_ASAP7_75t_R g7189 ( 
.A(n_6866),
.Y(n_7189)
);

BUFx6f_ASAP7_75t_L g7190 ( 
.A(n_7018),
.Y(n_7190)
);

BUFx6f_ASAP7_75t_L g7191 ( 
.A(n_7028),
.Y(n_7191)
);

CKINVDCx20_ASAP7_75t_R g7192 ( 
.A(n_6913),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_6530),
.Y(n_7193)
);

CKINVDCx5p33_ASAP7_75t_R g7194 ( 
.A(n_6758),
.Y(n_7194)
);

INVx1_ASAP7_75t_SL g7195 ( 
.A(n_6953),
.Y(n_7195)
);

INVx2_ASAP7_75t_L g7196 ( 
.A(n_6564),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_6531),
.Y(n_7197)
);

HB1xp67_ASAP7_75t_L g7198 ( 
.A(n_6665),
.Y(n_7198)
);

CKINVDCx5p33_ASAP7_75t_R g7199 ( 
.A(n_6769),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_6532),
.Y(n_7200)
);

INVx2_ASAP7_75t_L g7201 ( 
.A(n_6571),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6540),
.Y(n_7202)
);

NOR2xp33_ASAP7_75t_R g7203 ( 
.A(n_6703),
.B(n_5322),
.Y(n_7203)
);

BUFx6f_ASAP7_75t_L g7204 ( 
.A(n_7040),
.Y(n_7204)
);

BUFx3_ASAP7_75t_L g7205 ( 
.A(n_6556),
.Y(n_7205)
);

INVx1_ASAP7_75t_L g7206 ( 
.A(n_6553),
.Y(n_7206)
);

NOR2xp33_ASAP7_75t_R g7207 ( 
.A(n_6565),
.B(n_5337),
.Y(n_7207)
);

CKINVDCx16_ASAP7_75t_R g7208 ( 
.A(n_6605),
.Y(n_7208)
);

BUFx6f_ASAP7_75t_L g7209 ( 
.A(n_7042),
.Y(n_7209)
);

INVx2_ASAP7_75t_L g7210 ( 
.A(n_6578),
.Y(n_7210)
);

BUFx6f_ASAP7_75t_L g7211 ( 
.A(n_7047),
.Y(n_7211)
);

CKINVDCx5p33_ASAP7_75t_R g7212 ( 
.A(n_6843),
.Y(n_7212)
);

BUFx6f_ASAP7_75t_L g7213 ( 
.A(n_7065),
.Y(n_7213)
);

INVx1_ASAP7_75t_L g7214 ( 
.A(n_6557),
.Y(n_7214)
);

INVx2_ASAP7_75t_L g7215 ( 
.A(n_6585),
.Y(n_7215)
);

AND2x4_ASAP7_75t_L g7216 ( 
.A(n_6718),
.B(n_5389),
.Y(n_7216)
);

CKINVDCx5p33_ASAP7_75t_R g7217 ( 
.A(n_6844),
.Y(n_7217)
);

INVx1_ASAP7_75t_L g7218 ( 
.A(n_6569),
.Y(n_7218)
);

INVx1_ASAP7_75t_L g7219 ( 
.A(n_6574),
.Y(n_7219)
);

CKINVDCx5p33_ASAP7_75t_R g7220 ( 
.A(n_6905),
.Y(n_7220)
);

INVx1_ASAP7_75t_L g7221 ( 
.A(n_6576),
.Y(n_7221)
);

NAND2xp5_ASAP7_75t_SL g7222 ( 
.A(n_6666),
.B(n_4380),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_6577),
.Y(n_7223)
);

BUFx6f_ASAP7_75t_L g7224 ( 
.A(n_7070),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_6580),
.Y(n_7225)
);

INVx2_ASAP7_75t_L g7226 ( 
.A(n_6612),
.Y(n_7226)
);

INVx3_ASAP7_75t_L g7227 ( 
.A(n_6562),
.Y(n_7227)
);

CKINVDCx5p33_ASAP7_75t_R g7228 ( 
.A(n_6950),
.Y(n_7228)
);

BUFx2_ASAP7_75t_L g7229 ( 
.A(n_7090),
.Y(n_7229)
);

CKINVDCx5p33_ASAP7_75t_R g7230 ( 
.A(n_6979),
.Y(n_7230)
);

AND2x2_ASAP7_75t_SL g7231 ( 
.A(n_6630),
.B(n_4616),
.Y(n_7231)
);

NOR2xp33_ASAP7_75t_R g7232 ( 
.A(n_6724),
.B(n_6886),
.Y(n_7232)
);

INVx2_ASAP7_75t_L g7233 ( 
.A(n_6620),
.Y(n_7233)
);

CKINVDCx5p33_ASAP7_75t_R g7234 ( 
.A(n_6776),
.Y(n_7234)
);

CKINVDCx5p33_ASAP7_75t_R g7235 ( 
.A(n_6779),
.Y(n_7235)
);

OAI21x1_ASAP7_75t_L g7236 ( 
.A1(n_6809),
.A2(n_4640),
.B(n_4626),
.Y(n_7236)
);

HB1xp67_ASAP7_75t_L g7237 ( 
.A(n_6583),
.Y(n_7237)
);

CKINVDCx5p33_ASAP7_75t_R g7238 ( 
.A(n_6784),
.Y(n_7238)
);

HB1xp67_ASAP7_75t_L g7239 ( 
.A(n_7043),
.Y(n_7239)
);

BUFx6f_ASAP7_75t_L g7240 ( 
.A(n_7078),
.Y(n_7240)
);

INVx1_ASAP7_75t_SL g7241 ( 
.A(n_6563),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_6599),
.Y(n_7242)
);

CKINVDCx20_ASAP7_75t_R g7243 ( 
.A(n_7041),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_6601),
.Y(n_7244)
);

BUFx2_ASAP7_75t_L g7245 ( 
.A(n_6598),
.Y(n_7245)
);

NOR2xp33_ASAP7_75t_R g7246 ( 
.A(n_6897),
.B(n_5392),
.Y(n_7246)
);

NOR2xp33_ASAP7_75t_L g7247 ( 
.A(n_6674),
.B(n_5178),
.Y(n_7247)
);

CKINVDCx20_ASAP7_75t_R g7248 ( 
.A(n_6629),
.Y(n_7248)
);

AND2x4_ASAP7_75t_L g7249 ( 
.A(n_6719),
.B(n_5444),
.Y(n_7249)
);

INVxp67_ASAP7_75t_L g7250 ( 
.A(n_7062),
.Y(n_7250)
);

INVx2_ASAP7_75t_L g7251 ( 
.A(n_6622),
.Y(n_7251)
);

NAND2xp5_ASAP7_75t_L g7252 ( 
.A(n_7081),
.B(n_4381),
.Y(n_7252)
);

NAND2xp5_ASAP7_75t_L g7253 ( 
.A(n_6638),
.B(n_4384),
.Y(n_7253)
);

INVx2_ASAP7_75t_L g7254 ( 
.A(n_6626),
.Y(n_7254)
);

CKINVDCx20_ASAP7_75t_R g7255 ( 
.A(n_6757),
.Y(n_7255)
);

BUFx6f_ASAP7_75t_L g7256 ( 
.A(n_7080),
.Y(n_7256)
);

CKINVDCx5p33_ASAP7_75t_R g7257 ( 
.A(n_6786),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_6608),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_L g7259 ( 
.A(n_6643),
.B(n_6652),
.Y(n_7259)
);

NOR2xp33_ASAP7_75t_L g7260 ( 
.A(n_6763),
.B(n_5231),
.Y(n_7260)
);

NAND2xp5_ASAP7_75t_L g7261 ( 
.A(n_6663),
.B(n_4385),
.Y(n_7261)
);

HB1xp67_ASAP7_75t_L g7262 ( 
.A(n_7066),
.Y(n_7262)
);

CKINVDCx20_ASAP7_75t_R g7263 ( 
.A(n_6796),
.Y(n_7263)
);

INVx2_ASAP7_75t_L g7264 ( 
.A(n_6859),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_6609),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_6610),
.Y(n_7266)
);

CKINVDCx5p33_ASAP7_75t_R g7267 ( 
.A(n_6806),
.Y(n_7267)
);

INVx2_ASAP7_75t_SL g7268 ( 
.A(n_6582),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_6614),
.Y(n_7269)
);

NAND2xp33_ASAP7_75t_SL g7270 ( 
.A(n_6684),
.B(n_5482),
.Y(n_7270)
);

INVx2_ASAP7_75t_L g7271 ( 
.A(n_6864),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_6617),
.Y(n_7272)
);

NAND2xp5_ASAP7_75t_L g7273 ( 
.A(n_6678),
.B(n_4386),
.Y(n_7273)
);

AND2x4_ASAP7_75t_L g7274 ( 
.A(n_6807),
.B(n_6842),
.Y(n_7274)
);

XNOR2xp5_ASAP7_75t_L g7275 ( 
.A(n_7076),
.B(n_5494),
.Y(n_7275)
);

CKINVDCx20_ASAP7_75t_R g7276 ( 
.A(n_6810),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_6618),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_6621),
.Y(n_7278)
);

CKINVDCx20_ASAP7_75t_R g7279 ( 
.A(n_6831),
.Y(n_7279)
);

INVx2_ASAP7_75t_L g7280 ( 
.A(n_6890),
.Y(n_7280)
);

CKINVDCx5p33_ASAP7_75t_R g7281 ( 
.A(n_6818),
.Y(n_7281)
);

BUFx3_ASAP7_75t_L g7282 ( 
.A(n_6834),
.Y(n_7282)
);

INVx1_ASAP7_75t_L g7283 ( 
.A(n_6641),
.Y(n_7283)
);

CKINVDCx20_ASAP7_75t_R g7284 ( 
.A(n_6989),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_6646),
.Y(n_7285)
);

INVx3_ASAP7_75t_L g7286 ( 
.A(n_7012),
.Y(n_7286)
);

CKINVDCx5p33_ASAP7_75t_R g7287 ( 
.A(n_6822),
.Y(n_7287)
);

BUFx6f_ASAP7_75t_L g7288 ( 
.A(n_7086),
.Y(n_7288)
);

INVx1_ASAP7_75t_L g7289 ( 
.A(n_6649),
.Y(n_7289)
);

CKINVDCx20_ASAP7_75t_R g7290 ( 
.A(n_6861),
.Y(n_7290)
);

INVx1_ASAP7_75t_L g7291 ( 
.A(n_6679),
.Y(n_7291)
);

NAND2xp5_ASAP7_75t_L g7292 ( 
.A(n_6710),
.B(n_4387),
.Y(n_7292)
);

CKINVDCx5p33_ASAP7_75t_R g7293 ( 
.A(n_6836),
.Y(n_7293)
);

BUFx6f_ASAP7_75t_L g7294 ( 
.A(n_6521),
.Y(n_7294)
);

INVx5_ASAP7_75t_L g7295 ( 
.A(n_6879),
.Y(n_7295)
);

CKINVDCx5p33_ASAP7_75t_R g7296 ( 
.A(n_6840),
.Y(n_7296)
);

BUFx6f_ASAP7_75t_L g7297 ( 
.A(n_6526),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_6691),
.Y(n_7298)
);

NAND2xp5_ASAP7_75t_L g7299 ( 
.A(n_6721),
.B(n_4388),
.Y(n_7299)
);

AND2x2_ASAP7_75t_L g7300 ( 
.A(n_6513),
.B(n_5496),
.Y(n_7300)
);

CKINVDCx20_ASAP7_75t_R g7301 ( 
.A(n_6654),
.Y(n_7301)
);

OAI22xp5_ASAP7_75t_SL g7302 ( 
.A1(n_6570),
.A2(n_5501),
.B1(n_5504),
.B2(n_5500),
.Y(n_7302)
);

CKINVDCx20_ASAP7_75t_R g7303 ( 
.A(n_6668),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_6694),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_6709),
.Y(n_7305)
);

CKINVDCx5p33_ASAP7_75t_R g7306 ( 
.A(n_6850),
.Y(n_7306)
);

INVx2_ASAP7_75t_L g7307 ( 
.A(n_6899),
.Y(n_7307)
);

INVx1_ASAP7_75t_L g7308 ( 
.A(n_6720),
.Y(n_7308)
);

INVx1_ASAP7_75t_L g7309 ( 
.A(n_6732),
.Y(n_7309)
);

CKINVDCx20_ASAP7_75t_R g7310 ( 
.A(n_6690),
.Y(n_7310)
);

INVx1_ASAP7_75t_L g7311 ( 
.A(n_6738),
.Y(n_7311)
);

INVx6_ASAP7_75t_L g7312 ( 
.A(n_6693),
.Y(n_7312)
);

CKINVDCx5p33_ASAP7_75t_R g7313 ( 
.A(n_6869),
.Y(n_7313)
);

AND2x6_ASAP7_75t_L g7314 ( 
.A(n_6715),
.B(n_4815),
.Y(n_7314)
);

XNOR2xp5_ASAP7_75t_L g7315 ( 
.A(n_6868),
.B(n_5256),
.Y(n_7315)
);

CKINVDCx5p33_ASAP7_75t_R g7316 ( 
.A(n_6875),
.Y(n_7316)
);

INVx3_ASAP7_75t_L g7317 ( 
.A(n_7055),
.Y(n_7317)
);

INVx1_ASAP7_75t_L g7318 ( 
.A(n_6755),
.Y(n_7318)
);

INVxp67_ASAP7_75t_L g7319 ( 
.A(n_6589),
.Y(n_7319)
);

INVx1_ASAP7_75t_L g7320 ( 
.A(n_6767),
.Y(n_7320)
);

CKINVDCx5p33_ASAP7_75t_R g7321 ( 
.A(n_6889),
.Y(n_7321)
);

BUFx6f_ASAP7_75t_L g7322 ( 
.A(n_6529),
.Y(n_7322)
);

CKINVDCx5p33_ASAP7_75t_R g7323 ( 
.A(n_6916),
.Y(n_7323)
);

INVx2_ASAP7_75t_L g7324 ( 
.A(n_6918),
.Y(n_7324)
);

CKINVDCx5p33_ASAP7_75t_R g7325 ( 
.A(n_6923),
.Y(n_7325)
);

AND2x2_ASAP7_75t_L g7326 ( 
.A(n_6524),
.B(n_4890),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_6771),
.Y(n_7327)
);

NOR2xp33_ASAP7_75t_L g7328 ( 
.A(n_6930),
.B(n_5264),
.Y(n_7328)
);

HB1xp67_ASAP7_75t_L g7329 ( 
.A(n_6855),
.Y(n_7329)
);

BUFx6f_ASAP7_75t_L g7330 ( 
.A(n_6714),
.Y(n_7330)
);

CKINVDCx20_ASAP7_75t_R g7331 ( 
.A(n_6656),
.Y(n_7331)
);

INVx1_ASAP7_75t_L g7332 ( 
.A(n_6775),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6800),
.Y(n_7333)
);

CKINVDCx5p33_ASAP7_75t_R g7334 ( 
.A(n_6942),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_6817),
.Y(n_7335)
);

INVx1_ASAP7_75t_L g7336 ( 
.A(n_6826),
.Y(n_7336)
);

NOR2xp33_ASAP7_75t_R g7337 ( 
.A(n_6722),
.B(n_6726),
.Y(n_7337)
);

INVx3_ASAP7_75t_L g7338 ( 
.A(n_6512),
.Y(n_7338)
);

CKINVDCx5p33_ASAP7_75t_R g7339 ( 
.A(n_6944),
.Y(n_7339)
);

NAND2xp33_ASAP7_75t_L g7340 ( 
.A(n_6948),
.B(n_4390),
.Y(n_7340)
);

CKINVDCx20_ASAP7_75t_R g7341 ( 
.A(n_6670),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_SL g7342 ( 
.A(n_7051),
.B(n_4393),
.Y(n_7342)
);

CKINVDCx5p33_ASAP7_75t_R g7343 ( 
.A(n_6949),
.Y(n_7343)
);

CKINVDCx5p33_ASAP7_75t_R g7344 ( 
.A(n_6955),
.Y(n_7344)
);

NOR2xp33_ASAP7_75t_R g7345 ( 
.A(n_6736),
.B(n_4394),
.Y(n_7345)
);

INVx1_ASAP7_75t_L g7346 ( 
.A(n_6827),
.Y(n_7346)
);

CKINVDCx5p33_ASAP7_75t_R g7347 ( 
.A(n_6737),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_6846),
.Y(n_7348)
);

INVx2_ASAP7_75t_L g7349 ( 
.A(n_6921),
.Y(n_7349)
);

CKINVDCx5p33_ASAP7_75t_R g7350 ( 
.A(n_6756),
.Y(n_7350)
);

CKINVDCx5p33_ASAP7_75t_R g7351 ( 
.A(n_6768),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6847),
.Y(n_7352)
);

INVx3_ASAP7_75t_L g7353 ( 
.A(n_7026),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_6852),
.Y(n_7354)
);

CKINVDCx20_ASAP7_75t_R g7355 ( 
.A(n_6689),
.Y(n_7355)
);

CKINVDCx5p33_ASAP7_75t_R g7356 ( 
.A(n_7087),
.Y(n_7356)
);

CKINVDCx5p33_ASAP7_75t_R g7357 ( 
.A(n_6873),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_6853),
.Y(n_7358)
);

CKINVDCx11_ASAP7_75t_R g7359 ( 
.A(n_6702),
.Y(n_7359)
);

CKINVDCx20_ASAP7_75t_R g7360 ( 
.A(n_6717),
.Y(n_7360)
);

INVx2_ASAP7_75t_L g7361 ( 
.A(n_6928),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_6854),
.Y(n_7362)
);

CKINVDCx5p33_ASAP7_75t_R g7363 ( 
.A(n_6699),
.Y(n_7363)
);

INVx2_ASAP7_75t_L g7364 ( 
.A(n_6933),
.Y(n_7364)
);

CKINVDCx20_ASAP7_75t_R g7365 ( 
.A(n_6731),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_6935),
.Y(n_7366)
);

CKINVDCx20_ASAP7_75t_R g7367 ( 
.A(n_6830),
.Y(n_7367)
);

CKINVDCx5p33_ASAP7_75t_R g7368 ( 
.A(n_6723),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_6858),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_6860),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_6862),
.Y(n_7371)
);

CKINVDCx20_ASAP7_75t_R g7372 ( 
.A(n_6863),
.Y(n_7372)
);

INVx2_ASAP7_75t_L g7373 ( 
.A(n_6940),
.Y(n_7373)
);

INVxp67_ASAP7_75t_SL g7374 ( 
.A(n_6538),
.Y(n_7374)
);

NAND2xp33_ASAP7_75t_L g7375 ( 
.A(n_6799),
.B(n_4395),
.Y(n_7375)
);

INVx2_ASAP7_75t_L g7376 ( 
.A(n_6945),
.Y(n_7376)
);

CKINVDCx20_ASAP7_75t_R g7377 ( 
.A(n_6882),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_6865),
.Y(n_7378)
);

INVx2_ASAP7_75t_L g7379 ( 
.A(n_6965),
.Y(n_7379)
);

INVx1_ASAP7_75t_L g7380 ( 
.A(n_6870),
.Y(n_7380)
);

CKINVDCx5p33_ASAP7_75t_R g7381 ( 
.A(n_6804),
.Y(n_7381)
);

CKINVDCx5p33_ASAP7_75t_R g7382 ( 
.A(n_6816),
.Y(n_7382)
);

NAND2xp5_ASAP7_75t_L g7383 ( 
.A(n_6741),
.B(n_4396),
.Y(n_7383)
);

INVx1_ASAP7_75t_L g7384 ( 
.A(n_6871),
.Y(n_7384)
);

CKINVDCx5p33_ASAP7_75t_R g7385 ( 
.A(n_6872),
.Y(n_7385)
);

CKINVDCx20_ASAP7_75t_R g7386 ( 
.A(n_6895),
.Y(n_7386)
);

INVxp67_ASAP7_75t_L g7387 ( 
.A(n_6555),
.Y(n_7387)
);

INVx1_ASAP7_75t_L g7388 ( 
.A(n_6888),
.Y(n_7388)
);

CKINVDCx5p33_ASAP7_75t_R g7389 ( 
.A(n_6906),
.Y(n_7389)
);

CKINVDCx5p33_ASAP7_75t_R g7390 ( 
.A(n_6919),
.Y(n_7390)
);

NAND2xp5_ASAP7_75t_L g7391 ( 
.A(n_6761),
.B(n_4397),
.Y(n_7391)
);

CKINVDCx5p33_ASAP7_75t_R g7392 ( 
.A(n_6924),
.Y(n_7392)
);

INVx1_ASAP7_75t_L g7393 ( 
.A(n_6892),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_6783),
.B(n_4400),
.Y(n_7394)
);

CKINVDCx5p33_ASAP7_75t_R g7395 ( 
.A(n_6934),
.Y(n_7395)
);

NAND2xp5_ASAP7_75t_L g7396 ( 
.A(n_6819),
.B(n_4401),
.Y(n_7396)
);

CKINVDCx5p33_ASAP7_75t_R g7397 ( 
.A(n_6990),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6894),
.Y(n_7398)
);

INVx2_ASAP7_75t_L g7399 ( 
.A(n_6968),
.Y(n_7399)
);

HB1xp67_ASAP7_75t_L g7400 ( 
.A(n_6821),
.Y(n_7400)
);

CKINVDCx5p33_ASAP7_75t_R g7401 ( 
.A(n_6625),
.Y(n_7401)
);

INVx2_ASAP7_75t_L g7402 ( 
.A(n_6970),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_6896),
.Y(n_7403)
);

INVx3_ASAP7_75t_L g7404 ( 
.A(n_7035),
.Y(n_7404)
);

NAND2x1_ASAP7_75t_L g7405 ( 
.A(n_6591),
.B(n_4697),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_6911),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_6920),
.Y(n_7407)
);

CKINVDCx5p33_ASAP7_75t_R g7408 ( 
.A(n_6664),
.Y(n_7408)
);

NAND2xp5_ASAP7_75t_L g7409 ( 
.A(n_6828),
.B(n_4402),
.Y(n_7409)
);

INVx1_ASAP7_75t_L g7410 ( 
.A(n_6922),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_6925),
.Y(n_7411)
);

NOR2xp33_ASAP7_75t_L g7412 ( 
.A(n_6631),
.B(n_5267),
.Y(n_7412)
);

INVx1_ASAP7_75t_L g7413 ( 
.A(n_6926),
.Y(n_7413)
);

CKINVDCx5p33_ASAP7_75t_R g7414 ( 
.A(n_6688),
.Y(n_7414)
);

BUFx6f_ASAP7_75t_L g7415 ( 
.A(n_7046),
.Y(n_7415)
);

BUFx6f_ASAP7_75t_L g7416 ( 
.A(n_6999),
.Y(n_7416)
);

INVx2_ASAP7_75t_L g7417 ( 
.A(n_6982),
.Y(n_7417)
);

INVx2_ASAP7_75t_L g7418 ( 
.A(n_6983),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_6927),
.Y(n_7419)
);

NOR2xp33_ASAP7_75t_SL g7420 ( 
.A(n_6777),
.B(n_5307),
.Y(n_7420)
);

AND2x2_ASAP7_75t_L g7421 ( 
.A(n_6575),
.B(n_4890),
.Y(n_7421)
);

CKINVDCx5p33_ASAP7_75t_R g7422 ( 
.A(n_6914),
.Y(n_7422)
);

HB1xp67_ASAP7_75t_L g7423 ( 
.A(n_6829),
.Y(n_7423)
);

BUFx6f_ASAP7_75t_L g7424 ( 
.A(n_7007),
.Y(n_7424)
);

INVxp67_ASAP7_75t_L g7425 ( 
.A(n_6541),
.Y(n_7425)
);

CKINVDCx20_ASAP7_75t_R g7426 ( 
.A(n_6941),
.Y(n_7426)
);

NAND2xp33_ASAP7_75t_SL g7427 ( 
.A(n_6849),
.B(n_4403),
.Y(n_7427)
);

INVx3_ASAP7_75t_L g7428 ( 
.A(n_7083),
.Y(n_7428)
);

INVx1_ASAP7_75t_L g7429 ( 
.A(n_6938),
.Y(n_7429)
);

OAI21x1_ASAP7_75t_L g7430 ( 
.A1(n_6832),
.A2(n_4705),
.B(n_4657),
.Y(n_7430)
);

CKINVDCx5p33_ASAP7_75t_R g7431 ( 
.A(n_6998),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_6939),
.Y(n_7432)
);

HB1xp67_ASAP7_75t_L g7433 ( 
.A(n_6877),
.Y(n_7433)
);

NAND2xp5_ASAP7_75t_L g7434 ( 
.A(n_6841),
.B(n_4404),
.Y(n_7434)
);

INVx1_ASAP7_75t_L g7435 ( 
.A(n_6943),
.Y(n_7435)
);

INVxp67_ASAP7_75t_L g7436 ( 
.A(n_6541),
.Y(n_7436)
);

CKINVDCx5p33_ASAP7_75t_R g7437 ( 
.A(n_7091),
.Y(n_7437)
);

CKINVDCx20_ASAP7_75t_R g7438 ( 
.A(n_6974),
.Y(n_7438)
);

BUFx2_ASAP7_75t_L g7439 ( 
.A(n_7089),
.Y(n_7439)
);

CKINVDCx5p33_ASAP7_75t_R g7440 ( 
.A(n_7091),
.Y(n_7440)
);

BUFx6f_ASAP7_75t_L g7441 ( 
.A(n_6956),
.Y(n_7441)
);

NAND2xp5_ASAP7_75t_L g7442 ( 
.A(n_6885),
.B(n_4405),
.Y(n_7442)
);

CKINVDCx5p33_ASAP7_75t_R g7443 ( 
.A(n_6644),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_6952),
.Y(n_7444)
);

CKINVDCx5p33_ASAP7_75t_R g7445 ( 
.A(n_6671),
.Y(n_7445)
);

BUFx3_ASAP7_75t_L g7446 ( 
.A(n_6967),
.Y(n_7446)
);

INVx1_ASAP7_75t_L g7447 ( 
.A(n_6961),
.Y(n_7447)
);

CKINVDCx5p33_ASAP7_75t_R g7448 ( 
.A(n_6590),
.Y(n_7448)
);

INVx3_ASAP7_75t_L g7449 ( 
.A(n_6636),
.Y(n_7449)
);

INVx2_ASAP7_75t_L g7450 ( 
.A(n_6987),
.Y(n_7450)
);

CKINVDCx5p33_ASAP7_75t_R g7451 ( 
.A(n_6706),
.Y(n_7451)
);

INVx1_ASAP7_75t_L g7452 ( 
.A(n_6972),
.Y(n_7452)
);

OA21x2_ASAP7_75t_L g7453 ( 
.A1(n_6904),
.A2(n_4823),
.B(n_4819),
.Y(n_7453)
);

INVx1_ASAP7_75t_L g7454 ( 
.A(n_6976),
.Y(n_7454)
);

INVx2_ASAP7_75t_L g7455 ( 
.A(n_6991),
.Y(n_7455)
);

INVx1_ASAP7_75t_L g7456 ( 
.A(n_6980),
.Y(n_7456)
);

CKINVDCx5p33_ASAP7_75t_R g7457 ( 
.A(n_6794),
.Y(n_7457)
);

INVx3_ASAP7_75t_L g7458 ( 
.A(n_6637),
.Y(n_7458)
);

INVx1_ASAP7_75t_L g7459 ( 
.A(n_6981),
.Y(n_7459)
);

CKINVDCx20_ASAP7_75t_R g7460 ( 
.A(n_6985),
.Y(n_7460)
);

NOR2xp33_ASAP7_75t_R g7461 ( 
.A(n_6734),
.B(n_4409),
.Y(n_7461)
);

CKINVDCx20_ASAP7_75t_R g7462 ( 
.A(n_6937),
.Y(n_7462)
);

AND2x4_ASAP7_75t_L g7463 ( 
.A(n_6744),
.B(n_5355),
.Y(n_7463)
);

INVx1_ASAP7_75t_L g7464 ( 
.A(n_6628),
.Y(n_7464)
);

CKINVDCx5p33_ASAP7_75t_R g7465 ( 
.A(n_6659),
.Y(n_7465)
);

INVx3_ASAP7_75t_L g7466 ( 
.A(n_6647),
.Y(n_7466)
);

HB1xp67_ASAP7_75t_L g7467 ( 
.A(n_6639),
.Y(n_7467)
);

AND2x2_ASAP7_75t_SL g7468 ( 
.A(n_7021),
.B(n_4716),
.Y(n_7468)
);

CKINVDCx5p33_ASAP7_75t_R g7469 ( 
.A(n_7033),
.Y(n_7469)
);

CKINVDCx5p33_ASAP7_75t_R g7470 ( 
.A(n_6857),
.Y(n_7470)
);

CKINVDCx5p33_ASAP7_75t_R g7471 ( 
.A(n_6751),
.Y(n_7471)
);

INVx2_ASAP7_75t_L g7472 ( 
.A(n_6595),
.Y(n_7472)
);

AND2x2_ASAP7_75t_L g7473 ( 
.A(n_6891),
.B(n_4894),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_6645),
.Y(n_7474)
);

NAND2xp5_ASAP7_75t_L g7475 ( 
.A(n_6901),
.B(n_4411),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_6650),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_6657),
.Y(n_7477)
);

CKINVDCx5p33_ASAP7_75t_R g7478 ( 
.A(n_6792),
.Y(n_7478)
);

NOR2xp33_ASAP7_75t_R g7479 ( 
.A(n_6594),
.B(n_4412),
.Y(n_7479)
);

NAND2xp5_ASAP7_75t_L g7480 ( 
.A(n_6902),
.B(n_4415),
.Y(n_7480)
);

AND2x2_ASAP7_75t_L g7481 ( 
.A(n_6667),
.B(n_6603),
.Y(n_7481)
);

NAND2xp33_ASAP7_75t_R g7482 ( 
.A(n_6837),
.B(n_4416),
.Y(n_7482)
);

HB1xp67_ASAP7_75t_L g7483 ( 
.A(n_6653),
.Y(n_7483)
);

NOR2xp33_ASAP7_75t_L g7484 ( 
.A(n_6551),
.B(n_5427),
.Y(n_7484)
);

AND2x2_ASAP7_75t_L g7485 ( 
.A(n_6624),
.B(n_4894),
.Y(n_7485)
);

BUFx6f_ASAP7_75t_L g7486 ( 
.A(n_6973),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_L g7487 ( 
.A(n_6903),
.B(n_6908),
.Y(n_7487)
);

INVx2_ASAP7_75t_L g7488 ( 
.A(n_6600),
.Y(n_7488)
);

CKINVDCx5p33_ASAP7_75t_R g7489 ( 
.A(n_6739),
.Y(n_7489)
);

INVx1_ASAP7_75t_L g7490 ( 
.A(n_6658),
.Y(n_7490)
);

INVx1_ASAP7_75t_L g7491 ( 
.A(n_6669),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_L g7492 ( 
.A(n_6915),
.B(n_4417),
.Y(n_7492)
);

NOR3xp33_ASAP7_75t_L g7493 ( 
.A(n_6825),
.B(n_5503),
.C(n_4826),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_6673),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_6698),
.Y(n_7495)
);

BUFx6f_ASAP7_75t_L g7496 ( 
.A(n_6651),
.Y(n_7496)
);

INVx2_ASAP7_75t_L g7497 ( 
.A(n_6597),
.Y(n_7497)
);

NAND2xp5_ASAP7_75t_L g7498 ( 
.A(n_6936),
.B(n_4421),
.Y(n_7498)
);

INVx3_ASAP7_75t_L g7499 ( 
.A(n_6660),
.Y(n_7499)
);

AND2x4_ASAP7_75t_L g7500 ( 
.A(n_6519),
.B(n_4825),
.Y(n_7500)
);

NOR2xp33_ASAP7_75t_L g7501 ( 
.A(n_6743),
.B(n_4425),
.Y(n_7501)
);

CKINVDCx20_ASAP7_75t_R g7502 ( 
.A(n_7082),
.Y(n_7502)
);

CKINVDCx5p33_ASAP7_75t_R g7503 ( 
.A(n_6874),
.Y(n_7503)
);

NOR2xp33_ASAP7_75t_R g7504 ( 
.A(n_6963),
.B(n_4426),
.Y(n_7504)
);

CKINVDCx5p33_ASAP7_75t_R g7505 ( 
.A(n_6954),
.Y(n_7505)
);

INVx2_ASAP7_75t_L g7506 ( 
.A(n_6700),
.Y(n_7506)
);

CKINVDCx5p33_ASAP7_75t_R g7507 ( 
.A(n_6856),
.Y(n_7507)
);

AND2x2_ASAP7_75t_L g7508 ( 
.A(n_6801),
.B(n_4897),
.Y(n_7508)
);

NAND2xp5_ASAP7_75t_L g7509 ( 
.A(n_6977),
.B(n_6745),
.Y(n_7509)
);

NAND2xp5_ASAP7_75t_L g7510 ( 
.A(n_6701),
.B(n_4428),
.Y(n_7510)
);

HB1xp67_ASAP7_75t_L g7511 ( 
.A(n_6909),
.Y(n_7511)
);

CKINVDCx5p33_ASAP7_75t_R g7512 ( 
.A(n_7037),
.Y(n_7512)
);

INVx1_ASAP7_75t_L g7513 ( 
.A(n_6523),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_6525),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7011),
.Y(n_7515)
);

INVx2_ASAP7_75t_L g7516 ( 
.A(n_6995),
.Y(n_7516)
);

NAND2xp5_ASAP7_75t_L g7517 ( 
.A(n_6604),
.B(n_4431),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_7019),
.Y(n_7518)
);

BUFx6f_ASAP7_75t_L g7519 ( 
.A(n_6661),
.Y(n_7519)
);

NAND2xp5_ASAP7_75t_L g7520 ( 
.A(n_6623),
.B(n_4435),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7029),
.Y(n_7521)
);

INVx2_ASAP7_75t_L g7522 ( 
.A(n_7030),
.Y(n_7522)
);

INVx2_ASAP7_75t_L g7523 ( 
.A(n_7038),
.Y(n_7523)
);

CKINVDCx20_ASAP7_75t_R g7524 ( 
.A(n_6534),
.Y(n_7524)
);

INVx1_ASAP7_75t_L g7525 ( 
.A(n_7045),
.Y(n_7525)
);

BUFx6f_ASAP7_75t_L g7526 ( 
.A(n_6662),
.Y(n_7526)
);

AND2x2_ASAP7_75t_L g7527 ( 
.A(n_6812),
.B(n_6785),
.Y(n_7527)
);

CKINVDCx20_ASAP7_75t_R g7528 ( 
.A(n_7058),
.Y(n_7528)
);

INVx1_ASAP7_75t_L g7529 ( 
.A(n_7067),
.Y(n_7529)
);

INVx1_ASAP7_75t_L g7530 ( 
.A(n_7072),
.Y(n_7530)
);

INVx1_ASAP7_75t_L g7531 ( 
.A(n_7079),
.Y(n_7531)
);

CKINVDCx5p33_ASAP7_75t_R g7532 ( 
.A(n_6573),
.Y(n_7532)
);

NAND2xp5_ASAP7_75t_L g7533 ( 
.A(n_7085),
.B(n_4436),
.Y(n_7533)
);

INVx2_ASAP7_75t_L g7534 ( 
.A(n_7003),
.Y(n_7534)
);

NAND2xp5_ASAP7_75t_SL g7535 ( 
.A(n_6572),
.B(n_4437),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_6752),
.Y(n_7536)
);

CKINVDCx16_ASAP7_75t_R g7537 ( 
.A(n_6898),
.Y(n_7537)
);

NAND2xp33_ASAP7_75t_R g7538 ( 
.A(n_6900),
.B(n_4438),
.Y(n_7538)
);

BUFx6f_ASAP7_75t_L g7539 ( 
.A(n_6675),
.Y(n_7539)
);

CKINVDCx5p33_ASAP7_75t_R g7540 ( 
.A(n_6789),
.Y(n_7540)
);

BUFx10_ASAP7_75t_L g7541 ( 
.A(n_6971),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_6787),
.Y(n_7542)
);

CKINVDCx5p33_ASAP7_75t_R g7543 ( 
.A(n_6789),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_6753),
.Y(n_7544)
);

INVx2_ASAP7_75t_L g7545 ( 
.A(n_7005),
.Y(n_7545)
);

BUFx10_ASAP7_75t_L g7546 ( 
.A(n_6725),
.Y(n_7546)
);

HB1xp67_ASAP7_75t_L g7547 ( 
.A(n_6797),
.Y(n_7547)
);

CKINVDCx20_ASAP7_75t_R g7548 ( 
.A(n_6845),
.Y(n_7548)
);

BUFx6f_ASAP7_75t_L g7549 ( 
.A(n_6680),
.Y(n_7549)
);

CKINVDCx20_ASAP7_75t_R g7550 ( 
.A(n_6867),
.Y(n_7550)
);

INVx3_ASAP7_75t_L g7551 ( 
.A(n_6682),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_6880),
.Y(n_7552)
);

NAND2xp5_ASAP7_75t_L g7553 ( 
.A(n_7059),
.B(n_4439),
.Y(n_7553)
);

CKINVDCx5p33_ASAP7_75t_R g7554 ( 
.A(n_6907),
.Y(n_7554)
);

INVx2_ASAP7_75t_L g7555 ( 
.A(n_6996),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_6883),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_6931),
.Y(n_7557)
);

BUFx6f_ASAP7_75t_L g7558 ( 
.A(n_6687),
.Y(n_7558)
);

CKINVDCx5p33_ASAP7_75t_R g7559 ( 
.A(n_7006),
.Y(n_7559)
);

NAND2xp5_ASAP7_75t_L g7560 ( 
.A(n_6959),
.B(n_4440),
.Y(n_7560)
);

CKINVDCx16_ASAP7_75t_R g7561 ( 
.A(n_6835),
.Y(n_7561)
);

CKINVDCx5p33_ASAP7_75t_R g7562 ( 
.A(n_6543),
.Y(n_7562)
);

INVx1_ASAP7_75t_L g7563 ( 
.A(n_6957),
.Y(n_7563)
);

OA21x2_ASAP7_75t_L g7564 ( 
.A1(n_6932),
.A2(n_4832),
.B(n_4830),
.Y(n_7564)
);

BUFx6f_ASAP7_75t_L g7565 ( 
.A(n_6692),
.Y(n_7565)
);

CKINVDCx5p33_ASAP7_75t_R g7566 ( 
.A(n_6960),
.Y(n_7566)
);

INVx2_ASAP7_75t_L g7567 ( 
.A(n_7009),
.Y(n_7567)
);

CKINVDCx20_ASAP7_75t_R g7568 ( 
.A(n_6917),
.Y(n_7568)
);

CKINVDCx5p33_ASAP7_75t_R g7569 ( 
.A(n_6960),
.Y(n_7569)
);

CKINVDCx5p33_ASAP7_75t_R g7570 ( 
.A(n_6978),
.Y(n_7570)
);

INVx1_ASAP7_75t_L g7571 ( 
.A(n_6988),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_6735),
.Y(n_7572)
);

BUFx6f_ASAP7_75t_L g7573 ( 
.A(n_6695),
.Y(n_7573)
);

INVx5_ASAP7_75t_L g7574 ( 
.A(n_6978),
.Y(n_7574)
);

INVx5_ASAP7_75t_L g7575 ( 
.A(n_6803),
.Y(n_7575)
);

AND2x4_ASAP7_75t_L g7576 ( 
.A(n_6820),
.B(n_4836),
.Y(n_7576)
);

INVx3_ASAP7_75t_L g7577 ( 
.A(n_6713),
.Y(n_7577)
);

CKINVDCx20_ASAP7_75t_R g7578 ( 
.A(n_6805),
.Y(n_7578)
);

NOR2xp33_ASAP7_75t_R g7579 ( 
.A(n_7001),
.B(n_4441),
.Y(n_7579)
);

BUFx6f_ASAP7_75t_L g7580 ( 
.A(n_6587),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_6561),
.Y(n_7581)
);

CKINVDCx16_ASAP7_75t_R g7582 ( 
.A(n_7049),
.Y(n_7582)
);

INVx2_ASAP7_75t_L g7583 ( 
.A(n_6514),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_6579),
.Y(n_7584)
);

HB1xp67_ASAP7_75t_L g7585 ( 
.A(n_6568),
.Y(n_7585)
);

BUFx6f_ASAP7_75t_L g7586 ( 
.A(n_6593),
.Y(n_7586)
);

INVx1_ASAP7_75t_L g7587 ( 
.A(n_6615),
.Y(n_7587)
);

BUFx6f_ASAP7_75t_L g7588 ( 
.A(n_6696),
.Y(n_7588)
);

INVx2_ASAP7_75t_L g7589 ( 
.A(n_6518),
.Y(n_7589)
);

AO21x2_ASAP7_75t_L g7590 ( 
.A1(n_6549),
.A2(n_4847),
.B(n_4838),
.Y(n_7590)
);

CKINVDCx5p33_ASAP7_75t_R g7591 ( 
.A(n_6740),
.Y(n_7591)
);

AND2x2_ASAP7_75t_L g7592 ( 
.A(n_6764),
.B(n_4897),
.Y(n_7592)
);

INVx2_ASAP7_75t_L g7593 ( 
.A(n_6520),
.Y(n_7593)
);

CKINVDCx5p33_ASAP7_75t_R g7594 ( 
.A(n_6760),
.Y(n_7594)
);

CKINVDCx20_ASAP7_75t_R g7595 ( 
.A(n_7060),
.Y(n_7595)
);

INVx1_ASAP7_75t_L g7596 ( 
.A(n_6616),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_6672),
.Y(n_7597)
);

AND2x2_ASAP7_75t_L g7598 ( 
.A(n_6676),
.B(n_4948),
.Y(n_7598)
);

CKINVDCx16_ASAP7_75t_R g7599 ( 
.A(n_7077),
.Y(n_7599)
);

AOI22xp5_ASAP7_75t_L g7600 ( 
.A1(n_6635),
.A2(n_4442),
.B1(n_4448),
.B2(n_4444),
.Y(n_7600)
);

NAND2xp5_ASAP7_75t_L g7601 ( 
.A(n_7024),
.B(n_4452),
.Y(n_7601)
);

CKINVDCx20_ASAP7_75t_R g7602 ( 
.A(n_7027),
.Y(n_7602)
);

NOR2xp33_ASAP7_75t_R g7603 ( 
.A(n_6546),
.B(n_4455),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_6697),
.Y(n_7604)
);

CKINVDCx20_ASAP7_75t_R g7605 ( 
.A(n_7052),
.Y(n_7605)
);

INVx2_ASAP7_75t_L g7606 ( 
.A(n_7013),
.Y(n_7606)
);

INVx3_ASAP7_75t_L g7607 ( 
.A(n_6567),
.Y(n_7607)
);

CKINVDCx5p33_ASAP7_75t_R g7608 ( 
.A(n_6823),
.Y(n_7608)
);

CKINVDCx5p33_ASAP7_75t_R g7609 ( 
.A(n_6887),
.Y(n_7609)
);

BUFx2_ASAP7_75t_L g7610 ( 
.A(n_6711),
.Y(n_7610)
);

INVx1_ASAP7_75t_L g7611 ( 
.A(n_6704),
.Y(n_7611)
);

BUFx6f_ASAP7_75t_L g7612 ( 
.A(n_6707),
.Y(n_7612)
);

INVx2_ASAP7_75t_L g7613 ( 
.A(n_7015),
.Y(n_7613)
);

CKINVDCx5p33_ASAP7_75t_R g7614 ( 
.A(n_6640),
.Y(n_7614)
);

NOR2xp33_ASAP7_75t_L g7615 ( 
.A(n_6969),
.B(n_4456),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_6705),
.Y(n_7616)
);

CKINVDCx5p33_ASAP7_75t_R g7617 ( 
.A(n_7008),
.Y(n_7617)
);

CKINVDCx16_ASAP7_75t_R g7618 ( 
.A(n_6584),
.Y(n_7618)
);

BUFx2_ASAP7_75t_L g7619 ( 
.A(n_6602),
.Y(n_7619)
);

CKINVDCx5p33_ASAP7_75t_R g7620 ( 
.A(n_6648),
.Y(n_7620)
);

AND2x2_ASAP7_75t_L g7621 ( 
.A(n_7036),
.B(n_4948),
.Y(n_7621)
);

CKINVDCx5p33_ASAP7_75t_R g7622 ( 
.A(n_7004),
.Y(n_7622)
);

INVx2_ASAP7_75t_L g7623 ( 
.A(n_7016),
.Y(n_7623)
);

INVx1_ASAP7_75t_L g7624 ( 
.A(n_6833),
.Y(n_7624)
);

AND2x2_ASAP7_75t_L g7625 ( 
.A(n_7039),
.B(n_4989),
.Y(n_7625)
);

INVx1_ASAP7_75t_L g7626 ( 
.A(n_6848),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_6958),
.Y(n_7627)
);

NOR2xp33_ASAP7_75t_R g7628 ( 
.A(n_6642),
.B(n_4457),
.Y(n_7628)
);

CKINVDCx5p33_ASAP7_75t_R g7629 ( 
.A(n_6632),
.Y(n_7629)
);

INVx1_ASAP7_75t_L g7630 ( 
.A(n_6962),
.Y(n_7630)
);

AND3x1_ASAP7_75t_L g7631 ( 
.A(n_6606),
.B(n_4858),
.C(n_4851),
.Y(n_7631)
);

INVx1_ASAP7_75t_L g7632 ( 
.A(n_6778),
.Y(n_7632)
);

INVx1_ASAP7_75t_L g7633 ( 
.A(n_6780),
.Y(n_7633)
);

NAND2xp5_ASAP7_75t_SL g7634 ( 
.A(n_7044),
.B(n_4458),
.Y(n_7634)
);

INVx2_ASAP7_75t_L g7635 ( 
.A(n_7020),
.Y(n_7635)
);

CKINVDCx5p33_ASAP7_75t_R g7636 ( 
.A(n_7054),
.Y(n_7636)
);

HB1xp67_ASAP7_75t_L g7637 ( 
.A(n_7063),
.Y(n_7637)
);

INVx2_ASAP7_75t_L g7638 ( 
.A(n_7022),
.Y(n_7638)
);

INVx3_ASAP7_75t_L g7639 ( 
.A(n_7023),
.Y(n_7639)
);

CKINVDCx5p33_ASAP7_75t_R g7640 ( 
.A(n_7074),
.Y(n_7640)
);

CKINVDCx11_ASAP7_75t_R g7641 ( 
.A(n_6975),
.Y(n_7641)
);

INVxp67_ASAP7_75t_L g7642 ( 
.A(n_7002),
.Y(n_7642)
);

INVx2_ASAP7_75t_L g7643 ( 
.A(n_7025),
.Y(n_7643)
);

INVx1_ASAP7_75t_L g7644 ( 
.A(n_6984),
.Y(n_7644)
);

AND2x2_ASAP7_75t_L g7645 ( 
.A(n_7010),
.B(n_4989),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_6994),
.Y(n_7646)
);

INVx2_ASAP7_75t_L g7647 ( 
.A(n_7034),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_6993),
.Y(n_7648)
);

CKINVDCx5p33_ASAP7_75t_R g7649 ( 
.A(n_7031),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_6876),
.Y(n_7650)
);

NAND2xp33_ASAP7_75t_L g7651 ( 
.A(n_7032),
.B(n_4460),
.Y(n_7651)
);

INVx3_ASAP7_75t_L g7652 ( 
.A(n_7061),
.Y(n_7652)
);

INVx1_ASAP7_75t_L g7653 ( 
.A(n_7000),
.Y(n_7653)
);

NAND2xp5_ASAP7_75t_SL g7654 ( 
.A(n_7356),
.B(n_7048),
.Y(n_7654)
);

INVx3_ASAP7_75t_L g7655 ( 
.A(n_7295),
.Y(n_7655)
);

CKINVDCx6p67_ASAP7_75t_R g7656 ( 
.A(n_7295),
.Y(n_7656)
);

BUFx6f_ASAP7_75t_L g7657 ( 
.A(n_7312),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7182),
.Y(n_7658)
);

NOR2xp33_ASAP7_75t_L g7659 ( 
.A(n_7443),
.B(n_6992),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_7193),
.Y(n_7660)
);

INVx2_ASAP7_75t_L g7661 ( 
.A(n_7110),
.Y(n_7661)
);

INVx1_ASAP7_75t_L g7662 ( 
.A(n_7197),
.Y(n_7662)
);

NOR2xp33_ASAP7_75t_L g7663 ( 
.A(n_7152),
.B(n_7629),
.Y(n_7663)
);

NOR2x1p5_ASAP7_75t_L g7664 ( 
.A(n_7094),
.B(n_4461),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_7200),
.Y(n_7665)
);

AO21x2_ASAP7_75t_L g7666 ( 
.A1(n_7624),
.A2(n_7069),
.B(n_7068),
.Y(n_7666)
);

INVx2_ASAP7_75t_L g7667 ( 
.A(n_7122),
.Y(n_7667)
);

NAND2xp33_ASAP7_75t_SL g7668 ( 
.A(n_7232),
.B(n_4462),
.Y(n_7668)
);

NAND2xp5_ASAP7_75t_SL g7669 ( 
.A(n_7212),
.B(n_6762),
.Y(n_7669)
);

INVx1_ASAP7_75t_L g7670 ( 
.A(n_7202),
.Y(n_7670)
);

BUFx10_ASAP7_75t_L g7671 ( 
.A(n_7274),
.Y(n_7671)
);

INVx3_ASAP7_75t_L g7672 ( 
.A(n_7097),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_7206),
.Y(n_7673)
);

NOR2xp33_ASAP7_75t_L g7674 ( 
.A(n_7562),
.B(n_6811),
.Y(n_7674)
);

NAND2xp5_ASAP7_75t_L g7675 ( 
.A(n_7544),
.B(n_6607),
.Y(n_7675)
);

INVx2_ASAP7_75t_L g7676 ( 
.A(n_7131),
.Y(n_7676)
);

INVx6_ASAP7_75t_L g7677 ( 
.A(n_7330),
.Y(n_7677)
);

INVx2_ASAP7_75t_L g7678 ( 
.A(n_7134),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_7214),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_7218),
.Y(n_7680)
);

INVxp67_ASAP7_75t_L g7681 ( 
.A(n_7137),
.Y(n_7681)
);

INVx2_ASAP7_75t_L g7682 ( 
.A(n_7138),
.Y(n_7682)
);

INVx1_ASAP7_75t_L g7683 ( 
.A(n_7219),
.Y(n_7683)
);

NOR2xp33_ASAP7_75t_SL g7684 ( 
.A(n_7208),
.B(n_5068),
.Y(n_7684)
);

INVx2_ASAP7_75t_L g7685 ( 
.A(n_7145),
.Y(n_7685)
);

AOI22xp5_ASAP7_75t_SL g7686 ( 
.A1(n_7502),
.A2(n_4465),
.B1(n_5008),
.B2(n_4410),
.Y(n_7686)
);

INVx3_ASAP7_75t_L g7687 ( 
.A(n_7097),
.Y(n_7687)
);

INVx2_ASAP7_75t_L g7688 ( 
.A(n_7146),
.Y(n_7688)
);

INVx2_ASAP7_75t_L g7689 ( 
.A(n_7148),
.Y(n_7689)
);

INVx2_ASAP7_75t_L g7690 ( 
.A(n_7174),
.Y(n_7690)
);

INVx3_ASAP7_75t_L g7691 ( 
.A(n_7102),
.Y(n_7691)
);

INVx5_ASAP7_75t_L g7692 ( 
.A(n_7415),
.Y(n_7692)
);

INVx1_ASAP7_75t_L g7693 ( 
.A(n_7221),
.Y(n_7693)
);

INVx2_ASAP7_75t_L g7694 ( 
.A(n_7187),
.Y(n_7694)
);

BUFx6f_ASAP7_75t_SL g7695 ( 
.A(n_7415),
.Y(n_7695)
);

NAND2xp5_ASAP7_75t_SL g7696 ( 
.A(n_7217),
.B(n_6677),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7223),
.Y(n_7697)
);

INVx2_ASAP7_75t_L g7698 ( 
.A(n_7196),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7225),
.Y(n_7699)
);

INVx2_ASAP7_75t_L g7700 ( 
.A(n_7201),
.Y(n_7700)
);

NOR2x1p5_ASAP7_75t_L g7701 ( 
.A(n_7103),
.B(n_4463),
.Y(n_7701)
);

INVx2_ASAP7_75t_L g7702 ( 
.A(n_7210),
.Y(n_7702)
);

INVx3_ASAP7_75t_L g7703 ( 
.A(n_7102),
.Y(n_7703)
);

INVx2_ASAP7_75t_L g7704 ( 
.A(n_7215),
.Y(n_7704)
);

INVx2_ASAP7_75t_L g7705 ( 
.A(n_7226),
.Y(n_7705)
);

INVx2_ASAP7_75t_L g7706 ( 
.A(n_7233),
.Y(n_7706)
);

NOR2xp33_ASAP7_75t_L g7707 ( 
.A(n_7608),
.B(n_6878),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_7242),
.Y(n_7708)
);

INVx1_ASAP7_75t_L g7709 ( 
.A(n_7244),
.Y(n_7709)
);

INVx1_ASAP7_75t_L g7710 ( 
.A(n_7258),
.Y(n_7710)
);

INVx1_ASAP7_75t_L g7711 ( 
.A(n_7265),
.Y(n_7711)
);

BUFx6f_ASAP7_75t_SL g7712 ( 
.A(n_7216),
.Y(n_7712)
);

INVx2_ASAP7_75t_L g7713 ( 
.A(n_7251),
.Y(n_7713)
);

INVx2_ASAP7_75t_L g7714 ( 
.A(n_7254),
.Y(n_7714)
);

NOR2xp33_ASAP7_75t_L g7715 ( 
.A(n_7420),
.B(n_7071),
.Y(n_7715)
);

INVx5_ASAP7_75t_L g7716 ( 
.A(n_7330),
.Y(n_7716)
);

AND2x2_ASAP7_75t_L g7717 ( 
.A(n_7421),
.B(n_5068),
.Y(n_7717)
);

AOI22xp5_ASAP7_75t_L g7718 ( 
.A1(n_7614),
.A2(n_7017),
.B1(n_6627),
.B2(n_7073),
.Y(n_7718)
);

INVx2_ASAP7_75t_L g7719 ( 
.A(n_7264),
.Y(n_7719)
);

NAND2xp5_ASAP7_75t_SL g7720 ( 
.A(n_7220),
.B(n_7084),
.Y(n_7720)
);

INVx3_ASAP7_75t_L g7721 ( 
.A(n_7205),
.Y(n_7721)
);

INVxp67_ASAP7_75t_SL g7722 ( 
.A(n_7580),
.Y(n_7722)
);

INVx2_ASAP7_75t_L g7723 ( 
.A(n_7271),
.Y(n_7723)
);

NAND2xp5_ASAP7_75t_L g7724 ( 
.A(n_7646),
.B(n_7088),
.Y(n_7724)
);

NAND3xp33_ASAP7_75t_L g7725 ( 
.A(n_7247),
.B(n_4466),
.C(n_4464),
.Y(n_7725)
);

INVx1_ASAP7_75t_L g7726 ( 
.A(n_7266),
.Y(n_7726)
);

BUFx2_ASAP7_75t_L g7727 ( 
.A(n_7098),
.Y(n_7727)
);

INVx2_ASAP7_75t_L g7728 ( 
.A(n_7280),
.Y(n_7728)
);

BUFx3_ASAP7_75t_L g7729 ( 
.A(n_7290),
.Y(n_7729)
);

AND2x2_ASAP7_75t_L g7730 ( 
.A(n_7114),
.B(n_7112),
.Y(n_7730)
);

INVx2_ASAP7_75t_L g7731 ( 
.A(n_7307),
.Y(n_7731)
);

NAND3xp33_ASAP7_75t_L g7732 ( 
.A(n_7260),
.B(n_4472),
.C(n_4467),
.Y(n_7732)
);

BUFx6f_ASAP7_75t_L g7733 ( 
.A(n_7159),
.Y(n_7733)
);

AOI22xp33_ASAP7_75t_L g7734 ( 
.A1(n_7468),
.A2(n_7591),
.B1(n_7532),
.B2(n_7493),
.Y(n_7734)
);

INVx2_ASAP7_75t_L g7735 ( 
.A(n_7324),
.Y(n_7735)
);

INVx3_ASAP7_75t_L g7736 ( 
.A(n_7282),
.Y(n_7736)
);

NAND2xp33_ASAP7_75t_L g7737 ( 
.A(n_7228),
.B(n_4473),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_7269),
.Y(n_7738)
);

INVx2_ASAP7_75t_L g7739 ( 
.A(n_7349),
.Y(n_7739)
);

NOR2xp33_ASAP7_75t_L g7740 ( 
.A(n_7561),
.B(n_4475),
.Y(n_7740)
);

BUFx10_ASAP7_75t_L g7741 ( 
.A(n_7113),
.Y(n_7741)
);

INVx1_ASAP7_75t_L g7742 ( 
.A(n_7272),
.Y(n_7742)
);

INVx1_ASAP7_75t_L g7743 ( 
.A(n_7277),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_7278),
.Y(n_7744)
);

INVx8_ASAP7_75t_L g7745 ( 
.A(n_7301),
.Y(n_7745)
);

INVx2_ASAP7_75t_L g7746 ( 
.A(n_7361),
.Y(n_7746)
);

INVx2_ASAP7_75t_L g7747 ( 
.A(n_7364),
.Y(n_7747)
);

NAND3xp33_ASAP7_75t_L g7748 ( 
.A(n_7328),
.B(n_4479),
.C(n_4476),
.Y(n_7748)
);

INVx2_ASAP7_75t_L g7749 ( 
.A(n_7366),
.Y(n_7749)
);

INVx2_ASAP7_75t_L g7750 ( 
.A(n_7373),
.Y(n_7750)
);

OR2x6_ASAP7_75t_L g7751 ( 
.A(n_7268),
.B(n_5018),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7283),
.Y(n_7752)
);

BUFx3_ASAP7_75t_L g7753 ( 
.A(n_7303),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_7285),
.Y(n_7754)
);

AND2x4_ASAP7_75t_L g7755 ( 
.A(n_7310),
.B(n_7178),
.Y(n_7755)
);

NAND2xp5_ASAP7_75t_SL g7756 ( 
.A(n_7649),
.B(n_4480),
.Y(n_7756)
);

NAND2xp5_ASAP7_75t_SL g7757 ( 
.A(n_7431),
.B(n_4481),
.Y(n_7757)
);

NAND2xp5_ASAP7_75t_L g7758 ( 
.A(n_7653),
.B(n_4864),
.Y(n_7758)
);

NAND2xp5_ASAP7_75t_SL g7759 ( 
.A(n_7115),
.B(n_4482),
.Y(n_7759)
);

INVx2_ASAP7_75t_L g7760 ( 
.A(n_7376),
.Y(n_7760)
);

INVx2_ASAP7_75t_L g7761 ( 
.A(n_7379),
.Y(n_7761)
);

AND2x2_ASAP7_75t_L g7762 ( 
.A(n_7326),
.B(n_5147),
.Y(n_7762)
);

INVx4_ASAP7_75t_L g7763 ( 
.A(n_7234),
.Y(n_7763)
);

INVx2_ASAP7_75t_L g7764 ( 
.A(n_7399),
.Y(n_7764)
);

NAND2xp5_ASAP7_75t_SL g7765 ( 
.A(n_7119),
.B(n_7120),
.Y(n_7765)
);

NAND2xp5_ASAP7_75t_L g7766 ( 
.A(n_7509),
.B(n_4873),
.Y(n_7766)
);

NOR2xp33_ASAP7_75t_L g7767 ( 
.A(n_7642),
.B(n_4484),
.Y(n_7767)
);

INVx1_ASAP7_75t_L g7768 ( 
.A(n_7289),
.Y(n_7768)
);

NAND2xp33_ASAP7_75t_L g7769 ( 
.A(n_7126),
.B(n_4486),
.Y(n_7769)
);

AO21x2_ASAP7_75t_L g7770 ( 
.A1(n_7626),
.A2(n_4889),
.B(n_4875),
.Y(n_7770)
);

OAI22xp33_ASAP7_75t_L g7771 ( 
.A1(n_7594),
.A2(n_7554),
.B1(n_7617),
.B2(n_7605),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_7291),
.Y(n_7772)
);

INVx2_ASAP7_75t_L g7773 ( 
.A(n_7402),
.Y(n_7773)
);

INVx3_ASAP7_75t_L g7774 ( 
.A(n_7235),
.Y(n_7774)
);

NAND2xp5_ASAP7_75t_L g7775 ( 
.A(n_7092),
.B(n_4891),
.Y(n_7775)
);

AND2x2_ASAP7_75t_L g7776 ( 
.A(n_7300),
.B(n_5147),
.Y(n_7776)
);

INVxp67_ASAP7_75t_SL g7777 ( 
.A(n_7580),
.Y(n_7777)
);

INVx2_ASAP7_75t_L g7778 ( 
.A(n_7417),
.Y(n_7778)
);

NAND2xp33_ASAP7_75t_L g7779 ( 
.A(n_7127),
.B(n_7129),
.Y(n_7779)
);

NAND3xp33_ASAP7_75t_L g7780 ( 
.A(n_7167),
.B(n_4490),
.C(n_4489),
.Y(n_7780)
);

INVx3_ASAP7_75t_L g7781 ( 
.A(n_7238),
.Y(n_7781)
);

INVx2_ASAP7_75t_L g7782 ( 
.A(n_7418),
.Y(n_7782)
);

NAND2xp5_ASAP7_75t_L g7783 ( 
.A(n_7252),
.B(n_7412),
.Y(n_7783)
);

INVx1_ASAP7_75t_L g7784 ( 
.A(n_7298),
.Y(n_7784)
);

INVx2_ASAP7_75t_SL g7785 ( 
.A(n_7546),
.Y(n_7785)
);

INVx3_ASAP7_75t_L g7786 ( 
.A(n_7257),
.Y(n_7786)
);

BUFx2_ASAP7_75t_L g7787 ( 
.A(n_7116),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7304),
.Y(n_7788)
);

NAND2xp33_ASAP7_75t_L g7789 ( 
.A(n_7132),
.B(n_7141),
.Y(n_7789)
);

INVx2_ASAP7_75t_SL g7790 ( 
.A(n_7173),
.Y(n_7790)
);

NAND2xp5_ASAP7_75t_SL g7791 ( 
.A(n_7445),
.B(n_4491),
.Y(n_7791)
);

NOR2xp33_ASAP7_75t_L g7792 ( 
.A(n_7250),
.B(n_4492),
.Y(n_7792)
);

INVx2_ASAP7_75t_L g7793 ( 
.A(n_7450),
.Y(n_7793)
);

AND2x2_ASAP7_75t_L g7794 ( 
.A(n_7231),
.B(n_5203),
.Y(n_7794)
);

INVx1_ASAP7_75t_L g7795 ( 
.A(n_7305),
.Y(n_7795)
);

AOI22xp5_ASAP7_75t_L g7796 ( 
.A1(n_7602),
.A2(n_4497),
.B1(n_4498),
.B2(n_4494),
.Y(n_7796)
);

INVx2_ASAP7_75t_L g7797 ( 
.A(n_7455),
.Y(n_7797)
);

BUFx3_ASAP7_75t_L g7798 ( 
.A(n_7248),
.Y(n_7798)
);

NAND2xp5_ASAP7_75t_L g7799 ( 
.A(n_7516),
.B(n_4892),
.Y(n_7799)
);

INVx1_ASAP7_75t_L g7800 ( 
.A(n_7308),
.Y(n_7800)
);

NAND2xp5_ASAP7_75t_L g7801 ( 
.A(n_7522),
.B(n_4893),
.Y(n_7801)
);

INVx2_ASAP7_75t_L g7802 ( 
.A(n_7506),
.Y(n_7802)
);

OR2x6_ASAP7_75t_L g7803 ( 
.A(n_7096),
.B(n_5218),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7309),
.Y(n_7804)
);

OR2x6_ASAP7_75t_L g7805 ( 
.A(n_7104),
.B(n_5485),
.Y(n_7805)
);

INVx1_ASAP7_75t_L g7806 ( 
.A(n_7311),
.Y(n_7806)
);

INVx2_ASAP7_75t_L g7807 ( 
.A(n_7095),
.Y(n_7807)
);

NAND2xp5_ASAP7_75t_SL g7808 ( 
.A(n_7229),
.B(n_4499),
.Y(n_7808)
);

BUFx10_ASAP7_75t_L g7809 ( 
.A(n_7162),
.Y(n_7809)
);

BUFx6f_ASAP7_75t_L g7810 ( 
.A(n_7117),
.Y(n_7810)
);

INVx1_ASAP7_75t_L g7811 ( 
.A(n_7318),
.Y(n_7811)
);

NAND2xp5_ASAP7_75t_L g7812 ( 
.A(n_7523),
.B(n_4899),
.Y(n_7812)
);

BUFx6f_ASAP7_75t_SL g7813 ( 
.A(n_7249),
.Y(n_7813)
);

BUFx6f_ASAP7_75t_L g7814 ( 
.A(n_7117),
.Y(n_7814)
);

NAND2xp5_ASAP7_75t_L g7815 ( 
.A(n_7572),
.B(n_4905),
.Y(n_7815)
);

NAND2xp33_ASAP7_75t_L g7816 ( 
.A(n_7156),
.B(n_4500),
.Y(n_7816)
);

NAND3xp33_ASAP7_75t_L g7817 ( 
.A(n_7484),
.B(n_4502),
.C(n_4501),
.Y(n_7817)
);

BUFx3_ASAP7_75t_L g7818 ( 
.A(n_7255),
.Y(n_7818)
);

NAND2xp5_ASAP7_75t_L g7819 ( 
.A(n_7320),
.B(n_7327),
.Y(n_7819)
);

NAND2xp5_ASAP7_75t_L g7820 ( 
.A(n_7332),
.B(n_7333),
.Y(n_7820)
);

INVx2_ASAP7_75t_L g7821 ( 
.A(n_7472),
.Y(n_7821)
);

INVx2_ASAP7_75t_L g7822 ( 
.A(n_7488),
.Y(n_7822)
);

INVx3_ASAP7_75t_L g7823 ( 
.A(n_7267),
.Y(n_7823)
);

NAND2xp5_ASAP7_75t_L g7824 ( 
.A(n_7335),
.B(n_4906),
.Y(n_7824)
);

INVx1_ASAP7_75t_L g7825 ( 
.A(n_7336),
.Y(n_7825)
);

INVx2_ASAP7_75t_L g7826 ( 
.A(n_7534),
.Y(n_7826)
);

INVx1_ASAP7_75t_L g7827 ( 
.A(n_7346),
.Y(n_7827)
);

BUFx3_ASAP7_75t_L g7828 ( 
.A(n_7263),
.Y(n_7828)
);

NAND2xp5_ASAP7_75t_L g7829 ( 
.A(n_7348),
.B(n_4915),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7352),
.Y(n_7830)
);

NOR3xp33_ASAP7_75t_L g7831 ( 
.A(n_7319),
.B(n_4922),
.C(n_4918),
.Y(n_7831)
);

INVx8_ASAP7_75t_L g7832 ( 
.A(n_7276),
.Y(n_7832)
);

INVx1_ASAP7_75t_L g7833 ( 
.A(n_7354),
.Y(n_7833)
);

INVx1_ASAP7_75t_L g7834 ( 
.A(n_7358),
.Y(n_7834)
);

NOR2xp33_ASAP7_75t_L g7835 ( 
.A(n_7158),
.B(n_4503),
.Y(n_7835)
);

INVx2_ASAP7_75t_L g7836 ( 
.A(n_7545),
.Y(n_7836)
);

INVx2_ASAP7_75t_L g7837 ( 
.A(n_7464),
.Y(n_7837)
);

INVx2_ASAP7_75t_L g7838 ( 
.A(n_7474),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7362),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7369),
.Y(n_7840)
);

INVx1_ASAP7_75t_L g7841 ( 
.A(n_7370),
.Y(n_7841)
);

INVx1_ASAP7_75t_L g7842 ( 
.A(n_7371),
.Y(n_7842)
);

INVx2_ASAP7_75t_SL g7843 ( 
.A(n_7125),
.Y(n_7843)
);

BUFx10_ASAP7_75t_L g7844 ( 
.A(n_7166),
.Y(n_7844)
);

NOR2xp33_ASAP7_75t_L g7845 ( 
.A(n_7582),
.B(n_4505),
.Y(n_7845)
);

INVx2_ASAP7_75t_L g7846 ( 
.A(n_7476),
.Y(n_7846)
);

INVx1_ASAP7_75t_L g7847 ( 
.A(n_7378),
.Y(n_7847)
);

INVx4_ASAP7_75t_L g7848 ( 
.A(n_7281),
.Y(n_7848)
);

INVx2_ASAP7_75t_L g7849 ( 
.A(n_7477),
.Y(n_7849)
);

INVx3_ASAP7_75t_L g7850 ( 
.A(n_7287),
.Y(n_7850)
);

INVx1_ASAP7_75t_L g7851 ( 
.A(n_7380),
.Y(n_7851)
);

INVx2_ASAP7_75t_L g7852 ( 
.A(n_7490),
.Y(n_7852)
);

INVx1_ASAP7_75t_L g7853 ( 
.A(n_7384),
.Y(n_7853)
);

NAND2xp5_ASAP7_75t_L g7854 ( 
.A(n_7388),
.B(n_7393),
.Y(n_7854)
);

INVx2_ASAP7_75t_L g7855 ( 
.A(n_7491),
.Y(n_7855)
);

INVx2_ASAP7_75t_L g7856 ( 
.A(n_7494),
.Y(n_7856)
);

INVx2_ASAP7_75t_L g7857 ( 
.A(n_7495),
.Y(n_7857)
);

BUFx6f_ASAP7_75t_L g7858 ( 
.A(n_7136),
.Y(n_7858)
);

NOR2xp33_ASAP7_75t_L g7859 ( 
.A(n_7599),
.B(n_4506),
.Y(n_7859)
);

NAND2xp5_ASAP7_75t_L g7860 ( 
.A(n_7398),
.B(n_4923),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_7403),
.Y(n_7861)
);

INVx1_ASAP7_75t_L g7862 ( 
.A(n_7406),
.Y(n_7862)
);

INVx2_ASAP7_75t_L g7863 ( 
.A(n_7100),
.Y(n_7863)
);

INVx2_ASAP7_75t_L g7864 ( 
.A(n_7105),
.Y(n_7864)
);

INVx2_ASAP7_75t_SL g7865 ( 
.A(n_7541),
.Y(n_7865)
);

INVxp67_ASAP7_75t_L g7866 ( 
.A(n_7147),
.Y(n_7866)
);

INVx2_ASAP7_75t_L g7867 ( 
.A(n_7106),
.Y(n_7867)
);

INVx4_ASAP7_75t_L g7868 ( 
.A(n_7293),
.Y(n_7868)
);

AND2x2_ASAP7_75t_L g7869 ( 
.A(n_7186),
.B(n_7645),
.Y(n_7869)
);

INVx2_ASAP7_75t_SL g7870 ( 
.A(n_7575),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_7407),
.Y(n_7871)
);

INVx1_ASAP7_75t_L g7872 ( 
.A(n_7410),
.Y(n_7872)
);

INVx8_ASAP7_75t_L g7873 ( 
.A(n_7279),
.Y(n_7873)
);

INVx8_ASAP7_75t_L g7874 ( 
.A(n_7296),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_7411),
.Y(n_7875)
);

CKINVDCx5p33_ASAP7_75t_R g7876 ( 
.A(n_7337),
.Y(n_7876)
);

NAND2xp5_ASAP7_75t_L g7877 ( 
.A(n_7413),
.B(n_4925),
.Y(n_7877)
);

INVx3_ASAP7_75t_L g7878 ( 
.A(n_7306),
.Y(n_7878)
);

INVx1_ASAP7_75t_L g7879 ( 
.A(n_7419),
.Y(n_7879)
);

NOR2xp33_ASAP7_75t_L g7880 ( 
.A(n_7387),
.B(n_4508),
.Y(n_7880)
);

INVx2_ASAP7_75t_L g7881 ( 
.A(n_7107),
.Y(n_7881)
);

INVx2_ASAP7_75t_L g7882 ( 
.A(n_7108),
.Y(n_7882)
);

NAND2xp5_ASAP7_75t_L g7883 ( 
.A(n_7429),
.B(n_4926),
.Y(n_7883)
);

NAND2xp5_ASAP7_75t_SL g7884 ( 
.A(n_7259),
.B(n_4511),
.Y(n_7884)
);

NAND3xp33_ASAP7_75t_L g7885 ( 
.A(n_7237),
.B(n_4515),
.C(n_4513),
.Y(n_7885)
);

INVx2_ASAP7_75t_L g7886 ( 
.A(n_7118),
.Y(n_7886)
);

INVx8_ASAP7_75t_L g7887 ( 
.A(n_7313),
.Y(n_7887)
);

INVx2_ASAP7_75t_L g7888 ( 
.A(n_7121),
.Y(n_7888)
);

NAND2xp5_ASAP7_75t_SL g7889 ( 
.A(n_7487),
.B(n_4516),
.Y(n_7889)
);

INVx2_ASAP7_75t_L g7890 ( 
.A(n_7128),
.Y(n_7890)
);

AND2x2_ASAP7_75t_L g7891 ( 
.A(n_7157),
.B(n_5203),
.Y(n_7891)
);

OAI22xp33_ASAP7_75t_L g7892 ( 
.A1(n_7609),
.A2(n_4519),
.B1(n_4520),
.B2(n_4518),
.Y(n_7892)
);

NAND2xp5_ASAP7_75t_SL g7893 ( 
.A(n_7363),
.B(n_4522),
.Y(n_7893)
);

OAI22xp33_ASAP7_75t_L g7894 ( 
.A1(n_7600),
.A2(n_4524),
.B1(n_4527),
.B2(n_4523),
.Y(n_7894)
);

NAND2xp5_ASAP7_75t_SL g7895 ( 
.A(n_7368),
.B(n_4528),
.Y(n_7895)
);

NAND2xp5_ASAP7_75t_SL g7896 ( 
.A(n_7381),
.B(n_4529),
.Y(n_7896)
);

INVx2_ASAP7_75t_L g7897 ( 
.A(n_7133),
.Y(n_7897)
);

NAND2xp5_ASAP7_75t_L g7898 ( 
.A(n_7432),
.B(n_4927),
.Y(n_7898)
);

INVx2_ASAP7_75t_L g7899 ( 
.A(n_7139),
.Y(n_7899)
);

INVx2_ASAP7_75t_L g7900 ( 
.A(n_7144),
.Y(n_7900)
);

INVx1_ASAP7_75t_L g7901 ( 
.A(n_7435),
.Y(n_7901)
);

NAND2xp5_ASAP7_75t_SL g7902 ( 
.A(n_7382),
.B(n_7385),
.Y(n_7902)
);

INVx1_ASAP7_75t_L g7903 ( 
.A(n_7444),
.Y(n_7903)
);

INVx5_ASAP7_75t_L g7904 ( 
.A(n_7245),
.Y(n_7904)
);

BUFx10_ASAP7_75t_L g7905 ( 
.A(n_7170),
.Y(n_7905)
);

OAI22xp33_ASAP7_75t_SL g7906 ( 
.A1(n_7622),
.A2(n_7451),
.B1(n_7457),
.B2(n_7448),
.Y(n_7906)
);

NAND2xp5_ASAP7_75t_SL g7907 ( 
.A(n_7389),
.B(n_4531),
.Y(n_7907)
);

INVxp33_ASAP7_75t_L g7908 ( 
.A(n_7111),
.Y(n_7908)
);

BUFx6f_ASAP7_75t_L g7909 ( 
.A(n_7136),
.Y(n_7909)
);

NOR2x1p5_ASAP7_75t_L g7910 ( 
.A(n_7171),
.B(n_4532),
.Y(n_7910)
);

INVx1_ASAP7_75t_SL g7911 ( 
.A(n_7195),
.Y(n_7911)
);

AND2x2_ASAP7_75t_L g7912 ( 
.A(n_7527),
.B(n_7481),
.Y(n_7912)
);

INVx2_ASAP7_75t_L g7913 ( 
.A(n_7150),
.Y(n_7913)
);

INVx2_ASAP7_75t_L g7914 ( 
.A(n_7153),
.Y(n_7914)
);

NAND2xp5_ASAP7_75t_L g7915 ( 
.A(n_7447),
.B(n_4939),
.Y(n_7915)
);

NAND2xp5_ASAP7_75t_SL g7916 ( 
.A(n_7390),
.B(n_4533),
.Y(n_7916)
);

NOR2xp33_ASAP7_75t_L g7917 ( 
.A(n_7559),
.B(n_4536),
.Y(n_7917)
);

AND2x6_ASAP7_75t_L g7918 ( 
.A(n_7650),
.B(n_4940),
.Y(n_7918)
);

NOR2xp33_ASAP7_75t_L g7919 ( 
.A(n_7239),
.B(n_4537),
.Y(n_7919)
);

INVx3_ASAP7_75t_L g7920 ( 
.A(n_7316),
.Y(n_7920)
);

INVx2_ASAP7_75t_L g7921 ( 
.A(n_7154),
.Y(n_7921)
);

INVx1_ASAP7_75t_L g7922 ( 
.A(n_7452),
.Y(n_7922)
);

NAND2xp5_ASAP7_75t_SL g7923 ( 
.A(n_7392),
.B(n_4538),
.Y(n_7923)
);

NAND2xp5_ASAP7_75t_SL g7924 ( 
.A(n_7395),
.B(n_4541),
.Y(n_7924)
);

INVx2_ASAP7_75t_L g7925 ( 
.A(n_7160),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_7454),
.Y(n_7926)
);

INVx5_ASAP7_75t_L g7927 ( 
.A(n_7537),
.Y(n_7927)
);

CKINVDCx5p33_ASAP7_75t_R g7928 ( 
.A(n_7230),
.Y(n_7928)
);

INVxp33_ASAP7_75t_L g7929 ( 
.A(n_7246),
.Y(n_7929)
);

INVx2_ASAP7_75t_L g7930 ( 
.A(n_7161),
.Y(n_7930)
);

INVx2_ASAP7_75t_L g7931 ( 
.A(n_7164),
.Y(n_7931)
);

INVx2_ASAP7_75t_L g7932 ( 
.A(n_7165),
.Y(n_7932)
);

NAND2xp33_ASAP7_75t_SL g7933 ( 
.A(n_7357),
.B(n_4542),
.Y(n_7933)
);

INVx1_ASAP7_75t_L g7934 ( 
.A(n_7456),
.Y(n_7934)
);

BUFx10_ASAP7_75t_L g7935 ( 
.A(n_7172),
.Y(n_7935)
);

INVx3_ASAP7_75t_L g7936 ( 
.A(n_7321),
.Y(n_7936)
);

AOI22xp33_ASAP7_75t_L g7937 ( 
.A1(n_7555),
.A2(n_5223),
.B1(n_5233),
.B2(n_5217),
.Y(n_7937)
);

INVx2_ASAP7_75t_L g7938 ( 
.A(n_7168),
.Y(n_7938)
);

INVx1_ASAP7_75t_L g7939 ( 
.A(n_7459),
.Y(n_7939)
);

INVx1_ASAP7_75t_L g7940 ( 
.A(n_7513),
.Y(n_7940)
);

NAND3xp33_ASAP7_75t_L g7941 ( 
.A(n_7198),
.B(n_4545),
.C(n_4544),
.Y(n_7941)
);

INVx2_ASAP7_75t_L g7942 ( 
.A(n_7175),
.Y(n_7942)
);

NAND3xp33_ASAP7_75t_L g7943 ( 
.A(n_7615),
.B(n_4547),
.C(n_4546),
.Y(n_7943)
);

NAND2xp5_ASAP7_75t_L g7944 ( 
.A(n_7514),
.B(n_4945),
.Y(n_7944)
);

INVx2_ASAP7_75t_L g7945 ( 
.A(n_7181),
.Y(n_7945)
);

INVx2_ASAP7_75t_L g7946 ( 
.A(n_7567),
.Y(n_7946)
);

NAND2xp5_ASAP7_75t_L g7947 ( 
.A(n_7515),
.B(n_4946),
.Y(n_7947)
);

INVx4_ASAP7_75t_L g7948 ( 
.A(n_7323),
.Y(n_7948)
);

NAND2xp5_ASAP7_75t_L g7949 ( 
.A(n_7518),
.B(n_7521),
.Y(n_7949)
);

INVx2_ASAP7_75t_SL g7950 ( 
.A(n_7575),
.Y(n_7950)
);

INVx2_ASAP7_75t_L g7951 ( 
.A(n_7583),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7525),
.Y(n_7952)
);

NAND2xp5_ASAP7_75t_SL g7953 ( 
.A(n_7473),
.B(n_4554),
.Y(n_7953)
);

OAI22xp5_ASAP7_75t_L g7954 ( 
.A1(n_7529),
.A2(n_4561),
.B1(n_4563),
.B2(n_4560),
.Y(n_7954)
);

NAND2xp5_ASAP7_75t_SL g7955 ( 
.A(n_7586),
.B(n_7579),
.Y(n_7955)
);

INVx1_ASAP7_75t_L g7956 ( 
.A(n_7530),
.Y(n_7956)
);

INVx2_ASAP7_75t_L g7957 ( 
.A(n_7589),
.Y(n_7957)
);

BUFx6f_ASAP7_75t_L g7958 ( 
.A(n_7190),
.Y(n_7958)
);

BUFx2_ASAP7_75t_L g7959 ( 
.A(n_7331),
.Y(n_7959)
);

INVx2_ASAP7_75t_L g7960 ( 
.A(n_7593),
.Y(n_7960)
);

INVx3_ASAP7_75t_L g7961 ( 
.A(n_7325),
.Y(n_7961)
);

INVx2_ASAP7_75t_L g7962 ( 
.A(n_7606),
.Y(n_7962)
);

INVx1_ASAP7_75t_L g7963 ( 
.A(n_7531),
.Y(n_7963)
);

NAND2xp5_ASAP7_75t_SL g7964 ( 
.A(n_7586),
.B(n_4565),
.Y(n_7964)
);

INVx1_ASAP7_75t_L g7965 ( 
.A(n_7613),
.Y(n_7965)
);

NAND2xp5_ASAP7_75t_SL g7966 ( 
.A(n_7504),
.B(n_4566),
.Y(n_7966)
);

INVx2_ASAP7_75t_L g7967 ( 
.A(n_7623),
.Y(n_7967)
);

INVx2_ASAP7_75t_L g7968 ( 
.A(n_7635),
.Y(n_7968)
);

OR2x6_ASAP7_75t_L g7969 ( 
.A(n_7619),
.B(n_4760),
.Y(n_7969)
);

NAND2xp5_ASAP7_75t_SL g7970 ( 
.A(n_7508),
.B(n_4572),
.Y(n_7970)
);

OAI22xp33_ASAP7_75t_L g7971 ( 
.A1(n_7262),
.A2(n_4576),
.B1(n_4582),
.B2(n_4574),
.Y(n_7971)
);

INVx1_ASAP7_75t_L g7972 ( 
.A(n_7638),
.Y(n_7972)
);

INVx2_ASAP7_75t_L g7973 ( 
.A(n_7643),
.Y(n_7973)
);

NAND2xp5_ASAP7_75t_L g7974 ( 
.A(n_7517),
.B(n_4947),
.Y(n_7974)
);

NAND2xp5_ASAP7_75t_L g7975 ( 
.A(n_7520),
.B(n_4961),
.Y(n_7975)
);

NAND3xp33_ASAP7_75t_L g7976 ( 
.A(n_7093),
.B(n_4586),
.C(n_4584),
.Y(n_7976)
);

CKINVDCx5p33_ASAP7_75t_R g7977 ( 
.A(n_7179),
.Y(n_7977)
);

BUFx6f_ASAP7_75t_L g7978 ( 
.A(n_7190),
.Y(n_7978)
);

INVx2_ASAP7_75t_L g7979 ( 
.A(n_7647),
.Y(n_7979)
);

NAND2xp5_ASAP7_75t_SL g7980 ( 
.A(n_7207),
.B(n_4589),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_SL g7981 ( 
.A(n_7441),
.B(n_4592),
.Y(n_7981)
);

INVx2_ASAP7_75t_L g7982 ( 
.A(n_7588),
.Y(n_7982)
);

INVx1_ASAP7_75t_SL g7983 ( 
.A(n_7341),
.Y(n_7983)
);

NAND2xp5_ASAP7_75t_L g7984 ( 
.A(n_7374),
.B(n_4964),
.Y(n_7984)
);

BUFx6f_ASAP7_75t_L g7985 ( 
.A(n_7191),
.Y(n_7985)
);

NAND2xp5_ASAP7_75t_SL g7986 ( 
.A(n_7441),
.B(n_7486),
.Y(n_7986)
);

INVx2_ASAP7_75t_L g7987 ( 
.A(n_7588),
.Y(n_7987)
);

NOR2xp33_ASAP7_75t_SL g7988 ( 
.A(n_7185),
.B(n_5217),
.Y(n_7988)
);

INVx2_ASAP7_75t_L g7989 ( 
.A(n_7612),
.Y(n_7989)
);

INVx2_ASAP7_75t_L g7990 ( 
.A(n_7612),
.Y(n_7990)
);

NAND2xp5_ASAP7_75t_SL g7991 ( 
.A(n_7486),
.B(n_4594),
.Y(n_7991)
);

NAND2xp5_ASAP7_75t_L g7992 ( 
.A(n_7553),
.B(n_4968),
.Y(n_7992)
);

INVx2_ASAP7_75t_L g7993 ( 
.A(n_7497),
.Y(n_7993)
);

BUFx2_ASAP7_75t_L g7994 ( 
.A(n_7355),
.Y(n_7994)
);

INVx2_ASAP7_75t_L g7995 ( 
.A(n_7639),
.Y(n_7995)
);

INVx1_ASAP7_75t_L g7996 ( 
.A(n_7632),
.Y(n_7996)
);

INVx2_ASAP7_75t_SL g7997 ( 
.A(n_7334),
.Y(n_7997)
);

NAND2xp5_ASAP7_75t_L g7998 ( 
.A(n_7644),
.B(n_4973),
.Y(n_7998)
);

CKINVDCx5p33_ASAP7_75t_R g7999 ( 
.A(n_7194),
.Y(n_7999)
);

NAND2xp5_ASAP7_75t_SL g8000 ( 
.A(n_7339),
.B(n_4595),
.Y(n_8000)
);

AND2x2_ASAP7_75t_L g8001 ( 
.A(n_7618),
.B(n_5223),
.Y(n_8001)
);

NOR2xp33_ASAP7_75t_L g8002 ( 
.A(n_7101),
.B(n_4596),
.Y(n_8002)
);

INVx1_ASAP7_75t_L g8003 ( 
.A(n_7633),
.Y(n_8003)
);

INVx2_ASAP7_75t_L g8004 ( 
.A(n_7652),
.Y(n_8004)
);

OAI21xp33_ASAP7_75t_L g8005 ( 
.A1(n_7628),
.A2(n_4605),
.B(n_4597),
.Y(n_8005)
);

INVx2_ASAP7_75t_L g8006 ( 
.A(n_7627),
.Y(n_8006)
);

INVx1_ASAP7_75t_SL g8007 ( 
.A(n_7360),
.Y(n_8007)
);

INVx2_ASAP7_75t_L g8008 ( 
.A(n_7630),
.Y(n_8008)
);

INVx1_ASAP7_75t_L g8009 ( 
.A(n_7648),
.Y(n_8009)
);

INVx1_ASAP7_75t_L g8010 ( 
.A(n_7510),
.Y(n_8010)
);

INVx2_ASAP7_75t_L g8011 ( 
.A(n_7453),
.Y(n_8011)
);

INVx1_ASAP7_75t_L g8012 ( 
.A(n_7533),
.Y(n_8012)
);

AND2x2_ASAP7_75t_L g8013 ( 
.A(n_7463),
.B(n_5233),
.Y(n_8013)
);

INVx2_ASAP7_75t_L g8014 ( 
.A(n_7564),
.Y(n_8014)
);

AO21x2_ASAP7_75t_L g8015 ( 
.A1(n_7099),
.A2(n_4982),
.B(n_4979),
.Y(n_8015)
);

INVx2_ASAP7_75t_L g8016 ( 
.A(n_7607),
.Y(n_8016)
);

INVx1_ASAP7_75t_L g8017 ( 
.A(n_7590),
.Y(n_8017)
);

NAND2xp33_ASAP7_75t_L g8018 ( 
.A(n_7397),
.B(n_4606),
.Y(n_8018)
);

AND2x6_ASAP7_75t_L g8019 ( 
.A(n_7536),
.B(n_4994),
.Y(n_8019)
);

INVx1_ASAP7_75t_L g8020 ( 
.A(n_7542),
.Y(n_8020)
);

INVx2_ASAP7_75t_L g8021 ( 
.A(n_7109),
.Y(n_8021)
);

NAND2xp33_ASAP7_75t_SL g8022 ( 
.A(n_7169),
.B(n_4607),
.Y(n_8022)
);

NAND2xp5_ASAP7_75t_L g8023 ( 
.A(n_7501),
.B(n_4996),
.Y(n_8023)
);

NAND2xp5_ASAP7_75t_L g8024 ( 
.A(n_7135),
.B(n_4999),
.Y(n_8024)
);

NAND2xp5_ASAP7_75t_SL g8025 ( 
.A(n_7343),
.B(n_4608),
.Y(n_8025)
);

INVx2_ASAP7_75t_L g8026 ( 
.A(n_7236),
.Y(n_8026)
);

NOR2xp33_ASAP7_75t_L g8027 ( 
.A(n_7130),
.B(n_4609),
.Y(n_8027)
);

NAND2xp5_ASAP7_75t_SL g8028 ( 
.A(n_7344),
.B(n_4610),
.Y(n_8028)
);

INVx2_ASAP7_75t_L g8029 ( 
.A(n_7430),
.Y(n_8029)
);

INVx2_ASAP7_75t_L g8030 ( 
.A(n_7552),
.Y(n_8030)
);

INVx2_ASAP7_75t_L g8031 ( 
.A(n_7556),
.Y(n_8031)
);

NAND3xp33_ASAP7_75t_L g8032 ( 
.A(n_7375),
.B(n_4620),
.C(n_4618),
.Y(n_8032)
);

INVx2_ASAP7_75t_L g8033 ( 
.A(n_7557),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_7563),
.Y(n_8034)
);

OAI22xp5_ASAP7_75t_L g8035 ( 
.A1(n_7560),
.A2(n_4623),
.B1(n_4627),
.B2(n_4621),
.Y(n_8035)
);

INVx5_ASAP7_75t_L g8036 ( 
.A(n_7191),
.Y(n_8036)
);

INVx3_ASAP7_75t_L g8037 ( 
.A(n_7347),
.Y(n_8037)
);

NAND2xp5_ASAP7_75t_SL g8038 ( 
.A(n_7350),
.B(n_7351),
.Y(n_8038)
);

INVx2_ASAP7_75t_L g8039 ( 
.A(n_7571),
.Y(n_8039)
);

INVx3_ASAP7_75t_L g8040 ( 
.A(n_7204),
.Y(n_8040)
);

INVx2_ASAP7_75t_L g8041 ( 
.A(n_7581),
.Y(n_8041)
);

INVx1_ASAP7_75t_L g8042 ( 
.A(n_7584),
.Y(n_8042)
);

NAND2xp33_ASAP7_75t_L g8043 ( 
.A(n_7540),
.B(n_4630),
.Y(n_8043)
);

INVx1_ASAP7_75t_L g8044 ( 
.A(n_7587),
.Y(n_8044)
);

NAND2xp5_ASAP7_75t_L g8045 ( 
.A(n_7601),
.B(n_5003),
.Y(n_8045)
);

INVx2_ASAP7_75t_L g8046 ( 
.A(n_7596),
.Y(n_8046)
);

INVx2_ASAP7_75t_L g8047 ( 
.A(n_7597),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_7604),
.Y(n_8048)
);

NAND2xp5_ASAP7_75t_SL g8049 ( 
.A(n_7286),
.B(n_4632),
.Y(n_8049)
);

NAND2xp5_ASAP7_75t_L g8050 ( 
.A(n_7123),
.B(n_5010),
.Y(n_8050)
);

NAND2xp5_ASAP7_75t_L g8051 ( 
.A(n_7314),
.B(n_7253),
.Y(n_8051)
);

NAND2xp5_ASAP7_75t_L g8052 ( 
.A(n_7314),
.B(n_5021),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_7611),
.Y(n_8053)
);

INVx1_ASAP7_75t_L g8054 ( 
.A(n_7616),
.Y(n_8054)
);

INVx2_ASAP7_75t_L g8055 ( 
.A(n_7140),
.Y(n_8055)
);

INVx2_ASAP7_75t_L g8056 ( 
.A(n_7496),
.Y(n_8056)
);

INVx1_ASAP7_75t_L g8057 ( 
.A(n_7261),
.Y(n_8057)
);

OR2x2_ASAP7_75t_L g8058 ( 
.A(n_7329),
.B(n_5024),
.Y(n_8058)
);

INVx2_ASAP7_75t_L g8059 ( 
.A(n_7496),
.Y(n_8059)
);

INVx2_ASAP7_75t_L g8060 ( 
.A(n_7519),
.Y(n_8060)
);

INVx2_ASAP7_75t_L g8061 ( 
.A(n_7519),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_SL g8062 ( 
.A(n_7317),
.B(n_4633),
.Y(n_8062)
);

AOI21x1_ASAP7_75t_L g8063 ( 
.A1(n_7405),
.A2(n_5031),
.B(n_5029),
.Y(n_8063)
);

INVxp67_ASAP7_75t_L g8064 ( 
.A(n_7585),
.Y(n_8064)
);

INVx1_ASAP7_75t_SL g8065 ( 
.A(n_7365),
.Y(n_8065)
);

CKINVDCx5p33_ASAP7_75t_R g8066 ( 
.A(n_7199),
.Y(n_8066)
);

INVx2_ASAP7_75t_L g8067 ( 
.A(n_7526),
.Y(n_8067)
);

INVx2_ASAP7_75t_L g8068 ( 
.A(n_7526),
.Y(n_8068)
);

INVx2_ASAP7_75t_L g8069 ( 
.A(n_7539),
.Y(n_8069)
);

NAND2xp33_ASAP7_75t_L g8070 ( 
.A(n_7543),
.B(n_4636),
.Y(n_8070)
);

INVx2_ASAP7_75t_L g8071 ( 
.A(n_7539),
.Y(n_8071)
);

AND2x2_ASAP7_75t_L g8072 ( 
.A(n_7479),
.B(n_5272),
.Y(n_8072)
);

NAND2xp5_ASAP7_75t_SL g8073 ( 
.A(n_7270),
.B(n_4642),
.Y(n_8073)
);

INVx2_ASAP7_75t_L g8074 ( 
.A(n_7549),
.Y(n_8074)
);

INVx2_ASAP7_75t_L g8075 ( 
.A(n_7549),
.Y(n_8075)
);

INVx2_ASAP7_75t_L g8076 ( 
.A(n_7558),
.Y(n_8076)
);

NAND2xp5_ASAP7_75t_SL g8077 ( 
.A(n_7338),
.B(n_4644),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_7273),
.Y(n_8078)
);

INVx2_ASAP7_75t_L g8079 ( 
.A(n_7558),
.Y(n_8079)
);

NAND2xp5_ASAP7_75t_L g8080 ( 
.A(n_7314),
.B(n_5045),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_7292),
.Y(n_8081)
);

BUFx6f_ASAP7_75t_L g8082 ( 
.A(n_7204),
.Y(n_8082)
);

NOR2xp33_ASAP7_75t_L g8083 ( 
.A(n_7284),
.B(n_4646),
.Y(n_8083)
);

INVxp67_ASAP7_75t_L g8084 ( 
.A(n_7180),
.Y(n_8084)
);

NOR2xp33_ASAP7_75t_L g8085 ( 
.A(n_7595),
.B(n_4647),
.Y(n_8085)
);

NAND2xp5_ASAP7_75t_SL g8086 ( 
.A(n_7353),
.B(n_4649),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_7299),
.Y(n_8087)
);

INVx2_ASAP7_75t_L g8088 ( 
.A(n_7565),
.Y(n_8088)
);

INVx2_ASAP7_75t_L g8089 ( 
.A(n_7565),
.Y(n_8089)
);

INVx2_ASAP7_75t_L g8090 ( 
.A(n_7573),
.Y(n_8090)
);

NAND2xp5_ASAP7_75t_L g8091 ( 
.A(n_7383),
.B(n_5046),
.Y(n_8091)
);

INVx2_ASAP7_75t_L g8092 ( 
.A(n_7573),
.Y(n_8092)
);

INVx4_ASAP7_75t_L g8093 ( 
.A(n_7401),
.Y(n_8093)
);

OR2x6_ASAP7_75t_L g8094 ( 
.A(n_7439),
.B(n_4790),
.Y(n_8094)
);

AND2x2_ASAP7_75t_L g8095 ( 
.A(n_7485),
.B(n_5272),
.Y(n_8095)
);

BUFx6f_ASAP7_75t_L g8096 ( 
.A(n_7209),
.Y(n_8096)
);

AND2x2_ASAP7_75t_SL g8097 ( 
.A(n_7631),
.B(n_4813),
.Y(n_8097)
);

INVx2_ASAP7_75t_L g8098 ( 
.A(n_7416),
.Y(n_8098)
);

INVx1_ASAP7_75t_L g8099 ( 
.A(n_7391),
.Y(n_8099)
);

INVx2_ASAP7_75t_L g8100 ( 
.A(n_7416),
.Y(n_8100)
);

NAND2xp5_ASAP7_75t_SL g8101 ( 
.A(n_7404),
.B(n_4650),
.Y(n_8101)
);

NAND2xp33_ASAP7_75t_L g8102 ( 
.A(n_7422),
.B(n_4651),
.Y(n_8102)
);

INVx2_ASAP7_75t_L g8103 ( 
.A(n_7424),
.Y(n_8103)
);

AO22x2_ASAP7_75t_L g8104 ( 
.A1(n_7302),
.A2(n_5062),
.B1(n_5072),
.B2(n_5051),
.Y(n_8104)
);

NAND2xp5_ASAP7_75t_SL g8105 ( 
.A(n_7428),
.B(n_4652),
.Y(n_8105)
);

INVx2_ASAP7_75t_L g8106 ( 
.A(n_7424),
.Y(n_8106)
);

NAND2xp5_ASAP7_75t_L g8107 ( 
.A(n_7394),
.B(n_5076),
.Y(n_8107)
);

BUFx6f_ASAP7_75t_L g8108 ( 
.A(n_7209),
.Y(n_8108)
);

INVx2_ASAP7_75t_L g8109 ( 
.A(n_7449),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_7396),
.Y(n_8110)
);

NAND2xp5_ASAP7_75t_L g8111 ( 
.A(n_7409),
.B(n_5082),
.Y(n_8111)
);

INVx2_ASAP7_75t_L g8112 ( 
.A(n_7458),
.Y(n_8112)
);

INVx2_ASAP7_75t_L g8113 ( 
.A(n_7466),
.Y(n_8113)
);

AOI21x1_ASAP7_75t_L g8114 ( 
.A1(n_7434),
.A2(n_7475),
.B(n_7442),
.Y(n_8114)
);

NAND2xp5_ASAP7_75t_SL g8115 ( 
.A(n_7574),
.B(n_4653),
.Y(n_8115)
);

BUFx3_ASAP7_75t_L g8116 ( 
.A(n_7211),
.Y(n_8116)
);

INVx2_ASAP7_75t_L g8117 ( 
.A(n_7499),
.Y(n_8117)
);

INVx2_ASAP7_75t_L g8118 ( 
.A(n_7551),
.Y(n_8118)
);

INVx5_ASAP7_75t_L g8119 ( 
.A(n_7211),
.Y(n_8119)
);

INVx1_ASAP7_75t_L g8120 ( 
.A(n_7480),
.Y(n_8120)
);

NAND2xp5_ASAP7_75t_L g8121 ( 
.A(n_7492),
.B(n_5089),
.Y(n_8121)
);

INVx4_ASAP7_75t_L g8122 ( 
.A(n_7408),
.Y(n_8122)
);

INVx1_ASAP7_75t_L g8123 ( 
.A(n_7498),
.Y(n_8123)
);

INVx2_ASAP7_75t_L g8124 ( 
.A(n_7577),
.Y(n_8124)
);

NAND2xp5_ASAP7_75t_SL g8125 ( 
.A(n_7574),
.B(n_4656),
.Y(n_8125)
);

INVx1_ASAP7_75t_L g8126 ( 
.A(n_7446),
.Y(n_8126)
);

INVx1_ASAP7_75t_SL g8127 ( 
.A(n_7367),
.Y(n_8127)
);

NAND2xp5_ASAP7_75t_L g8128 ( 
.A(n_7592),
.B(n_5095),
.Y(n_8128)
);

INVx4_ASAP7_75t_L g8129 ( 
.A(n_7414),
.Y(n_8129)
);

INVx1_ASAP7_75t_L g8130 ( 
.A(n_7576),
.Y(n_8130)
);

BUFx6f_ASAP7_75t_L g8131 ( 
.A(n_7213),
.Y(n_8131)
);

NAND2xp5_ASAP7_75t_SL g8132 ( 
.A(n_7636),
.B(n_4660),
.Y(n_8132)
);

INVx2_ASAP7_75t_L g8133 ( 
.A(n_7294),
.Y(n_8133)
);

OAI21xp33_ASAP7_75t_SL g8134 ( 
.A1(n_7535),
.A2(n_5097),
.B(n_5096),
.Y(n_8134)
);

INVx2_ASAP7_75t_L g8135 ( 
.A(n_7294),
.Y(n_8135)
);

NAND3xp33_ASAP7_75t_L g8136 ( 
.A(n_7538),
.B(n_4662),
.C(n_4661),
.Y(n_8136)
);

NAND2xp5_ASAP7_75t_SL g8137 ( 
.A(n_7640),
.B(n_7461),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_7297),
.Y(n_8138)
);

NOR2x1p5_ASAP7_75t_L g8139 ( 
.A(n_7124),
.B(n_4664),
.Y(n_8139)
);

INVx1_ASAP7_75t_L g8140 ( 
.A(n_7651),
.Y(n_8140)
);

INVx2_ASAP7_75t_L g8141 ( 
.A(n_7297),
.Y(n_8141)
);

INVx1_ASAP7_75t_L g8142 ( 
.A(n_7637),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_7547),
.Y(n_8143)
);

INVx3_ASAP7_75t_L g8144 ( 
.A(n_7213),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_7467),
.Y(n_8145)
);

INVx2_ASAP7_75t_L g8146 ( 
.A(n_7322),
.Y(n_8146)
);

INVx2_ASAP7_75t_SL g8147 ( 
.A(n_7372),
.Y(n_8147)
);

NAND3xp33_ASAP7_75t_L g8148 ( 
.A(n_7340),
.B(n_4666),
.C(n_4665),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7483),
.Y(n_8149)
);

INVx2_ASAP7_75t_L g8150 ( 
.A(n_7322),
.Y(n_8150)
);

INVx2_ASAP7_75t_SL g8151 ( 
.A(n_7377),
.Y(n_8151)
);

INVx2_ASAP7_75t_L g8152 ( 
.A(n_7224),
.Y(n_8152)
);

INVx2_ASAP7_75t_L g8153 ( 
.A(n_7224),
.Y(n_8153)
);

NOR2xp33_ASAP7_75t_L g8154 ( 
.A(n_7548),
.B(n_4671),
.Y(n_8154)
);

NAND2xp5_ASAP7_75t_SL g8155 ( 
.A(n_7345),
.B(n_4673),
.Y(n_8155)
);

INVx1_ASAP7_75t_L g8156 ( 
.A(n_7500),
.Y(n_8156)
);

AOI21x1_ASAP7_75t_L g8157 ( 
.A1(n_7149),
.A2(n_5104),
.B(n_5102),
.Y(n_8157)
);

INVx2_ASAP7_75t_SL g8158 ( 
.A(n_7240),
.Y(n_8158)
);

NAND2xp33_ASAP7_75t_L g8159 ( 
.A(n_7188),
.B(n_4675),
.Y(n_8159)
);

INVx2_ASAP7_75t_L g8160 ( 
.A(n_7240),
.Y(n_8160)
);

INVx2_ASAP7_75t_L g8161 ( 
.A(n_7256),
.Y(n_8161)
);

NAND3xp33_ASAP7_75t_L g8162 ( 
.A(n_7621),
.B(n_4677),
.C(n_4676),
.Y(n_8162)
);

INVx1_ASAP7_75t_L g8163 ( 
.A(n_7610),
.Y(n_8163)
);

INVx1_ASAP7_75t_L g8164 ( 
.A(n_7256),
.Y(n_8164)
);

NAND2xp5_ASAP7_75t_SL g8165 ( 
.A(n_7151),
.B(n_4678),
.Y(n_8165)
);

INVx2_ASAP7_75t_L g8166 ( 
.A(n_7288),
.Y(n_8166)
);

BUFx6f_ASAP7_75t_L g8167 ( 
.A(n_7288),
.Y(n_8167)
);

INVx2_ASAP7_75t_L g8168 ( 
.A(n_7155),
.Y(n_8168)
);

INVx3_ASAP7_75t_L g8169 ( 
.A(n_7227),
.Y(n_8169)
);

NAND2xp5_ASAP7_75t_L g8170 ( 
.A(n_7315),
.B(n_5105),
.Y(n_8170)
);

INVx1_ASAP7_75t_L g8171 ( 
.A(n_7400),
.Y(n_8171)
);

NOR2xp33_ASAP7_75t_L g8172 ( 
.A(n_7550),
.B(n_4680),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7423),
.Y(n_8173)
);

INVx1_ASAP7_75t_L g8174 ( 
.A(n_7433),
.Y(n_8174)
);

NOR2xp33_ASAP7_75t_L g8175 ( 
.A(n_7568),
.B(n_7511),
.Y(n_8175)
);

INVx1_ASAP7_75t_L g8176 ( 
.A(n_7163),
.Y(n_8176)
);

INVx4_ASAP7_75t_L g8177 ( 
.A(n_7489),
.Y(n_8177)
);

INVx2_ASAP7_75t_L g8178 ( 
.A(n_7625),
.Y(n_8178)
);

INVx2_ASAP7_75t_L g8179 ( 
.A(n_7598),
.Y(n_8179)
);

INVx2_ASAP7_75t_L g8180 ( 
.A(n_7222),
.Y(n_8180)
);

INVx2_ASAP7_75t_L g8181 ( 
.A(n_7342),
.Y(n_8181)
);

NAND2xp5_ASAP7_75t_SL g8182 ( 
.A(n_7241),
.B(n_4682),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_7425),
.Y(n_8183)
);

NAND2xp5_ASAP7_75t_SL g8184 ( 
.A(n_7603),
.B(n_4683),
.Y(n_8184)
);

INVx1_ASAP7_75t_L g8185 ( 
.A(n_7436),
.Y(n_8185)
);

INVx2_ASAP7_75t_L g8186 ( 
.A(n_7634),
.Y(n_8186)
);

INVx3_ASAP7_75t_L g8187 ( 
.A(n_7359),
.Y(n_8187)
);

BUFx3_ASAP7_75t_L g8188 ( 
.A(n_7177),
.Y(n_8188)
);

CKINVDCx11_ASAP7_75t_R g8189 ( 
.A(n_7184),
.Y(n_8189)
);

NAND2xp5_ASAP7_75t_L g8190 ( 
.A(n_7465),
.B(n_5106),
.Y(n_8190)
);

INVx1_ASAP7_75t_L g8191 ( 
.A(n_7469),
.Y(n_8191)
);

INVx1_ASAP7_75t_L g8192 ( 
.A(n_7142),
.Y(n_8192)
);

BUFx2_ASAP7_75t_L g8193 ( 
.A(n_7386),
.Y(n_8193)
);

NAND2xp33_ASAP7_75t_L g8194 ( 
.A(n_7427),
.B(n_4684),
.Y(n_8194)
);

NAND2xp5_ASAP7_75t_SL g8195 ( 
.A(n_7143),
.B(n_4685),
.Y(n_8195)
);

INVx2_ASAP7_75t_L g8196 ( 
.A(n_7578),
.Y(n_8196)
);

INVx1_ASAP7_75t_L g8197 ( 
.A(n_7566),
.Y(n_8197)
);

AND3x1_ASAP7_75t_L g8198 ( 
.A(n_7641),
.B(n_5124),
.C(n_5121),
.Y(n_8198)
);

BUFx2_ASAP7_75t_L g8199 ( 
.A(n_7183),
.Y(n_8199)
);

INVx1_ASAP7_75t_L g8200 ( 
.A(n_7569),
.Y(n_8200)
);

INVx2_ASAP7_75t_L g8201 ( 
.A(n_7620),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_7570),
.Y(n_8202)
);

INVx2_ASAP7_75t_L g8203 ( 
.A(n_7437),
.Y(n_8203)
);

NAND2xp5_ASAP7_75t_SL g8204 ( 
.A(n_7440),
.B(n_4686),
.Y(n_8204)
);

INVx2_ASAP7_75t_SL g8205 ( 
.A(n_7203),
.Y(n_8205)
);

INVx3_ASAP7_75t_L g8206 ( 
.A(n_7503),
.Y(n_8206)
);

INVx2_ASAP7_75t_L g8207 ( 
.A(n_7189),
.Y(n_8207)
);

INVx2_ASAP7_75t_SL g8208 ( 
.A(n_7874),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_7658),
.Y(n_8209)
);

AND2x2_ASAP7_75t_SL g8210 ( 
.A(n_7663),
.B(n_7734),
.Y(n_8210)
);

INVx1_ASAP7_75t_L g8211 ( 
.A(n_7660),
.Y(n_8211)
);

INVxp67_ASAP7_75t_L g8212 ( 
.A(n_7790),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_SL g8213 ( 
.A(n_7904),
.B(n_7176),
.Y(n_8213)
);

BUFx6f_ASAP7_75t_SL g8214 ( 
.A(n_7733),
.Y(n_8214)
);

NAND2xp5_ASAP7_75t_SL g8215 ( 
.A(n_7904),
.B(n_7505),
.Y(n_8215)
);

OR2x2_ASAP7_75t_L g8216 ( 
.A(n_7983),
.B(n_8007),
.Y(n_8216)
);

BUFx6f_ASAP7_75t_L g8217 ( 
.A(n_7657),
.Y(n_8217)
);

INVx2_ASAP7_75t_L g8218 ( 
.A(n_7946),
.Y(n_8218)
);

INVx1_ASAP7_75t_L g8219 ( 
.A(n_7662),
.Y(n_8219)
);

NAND2xp33_ASAP7_75t_L g8220 ( 
.A(n_7928),
.B(n_7192),
.Y(n_8220)
);

AND2x6_ASAP7_75t_L g8221 ( 
.A(n_7774),
.B(n_7243),
.Y(n_8221)
);

INVx1_ASAP7_75t_L g8222 ( 
.A(n_7665),
.Y(n_8222)
);

NOR2xp33_ASAP7_75t_L g8223 ( 
.A(n_7674),
.B(n_7275),
.Y(n_8223)
);

INVx1_ASAP7_75t_L g8224 ( 
.A(n_7670),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_7673),
.Y(n_8225)
);

AND2x2_ASAP7_75t_SL g8226 ( 
.A(n_7684),
.B(n_7462),
.Y(n_8226)
);

XNOR2x2_ASAP7_75t_L g8227 ( 
.A(n_8104),
.B(n_7438),
.Y(n_8227)
);

INVx1_ASAP7_75t_L g8228 ( 
.A(n_7679),
.Y(n_8228)
);

CKINVDCx20_ASAP7_75t_R g8229 ( 
.A(n_8189),
.Y(n_8229)
);

BUFx6f_ASAP7_75t_L g8230 ( 
.A(n_7657),
.Y(n_8230)
);

INVx2_ASAP7_75t_L g8231 ( 
.A(n_7837),
.Y(n_8231)
);

AOI22xp5_ASAP7_75t_L g8232 ( 
.A1(n_7659),
.A2(n_7482),
.B1(n_7426),
.B2(n_7524),
.Y(n_8232)
);

INVx1_ASAP7_75t_L g8233 ( 
.A(n_7680),
.Y(n_8233)
);

INVx3_ASAP7_75t_L g8234 ( 
.A(n_7874),
.Y(n_8234)
);

INVx2_ASAP7_75t_SL g8235 ( 
.A(n_7887),
.Y(n_8235)
);

AND2x2_ASAP7_75t_SL g8236 ( 
.A(n_8097),
.B(n_7460),
.Y(n_8236)
);

INVx1_ASAP7_75t_SL g8237 ( 
.A(n_8065),
.Y(n_8237)
);

INVx4_ASAP7_75t_L g8238 ( 
.A(n_7887),
.Y(n_8238)
);

NOR2xp33_ASAP7_75t_SL g8239 ( 
.A(n_7876),
.B(n_7471),
.Y(n_8239)
);

BUFx10_ASAP7_75t_L g8240 ( 
.A(n_7695),
.Y(n_8240)
);

NOR2xp33_ASAP7_75t_L g8241 ( 
.A(n_7783),
.B(n_7478),
.Y(n_8241)
);

NOR2xp33_ASAP7_75t_L g8242 ( 
.A(n_7771),
.B(n_7470),
.Y(n_8242)
);

NOR2xp33_ASAP7_75t_L g8243 ( 
.A(n_7681),
.B(n_4687),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_7683),
.Y(n_8244)
);

NAND2xp5_ASAP7_75t_L g8245 ( 
.A(n_7730),
.B(n_4689),
.Y(n_8245)
);

HB1xp67_ASAP7_75t_L g8246 ( 
.A(n_8064),
.Y(n_8246)
);

NAND2xp5_ASAP7_75t_SL g8247 ( 
.A(n_8036),
.B(n_4690),
.Y(n_8247)
);

AND2x4_ASAP7_75t_L g8248 ( 
.A(n_7927),
.B(n_7528),
.Y(n_8248)
);

INVx2_ASAP7_75t_L g8249 ( 
.A(n_7838),
.Y(n_8249)
);

NAND2xp5_ASAP7_75t_L g8250 ( 
.A(n_8012),
.B(n_4691),
.Y(n_8250)
);

CKINVDCx5p33_ASAP7_75t_R g8251 ( 
.A(n_7977),
.Y(n_8251)
);

BUFx2_ASAP7_75t_L g8252 ( 
.A(n_7959),
.Y(n_8252)
);

BUFx6f_ASAP7_75t_L g8253 ( 
.A(n_7716),
.Y(n_8253)
);

INVx2_ASAP7_75t_L g8254 ( 
.A(n_7846),
.Y(n_8254)
);

AOI22xp5_ASAP7_75t_L g8255 ( 
.A1(n_8085),
.A2(n_4700),
.B1(n_4701),
.B2(n_4695),
.Y(n_8255)
);

INVx1_ASAP7_75t_L g8256 ( 
.A(n_7693),
.Y(n_8256)
);

BUFx6f_ASAP7_75t_L g8257 ( 
.A(n_7716),
.Y(n_8257)
);

AND2x2_ASAP7_75t_SL g8258 ( 
.A(n_8199),
.B(n_4841),
.Y(n_8258)
);

CKINVDCx6p67_ASAP7_75t_R g8259 ( 
.A(n_7927),
.Y(n_8259)
);

BUFx4f_ASAP7_75t_L g8260 ( 
.A(n_7656),
.Y(n_8260)
);

INVx2_ASAP7_75t_L g8261 ( 
.A(n_7849),
.Y(n_8261)
);

NAND2xp5_ASAP7_75t_SL g8262 ( 
.A(n_8036),
.B(n_4706),
.Y(n_8262)
);

INVx4_ASAP7_75t_L g8263 ( 
.A(n_7692),
.Y(n_8263)
);

NAND2xp5_ASAP7_75t_SL g8264 ( 
.A(n_8119),
.B(n_4707),
.Y(n_8264)
);

AND2x6_ASAP7_75t_L g8265 ( 
.A(n_7781),
.B(n_5127),
.Y(n_8265)
);

NAND2xp5_ASAP7_75t_L g8266 ( 
.A(n_7918),
.B(n_4709),
.Y(n_8266)
);

INVx4_ASAP7_75t_L g8267 ( 
.A(n_7692),
.Y(n_8267)
);

NAND2xp5_ASAP7_75t_L g8268 ( 
.A(n_7918),
.B(n_4711),
.Y(n_8268)
);

INVx1_ASAP7_75t_L g8269 ( 
.A(n_7697),
.Y(n_8269)
);

INVx4_ASAP7_75t_L g8270 ( 
.A(n_7745),
.Y(n_8270)
);

NOR2xp33_ASAP7_75t_L g8271 ( 
.A(n_7845),
.B(n_4714),
.Y(n_8271)
);

BUFx6f_ASAP7_75t_L g8272 ( 
.A(n_8119),
.Y(n_8272)
);

INVxp67_ASAP7_75t_L g8273 ( 
.A(n_8193),
.Y(n_8273)
);

INVx2_ASAP7_75t_L g8274 ( 
.A(n_7852),
.Y(n_8274)
);

AND2x4_ASAP7_75t_SL g8275 ( 
.A(n_7763),
.B(n_5313),
.Y(n_8275)
);

AND2x2_ASAP7_75t_L g8276 ( 
.A(n_8154),
.B(n_5313),
.Y(n_8276)
);

INVx2_ASAP7_75t_L g8277 ( 
.A(n_7855),
.Y(n_8277)
);

INVx1_ASAP7_75t_L g8278 ( 
.A(n_7699),
.Y(n_8278)
);

INVx2_ASAP7_75t_L g8279 ( 
.A(n_7856),
.Y(n_8279)
);

NAND2xp5_ASAP7_75t_L g8280 ( 
.A(n_7918),
.B(n_4715),
.Y(n_8280)
);

AND2x6_ASAP7_75t_L g8281 ( 
.A(n_7786),
.B(n_5128),
.Y(n_8281)
);

BUFx6f_ASAP7_75t_L g8282 ( 
.A(n_7810),
.Y(n_8282)
);

INVx1_ASAP7_75t_L g8283 ( 
.A(n_7708),
.Y(n_8283)
);

INVx2_ASAP7_75t_L g8284 ( 
.A(n_7857),
.Y(n_8284)
);

INVx2_ASAP7_75t_SL g8285 ( 
.A(n_7745),
.Y(n_8285)
);

CKINVDCx5p33_ASAP7_75t_R g8286 ( 
.A(n_7999),
.Y(n_8286)
);

INVx1_ASAP7_75t_L g8287 ( 
.A(n_7709),
.Y(n_8287)
);

BUFx2_ASAP7_75t_L g8288 ( 
.A(n_7994),
.Y(n_8288)
);

AND2x2_ASAP7_75t_L g8289 ( 
.A(n_8172),
.B(n_5333),
.Y(n_8289)
);

INVx4_ASAP7_75t_SL g8290 ( 
.A(n_7733),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_7710),
.Y(n_8291)
);

INVx2_ASAP7_75t_L g8292 ( 
.A(n_7863),
.Y(n_8292)
);

INVx2_ASAP7_75t_L g8293 ( 
.A(n_7864),
.Y(n_8293)
);

AOI22xp33_ASAP7_75t_L g8294 ( 
.A1(n_7859),
.A2(n_7512),
.B1(n_7507),
.B2(n_5383),
.Y(n_8294)
);

INVx1_ASAP7_75t_L g8295 ( 
.A(n_7711),
.Y(n_8295)
);

BUFx6f_ASAP7_75t_L g8296 ( 
.A(n_7810),
.Y(n_8296)
);

INVx2_ASAP7_75t_L g8297 ( 
.A(n_7867),
.Y(n_8297)
);

INVx1_ASAP7_75t_L g8298 ( 
.A(n_7726),
.Y(n_8298)
);

INVx2_ASAP7_75t_L g8299 ( 
.A(n_7881),
.Y(n_8299)
);

NAND2xp5_ASAP7_75t_L g8300 ( 
.A(n_8019),
.B(n_7717),
.Y(n_8300)
);

INVx4_ASAP7_75t_L g8301 ( 
.A(n_7832),
.Y(n_8301)
);

INVx1_ASAP7_75t_L g8302 ( 
.A(n_7738),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7742),
.Y(n_8303)
);

INVx1_ASAP7_75t_L g8304 ( 
.A(n_7743),
.Y(n_8304)
);

AND2x6_ASAP7_75t_L g8305 ( 
.A(n_7823),
.B(n_5136),
.Y(n_8305)
);

INVx4_ASAP7_75t_L g8306 ( 
.A(n_7832),
.Y(n_8306)
);

INVx2_ASAP7_75t_L g8307 ( 
.A(n_7882),
.Y(n_8307)
);

AND2x6_ASAP7_75t_L g8308 ( 
.A(n_7850),
.B(n_5144),
.Y(n_8308)
);

INVx5_ASAP7_75t_L g8309 ( 
.A(n_7873),
.Y(n_8309)
);

BUFx8_ASAP7_75t_SL g8310 ( 
.A(n_8066),
.Y(n_8310)
);

NAND2xp5_ASAP7_75t_L g8311 ( 
.A(n_8019),
.B(n_4717),
.Y(n_8311)
);

BUFx2_ASAP7_75t_L g8312 ( 
.A(n_8147),
.Y(n_8312)
);

BUFx3_ASAP7_75t_L g8313 ( 
.A(n_7873),
.Y(n_8313)
);

BUFx3_ASAP7_75t_L g8314 ( 
.A(n_7729),
.Y(n_8314)
);

AND2x2_ASAP7_75t_L g8315 ( 
.A(n_7912),
.B(n_5333),
.Y(n_8315)
);

AND2x4_ASAP7_75t_L g8316 ( 
.A(n_7753),
.B(n_5157),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_7744),
.Y(n_8317)
);

INVx2_ASAP7_75t_L g8318 ( 
.A(n_7886),
.Y(n_8318)
);

NAND2xp5_ASAP7_75t_L g8319 ( 
.A(n_8019),
.B(n_4718),
.Y(n_8319)
);

BUFx6f_ASAP7_75t_L g8320 ( 
.A(n_7814),
.Y(n_8320)
);

NOR2xp33_ASAP7_75t_L g8321 ( 
.A(n_7740),
.B(n_4722),
.Y(n_8321)
);

INVx1_ASAP7_75t_L g8322 ( 
.A(n_7752),
.Y(n_8322)
);

INVx1_ASAP7_75t_L g8323 ( 
.A(n_7754),
.Y(n_8323)
);

NOR2xp33_ASAP7_75t_L g8324 ( 
.A(n_7917),
.B(n_4724),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_7768),
.Y(n_8325)
);

INVx3_ASAP7_75t_L g8326 ( 
.A(n_7848),
.Y(n_8326)
);

NAND2xp5_ASAP7_75t_L g8327 ( 
.A(n_7819),
.B(n_4725),
.Y(n_8327)
);

BUFx6f_ASAP7_75t_L g8328 ( 
.A(n_7814),
.Y(n_8328)
);

AND2x2_ASAP7_75t_L g8329 ( 
.A(n_7869),
.B(n_5383),
.Y(n_8329)
);

AND2x4_ASAP7_75t_L g8330 ( 
.A(n_7798),
.B(n_5177),
.Y(n_8330)
);

INVx2_ASAP7_75t_L g8331 ( 
.A(n_7888),
.Y(n_8331)
);

BUFx3_ASAP7_75t_L g8332 ( 
.A(n_7818),
.Y(n_8332)
);

NAND2xp5_ASAP7_75t_SL g8333 ( 
.A(n_7858),
.B(n_4726),
.Y(n_8333)
);

AND2x2_ASAP7_75t_L g8334 ( 
.A(n_7776),
.B(n_5468),
.Y(n_8334)
);

INVx2_ASAP7_75t_L g8335 ( 
.A(n_7890),
.Y(n_8335)
);

NOR2xp33_ASAP7_75t_L g8336 ( 
.A(n_7707),
.B(n_4728),
.Y(n_8336)
);

NAND2xp5_ASAP7_75t_SL g8337 ( 
.A(n_7858),
.B(n_4729),
.Y(n_8337)
);

BUFx6f_ASAP7_75t_L g8338 ( 
.A(n_7909),
.Y(n_8338)
);

INVx1_ASAP7_75t_SL g8339 ( 
.A(n_8127),
.Y(n_8339)
);

BUFx6f_ASAP7_75t_L g8340 ( 
.A(n_7909),
.Y(n_8340)
);

NAND2xp5_ASAP7_75t_SL g8341 ( 
.A(n_7958),
.B(n_4730),
.Y(n_8341)
);

CKINVDCx5p33_ASAP7_75t_R g8342 ( 
.A(n_7741),
.Y(n_8342)
);

NAND2xp5_ASAP7_75t_L g8343 ( 
.A(n_7820),
.B(n_4732),
.Y(n_8343)
);

AND2x2_ASAP7_75t_SL g8344 ( 
.A(n_8198),
.B(n_4866),
.Y(n_8344)
);

AND2x4_ASAP7_75t_L g8345 ( 
.A(n_7828),
.B(n_5182),
.Y(n_8345)
);

INVx2_ASAP7_75t_L g8346 ( 
.A(n_7897),
.Y(n_8346)
);

INVx2_ASAP7_75t_L g8347 ( 
.A(n_7899),
.Y(n_8347)
);

BUFx6f_ASAP7_75t_L g8348 ( 
.A(n_7958),
.Y(n_8348)
);

INVx3_ASAP7_75t_L g8349 ( 
.A(n_7868),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_7772),
.Y(n_8350)
);

INVx1_ASAP7_75t_L g8351 ( 
.A(n_7784),
.Y(n_8351)
);

INVx4_ASAP7_75t_SL g8352 ( 
.A(n_7712),
.Y(n_8352)
);

CKINVDCx5p33_ASAP7_75t_R g8353 ( 
.A(n_7809),
.Y(n_8353)
);

INVx2_ASAP7_75t_L g8354 ( 
.A(n_7900),
.Y(n_8354)
);

BUFx3_ASAP7_75t_L g8355 ( 
.A(n_7677),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_7788),
.Y(n_8356)
);

AO22x2_ASAP7_75t_L g8357 ( 
.A1(n_7794),
.A2(n_5196),
.B1(n_5197),
.B2(n_5194),
.Y(n_8357)
);

INVx1_ASAP7_75t_L g8358 ( 
.A(n_7795),
.Y(n_8358)
);

BUFx6f_ASAP7_75t_L g8359 ( 
.A(n_7978),
.Y(n_8359)
);

BUFx6f_ASAP7_75t_L g8360 ( 
.A(n_7978),
.Y(n_8360)
);

INVx2_ASAP7_75t_L g8361 ( 
.A(n_7913),
.Y(n_8361)
);

AND2x4_ASAP7_75t_L g8362 ( 
.A(n_7755),
.B(n_5207),
.Y(n_8362)
);

INVx2_ASAP7_75t_L g8363 ( 
.A(n_7914),
.Y(n_8363)
);

AND2x2_ASAP7_75t_L g8364 ( 
.A(n_7762),
.B(n_8095),
.Y(n_8364)
);

INVx1_ASAP7_75t_L g8365 ( 
.A(n_7800),
.Y(n_8365)
);

AND2x4_ASAP7_75t_L g8366 ( 
.A(n_8116),
.B(n_5209),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_7804),
.Y(n_8367)
);

INVx2_ASAP7_75t_L g8368 ( 
.A(n_7921),
.Y(n_8368)
);

INVx1_ASAP7_75t_SL g8369 ( 
.A(n_7911),
.Y(n_8369)
);

AOI22xp5_ASAP7_75t_L g8370 ( 
.A1(n_7835),
.A2(n_4737),
.B1(n_4738),
.B2(n_4733),
.Y(n_8370)
);

BUFx2_ASAP7_75t_L g8371 ( 
.A(n_8151),
.Y(n_8371)
);

INVx1_ASAP7_75t_L g8372 ( 
.A(n_7806),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7811),
.Y(n_8373)
);

INVx1_ASAP7_75t_L g8374 ( 
.A(n_7825),
.Y(n_8374)
);

NAND2xp5_ASAP7_75t_L g8375 ( 
.A(n_7854),
.B(n_4739),
.Y(n_8375)
);

AND2x2_ASAP7_75t_L g8376 ( 
.A(n_8175),
.B(n_5468),
.Y(n_8376)
);

INVx1_ASAP7_75t_L g8377 ( 
.A(n_7827),
.Y(n_8377)
);

BUFx6f_ASAP7_75t_L g8378 ( 
.A(n_7985),
.Y(n_8378)
);

INVx3_ASAP7_75t_L g8379 ( 
.A(n_7948),
.Y(n_8379)
);

OAI22xp5_ASAP7_75t_L g8380 ( 
.A1(n_7949),
.A2(n_4745),
.B1(n_4751),
.B2(n_4744),
.Y(n_8380)
);

BUFx3_ASAP7_75t_L g8381 ( 
.A(n_7878),
.Y(n_8381)
);

INVx3_ASAP7_75t_L g8382 ( 
.A(n_7671),
.Y(n_8382)
);

AND2x6_ASAP7_75t_L g8383 ( 
.A(n_7920),
.B(n_7936),
.Y(n_8383)
);

INVx1_ASAP7_75t_L g8384 ( 
.A(n_7830),
.Y(n_8384)
);

NOR2xp33_ASAP7_75t_SL g8385 ( 
.A(n_8177),
.B(n_5472),
.Y(n_8385)
);

NAND2xp5_ASAP7_75t_SL g8386 ( 
.A(n_7985),
.B(n_4754),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_7833),
.Y(n_8387)
);

BUFx6f_ASAP7_75t_L g8388 ( 
.A(n_8082),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_7834),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_7839),
.Y(n_8390)
);

INVx2_ASAP7_75t_L g8391 ( 
.A(n_7925),
.Y(n_8391)
);

INVx2_ASAP7_75t_SL g8392 ( 
.A(n_7961),
.Y(n_8392)
);

INVx2_ASAP7_75t_L g8393 ( 
.A(n_7930),
.Y(n_8393)
);

BUFx2_ASAP7_75t_L g8394 ( 
.A(n_7727),
.Y(n_8394)
);

CKINVDCx5p33_ASAP7_75t_R g8395 ( 
.A(n_7844),
.Y(n_8395)
);

INVx1_ASAP7_75t_L g8396 ( 
.A(n_7840),
.Y(n_8396)
);

AND2x4_ASAP7_75t_L g8397 ( 
.A(n_8037),
.B(n_5213),
.Y(n_8397)
);

NOR2xp33_ASAP7_75t_L g8398 ( 
.A(n_7866),
.B(n_4758),
.Y(n_8398)
);

INVx3_ASAP7_75t_L g8399 ( 
.A(n_7655),
.Y(n_8399)
);

INVx1_ASAP7_75t_L g8400 ( 
.A(n_7841),
.Y(n_8400)
);

INVx1_ASAP7_75t_L g8401 ( 
.A(n_7842),
.Y(n_8401)
);

INVx2_ASAP7_75t_L g8402 ( 
.A(n_7931),
.Y(n_8402)
);

AND2x2_ASAP7_75t_L g8403 ( 
.A(n_8072),
.B(n_5472),
.Y(n_8403)
);

BUFx3_ASAP7_75t_L g8404 ( 
.A(n_7721),
.Y(n_8404)
);

INVx2_ASAP7_75t_L g8405 ( 
.A(n_7932),
.Y(n_8405)
);

BUFx2_ASAP7_75t_L g8406 ( 
.A(n_7787),
.Y(n_8406)
);

INVx4_ASAP7_75t_L g8407 ( 
.A(n_8082),
.Y(n_8407)
);

AND2x4_ASAP7_75t_L g8408 ( 
.A(n_7997),
.B(n_5214),
.Y(n_8408)
);

AND2x6_ASAP7_75t_L g8409 ( 
.A(n_7736),
.B(n_5220),
.Y(n_8409)
);

INVx4_ASAP7_75t_L g8410 ( 
.A(n_8096),
.Y(n_8410)
);

INVx1_ASAP7_75t_L g8411 ( 
.A(n_7847),
.Y(n_8411)
);

INVx5_ASAP7_75t_L g8412 ( 
.A(n_8187),
.Y(n_8412)
);

NAND2xp5_ASAP7_75t_SL g8413 ( 
.A(n_8096),
.B(n_4759),
.Y(n_8413)
);

NAND2xp5_ASAP7_75t_L g8414 ( 
.A(n_8020),
.B(n_8034),
.Y(n_8414)
);

CKINVDCx16_ASAP7_75t_R g8415 ( 
.A(n_7988),
.Y(n_8415)
);

INVx3_ASAP7_75t_L g8416 ( 
.A(n_8108),
.Y(n_8416)
);

AND2x2_ASAP7_75t_L g8417 ( 
.A(n_7891),
.B(n_4762),
.Y(n_8417)
);

NOR2xp33_ASAP7_75t_L g8418 ( 
.A(n_8084),
.B(n_4763),
.Y(n_8418)
);

INVx6_ASAP7_75t_L g8419 ( 
.A(n_7905),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_7851),
.Y(n_8420)
);

NOR2xp33_ASAP7_75t_L g8421 ( 
.A(n_7902),
.B(n_4764),
.Y(n_8421)
);

AND2x4_ASAP7_75t_L g8422 ( 
.A(n_8158),
.B(n_7865),
.Y(n_8422)
);

OR2x2_ASAP7_75t_L g8423 ( 
.A(n_8196),
.B(n_4766),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_7853),
.Y(n_8424)
);

INVx1_ASAP7_75t_L g8425 ( 
.A(n_7861),
.Y(n_8425)
);

INVx5_ASAP7_75t_L g8426 ( 
.A(n_7935),
.Y(n_8426)
);

CKINVDCx5p33_ASAP7_75t_R g8427 ( 
.A(n_8188),
.Y(n_8427)
);

INVx2_ASAP7_75t_L g8428 ( 
.A(n_7938),
.Y(n_8428)
);

INVx2_ASAP7_75t_L g8429 ( 
.A(n_7942),
.Y(n_8429)
);

NOR2xp33_ASAP7_75t_L g8430 ( 
.A(n_8083),
.B(n_4767),
.Y(n_8430)
);

INVxp67_ASAP7_75t_SL g8431 ( 
.A(n_7843),
.Y(n_8431)
);

INVx4_ASAP7_75t_L g8432 ( 
.A(n_8108),
.Y(n_8432)
);

OR2x6_ASAP7_75t_L g8433 ( 
.A(n_8205),
.B(n_4883),
.Y(n_8433)
);

NAND2xp5_ASAP7_75t_L g8434 ( 
.A(n_8042),
.B(n_4769),
.Y(n_8434)
);

INVx3_ASAP7_75t_L g8435 ( 
.A(n_8131),
.Y(n_8435)
);

NOR2xp33_ASAP7_75t_L g8436 ( 
.A(n_8057),
.B(n_8078),
.Y(n_8436)
);

NOR2xp33_ASAP7_75t_L g8437 ( 
.A(n_8081),
.B(n_4771),
.Y(n_8437)
);

AND2x4_ASAP7_75t_L g8438 ( 
.A(n_7785),
.B(n_5230),
.Y(n_8438)
);

BUFx6f_ASAP7_75t_SL g8439 ( 
.A(n_8093),
.Y(n_8439)
);

NAND2xp5_ASAP7_75t_L g8440 ( 
.A(n_8044),
.B(n_4775),
.Y(n_8440)
);

NAND3xp33_ASAP7_75t_L g8441 ( 
.A(n_8023),
.B(n_4777),
.C(n_4776),
.Y(n_8441)
);

AND2x4_ASAP7_75t_L g8442 ( 
.A(n_8040),
.B(n_5236),
.Y(n_8442)
);

BUFx6f_ASAP7_75t_L g8443 ( 
.A(n_8131),
.Y(n_8443)
);

INVx1_ASAP7_75t_L g8444 ( 
.A(n_7862),
.Y(n_8444)
);

INVx5_ASAP7_75t_L g8445 ( 
.A(n_8167),
.Y(n_8445)
);

BUFx10_ASAP7_75t_L g8446 ( 
.A(n_8002),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_7871),
.Y(n_8447)
);

CKINVDCx20_ASAP7_75t_R g8448 ( 
.A(n_8022),
.Y(n_8448)
);

NAND2xp5_ASAP7_75t_SL g8449 ( 
.A(n_8167),
.B(n_8179),
.Y(n_8449)
);

NAND2x1p5_ASAP7_75t_L g8450 ( 
.A(n_8038),
.B(n_5238),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_7872),
.Y(n_8451)
);

INVx1_ASAP7_75t_L g8452 ( 
.A(n_7875),
.Y(n_8452)
);

INVx2_ASAP7_75t_L g8453 ( 
.A(n_7945),
.Y(n_8453)
);

INVx3_ASAP7_75t_L g8454 ( 
.A(n_8122),
.Y(n_8454)
);

INVx2_ASAP7_75t_L g8455 ( 
.A(n_7826),
.Y(n_8455)
);

BUFx2_ASAP7_75t_L g8456 ( 
.A(n_7969),
.Y(n_8456)
);

NAND2xp33_ASAP7_75t_SL g8457 ( 
.A(n_8180),
.B(n_4778),
.Y(n_8457)
);

INVx3_ASAP7_75t_L g8458 ( 
.A(n_8129),
.Y(n_8458)
);

HB1xp67_ASAP7_75t_L g8459 ( 
.A(n_8156),
.Y(n_8459)
);

NAND2xp5_ASAP7_75t_SL g8460 ( 
.A(n_8178),
.B(n_4782),
.Y(n_8460)
);

OR2x2_ASAP7_75t_L g8461 ( 
.A(n_8190),
.B(n_4783),
.Y(n_8461)
);

INVxp67_ASAP7_75t_SL g8462 ( 
.A(n_8142),
.Y(n_8462)
);

BUFx3_ASAP7_75t_L g8463 ( 
.A(n_7672),
.Y(n_8463)
);

INVxp67_ASAP7_75t_L g8464 ( 
.A(n_8163),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_7879),
.Y(n_8465)
);

INVx1_ASAP7_75t_L g8466 ( 
.A(n_7901),
.Y(n_8466)
);

INVx2_ASAP7_75t_L g8467 ( 
.A(n_7836),
.Y(n_8467)
);

INVx3_ASAP7_75t_L g8468 ( 
.A(n_7687),
.Y(n_8468)
);

AND2x6_ASAP7_75t_L g8469 ( 
.A(n_8206),
.B(n_5240),
.Y(n_8469)
);

NAND2xp5_ASAP7_75t_L g8470 ( 
.A(n_8048),
.B(n_4784),
.Y(n_8470)
);

AND2x4_ASAP7_75t_L g8471 ( 
.A(n_8144),
.B(n_7722),
.Y(n_8471)
);

INVx1_ASAP7_75t_L g8472 ( 
.A(n_7903),
.Y(n_8472)
);

INVx1_ASAP7_75t_L g8473 ( 
.A(n_7922),
.Y(n_8473)
);

INVx1_ASAP7_75t_L g8474 ( 
.A(n_7926),
.Y(n_8474)
);

AND2x4_ASAP7_75t_L g8475 ( 
.A(n_7777),
.B(n_5245),
.Y(n_8475)
);

INVx8_ASAP7_75t_L g8476 ( 
.A(n_7813),
.Y(n_8476)
);

NAND2xp5_ASAP7_75t_L g8477 ( 
.A(n_8053),
.B(n_4786),
.Y(n_8477)
);

INVx5_ASAP7_75t_L g8478 ( 
.A(n_7803),
.Y(n_8478)
);

AND2x4_ASAP7_75t_L g8479 ( 
.A(n_7870),
.B(n_5252),
.Y(n_8479)
);

AND2x4_ASAP7_75t_L g8480 ( 
.A(n_7950),
.B(n_5254),
.Y(n_8480)
);

OAI22xp5_ASAP7_75t_L g8481 ( 
.A1(n_8087),
.A2(n_4789),
.B1(n_4791),
.B2(n_4787),
.Y(n_8481)
);

INVx1_ASAP7_75t_L g8482 ( 
.A(n_7934),
.Y(n_8482)
);

NOR2xp33_ASAP7_75t_L g8483 ( 
.A(n_8099),
.B(n_4798),
.Y(n_8483)
);

INVx4_ASAP7_75t_L g8484 ( 
.A(n_7691),
.Y(n_8484)
);

INVx3_ASAP7_75t_L g8485 ( 
.A(n_7703),
.Y(n_8485)
);

NAND2xp5_ASAP7_75t_SL g8486 ( 
.A(n_8051),
.B(n_4801),
.Y(n_8486)
);

INVx1_ASAP7_75t_L g8487 ( 
.A(n_7939),
.Y(n_8487)
);

OR2x2_ASAP7_75t_L g8488 ( 
.A(n_8058),
.B(n_4802),
.Y(n_8488)
);

NAND2xp5_ASAP7_75t_L g8489 ( 
.A(n_8054),
.B(n_4805),
.Y(n_8489)
);

NAND2xp5_ASAP7_75t_SL g8490 ( 
.A(n_7906),
.B(n_4806),
.Y(n_8490)
);

BUFx3_ASAP7_75t_L g8491 ( 
.A(n_8133),
.Y(n_8491)
);

BUFx2_ASAP7_75t_L g8492 ( 
.A(n_7969),
.Y(n_8492)
);

INVx1_ASAP7_75t_L g8493 ( 
.A(n_7940),
.Y(n_8493)
);

INVx1_ASAP7_75t_L g8494 ( 
.A(n_7952),
.Y(n_8494)
);

INVx1_ASAP7_75t_L g8495 ( 
.A(n_7956),
.Y(n_8495)
);

BUFx6f_ASAP7_75t_L g8496 ( 
.A(n_8169),
.Y(n_8496)
);

NOR2xp33_ASAP7_75t_L g8497 ( 
.A(n_8110),
.B(n_4807),
.Y(n_8497)
);

INVx1_ASAP7_75t_SL g8498 ( 
.A(n_8001),
.Y(n_8498)
);

INVx2_ASAP7_75t_L g8499 ( 
.A(n_7676),
.Y(n_8499)
);

NAND3xp33_ASAP7_75t_L g8500 ( 
.A(n_7748),
.B(n_4817),
.C(n_4809),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_7963),
.Y(n_8501)
);

INVx2_ASAP7_75t_L g8502 ( 
.A(n_7678),
.Y(n_8502)
);

HB1xp67_ASAP7_75t_L g8503 ( 
.A(n_8145),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_8030),
.Y(n_8504)
);

NAND2xp5_ASAP7_75t_SL g8505 ( 
.A(n_7765),
.B(n_4818),
.Y(n_8505)
);

INVx2_ASAP7_75t_SL g8506 ( 
.A(n_8135),
.Y(n_8506)
);

INVx1_ASAP7_75t_L g8507 ( 
.A(n_8031),
.Y(n_8507)
);

INVx2_ASAP7_75t_L g8508 ( 
.A(n_7682),
.Y(n_8508)
);

BUFx10_ASAP7_75t_L g8509 ( 
.A(n_8027),
.Y(n_8509)
);

OR2x2_ASAP7_75t_L g8510 ( 
.A(n_8191),
.B(n_4820),
.Y(n_8510)
);

OR2x2_ASAP7_75t_L g8511 ( 
.A(n_8170),
.B(n_4821),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_8033),
.Y(n_8512)
);

NAND2xp5_ASAP7_75t_SL g8513 ( 
.A(n_7971),
.B(n_4827),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_8039),
.Y(n_8514)
);

INVx1_ASAP7_75t_L g8515 ( 
.A(n_8041),
.Y(n_8515)
);

NAND3xp33_ASAP7_75t_L g8516 ( 
.A(n_7769),
.B(n_4833),
.C(n_4829),
.Y(n_8516)
);

INVx2_ASAP7_75t_L g8517 ( 
.A(n_7685),
.Y(n_8517)
);

AND2x6_ASAP7_75t_L g8518 ( 
.A(n_8203),
.B(n_5259),
.Y(n_8518)
);

BUFx6f_ASAP7_75t_L g8519 ( 
.A(n_8138),
.Y(n_8519)
);

BUFx3_ASAP7_75t_L g8520 ( 
.A(n_8141),
.Y(n_8520)
);

INVx1_ASAP7_75t_SL g8521 ( 
.A(n_8094),
.Y(n_8521)
);

NAND2xp5_ASAP7_75t_SL g8522 ( 
.A(n_7892),
.B(n_4835),
.Y(n_8522)
);

INVx2_ASAP7_75t_L g8523 ( 
.A(n_7688),
.Y(n_8523)
);

BUFx2_ASAP7_75t_L g8524 ( 
.A(n_8094),
.Y(n_8524)
);

INVx2_ASAP7_75t_L g8525 ( 
.A(n_7689),
.Y(n_8525)
);

INVx5_ASAP7_75t_L g8526 ( 
.A(n_7803),
.Y(n_8526)
);

INVx5_ASAP7_75t_L g8527 ( 
.A(n_7805),
.Y(n_8527)
);

INVx2_ASAP7_75t_L g8528 ( 
.A(n_7690),
.Y(n_8528)
);

INVx1_ASAP7_75t_SL g8529 ( 
.A(n_7779),
.Y(n_8529)
);

INVx2_ASAP7_75t_L g8530 ( 
.A(n_7694),
.Y(n_8530)
);

AOI22xp5_ASAP7_75t_L g8531 ( 
.A1(n_7816),
.A2(n_4840),
.B1(n_4842),
.B2(n_4839),
.Y(n_8531)
);

BUFx10_ASAP7_75t_L g8532 ( 
.A(n_7910),
.Y(n_8532)
);

INVx2_ASAP7_75t_L g8533 ( 
.A(n_7698),
.Y(n_8533)
);

NAND2xp5_ASAP7_75t_SL g8534 ( 
.A(n_7669),
.B(n_7668),
.Y(n_8534)
);

INVx1_ASAP7_75t_L g8535 ( 
.A(n_8046),
.Y(n_8535)
);

INVx1_ASAP7_75t_L g8536 ( 
.A(n_8047),
.Y(n_8536)
);

INVx1_ASAP7_75t_L g8537 ( 
.A(n_7724),
.Y(n_8537)
);

INVx1_ASAP7_75t_L g8538 ( 
.A(n_7700),
.Y(n_8538)
);

INVx4_ASAP7_75t_L g8539 ( 
.A(n_7751),
.Y(n_8539)
);

INVx3_ASAP7_75t_L g8540 ( 
.A(n_8146),
.Y(n_8540)
);

INVx1_ASAP7_75t_L g8541 ( 
.A(n_7702),
.Y(n_8541)
);

NAND2xp5_ASAP7_75t_SL g8542 ( 
.A(n_7780),
.B(n_4844),
.Y(n_8542)
);

NOR2xp33_ASAP7_75t_L g8543 ( 
.A(n_8120),
.B(n_4846),
.Y(n_8543)
);

BUFx3_ASAP7_75t_L g8544 ( 
.A(n_8150),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_7704),
.Y(n_8545)
);

NOR2xp33_ASAP7_75t_L g8546 ( 
.A(n_8123),
.B(n_4850),
.Y(n_8546)
);

INVx2_ASAP7_75t_L g8547 ( 
.A(n_7705),
.Y(n_8547)
);

INVx4_ASAP7_75t_L g8548 ( 
.A(n_7751),
.Y(n_8548)
);

NOR2xp33_ASAP7_75t_L g8549 ( 
.A(n_7908),
.B(n_4854),
.Y(n_8549)
);

INVx1_ASAP7_75t_L g8550 ( 
.A(n_7706),
.Y(n_8550)
);

NAND2xp33_ASAP7_75t_L g8551 ( 
.A(n_8140),
.B(n_4855),
.Y(n_8551)
);

INVx2_ASAP7_75t_L g8552 ( 
.A(n_7713),
.Y(n_8552)
);

NAND2xp5_ASAP7_75t_SL g8553 ( 
.A(n_8010),
.B(n_4859),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_7714),
.Y(n_8554)
);

INVx1_ASAP7_75t_L g8555 ( 
.A(n_7719),
.Y(n_8555)
);

INVx2_ASAP7_75t_L g8556 ( 
.A(n_7723),
.Y(n_8556)
);

INVxp33_ASAP7_75t_L g8557 ( 
.A(n_8013),
.Y(n_8557)
);

AND2x2_ASAP7_75t_L g8558 ( 
.A(n_7919),
.B(n_7796),
.Y(n_8558)
);

INVx1_ASAP7_75t_L g8559 ( 
.A(n_7728),
.Y(n_8559)
);

INVx1_ASAP7_75t_L g8560 ( 
.A(n_7731),
.Y(n_8560)
);

INVx1_ASAP7_75t_L g8561 ( 
.A(n_7735),
.Y(n_8561)
);

INVx1_ASAP7_75t_L g8562 ( 
.A(n_7739),
.Y(n_8562)
);

OAI21xp33_ASAP7_75t_L g8563 ( 
.A1(n_7767),
.A2(n_4861),
.B(n_4860),
.Y(n_8563)
);

INVx1_ASAP7_75t_L g8564 ( 
.A(n_7746),
.Y(n_8564)
);

BUFx6f_ASAP7_75t_L g8565 ( 
.A(n_8152),
.Y(n_8565)
);

INVx2_ASAP7_75t_SL g8566 ( 
.A(n_8153),
.Y(n_8566)
);

AOI22xp5_ASAP7_75t_L g8567 ( 
.A1(n_7880),
.A2(n_4863),
.B1(n_4867),
.B2(n_4862),
.Y(n_8567)
);

NAND2xp5_ASAP7_75t_L g8568 ( 
.A(n_7766),
.B(n_4868),
.Y(n_8568)
);

NOR2xp33_ASAP7_75t_L g8569 ( 
.A(n_7929),
.B(n_4871),
.Y(n_8569)
);

INVx5_ASAP7_75t_L g8570 ( 
.A(n_7805),
.Y(n_8570)
);

INVx3_ASAP7_75t_L g8571 ( 
.A(n_8160),
.Y(n_8571)
);

NAND2x1p5_ASAP7_75t_L g8572 ( 
.A(n_8137),
.B(n_5261),
.Y(n_8572)
);

OAI22xp5_ASAP7_75t_L g8573 ( 
.A1(n_7992),
.A2(n_4878),
.B1(n_4879),
.B2(n_4874),
.Y(n_8573)
);

INVx2_ASAP7_75t_SL g8574 ( 
.A(n_8161),
.Y(n_8574)
);

INVx3_ASAP7_75t_L g8575 ( 
.A(n_8166),
.Y(n_8575)
);

INVx4_ASAP7_75t_L g8576 ( 
.A(n_8207),
.Y(n_8576)
);

INVx4_ASAP7_75t_L g8577 ( 
.A(n_8098),
.Y(n_8577)
);

BUFx10_ASAP7_75t_L g8578 ( 
.A(n_7664),
.Y(n_8578)
);

INVx1_ASAP7_75t_L g8579 ( 
.A(n_7747),
.Y(n_8579)
);

INVx2_ASAP7_75t_L g8580 ( 
.A(n_7749),
.Y(n_8580)
);

INVx1_ASAP7_75t_L g8581 ( 
.A(n_7750),
.Y(n_8581)
);

INVx2_ASAP7_75t_L g8582 ( 
.A(n_7760),
.Y(n_8582)
);

AND2x2_ASAP7_75t_L g8583 ( 
.A(n_8130),
.B(n_4880),
.Y(n_8583)
);

NOR2xp33_ASAP7_75t_L g8584 ( 
.A(n_8005),
.B(n_4882),
.Y(n_8584)
);

NAND2xp5_ASAP7_75t_L g8585 ( 
.A(n_7974),
.B(n_4888),
.Y(n_8585)
);

AND2x4_ASAP7_75t_L g8586 ( 
.A(n_7955),
.B(n_5262),
.Y(n_8586)
);

INVx4_ASAP7_75t_L g8587 ( 
.A(n_8100),
.Y(n_8587)
);

INVx4_ASAP7_75t_L g8588 ( 
.A(n_8103),
.Y(n_8588)
);

AND2x4_ASAP7_75t_L g8589 ( 
.A(n_8176),
.B(n_5271),
.Y(n_8589)
);

NOR2xp33_ASAP7_75t_L g8590 ( 
.A(n_8192),
.B(n_4895),
.Y(n_8590)
);

BUFx10_ASAP7_75t_L g8591 ( 
.A(n_7701),
.Y(n_8591)
);

INVx2_ASAP7_75t_L g8592 ( 
.A(n_7761),
.Y(n_8592)
);

AND2x2_ASAP7_75t_L g8593 ( 
.A(n_7831),
.B(n_4896),
.Y(n_8593)
);

NAND2xp5_ASAP7_75t_SL g8594 ( 
.A(n_7817),
.B(n_4903),
.Y(n_8594)
);

INVx2_ASAP7_75t_L g8595 ( 
.A(n_7764),
.Y(n_8595)
);

BUFx6f_ASAP7_75t_L g8596 ( 
.A(n_8106),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_7773),
.Y(n_8597)
);

NAND2xp5_ASAP7_75t_L g8598 ( 
.A(n_7975),
.B(n_4908),
.Y(n_8598)
);

BUFx6f_ASAP7_75t_L g8599 ( 
.A(n_8056),
.Y(n_8599)
);

INVx2_ASAP7_75t_L g8600 ( 
.A(n_7778),
.Y(n_8600)
);

INVx1_ASAP7_75t_SL g8601 ( 
.A(n_7789),
.Y(n_8601)
);

INVx1_ASAP7_75t_L g8602 ( 
.A(n_7782),
.Y(n_8602)
);

AOI22xp33_ASAP7_75t_L g8603 ( 
.A1(n_8201),
.A2(n_4910),
.B1(n_4912),
.B2(n_4909),
.Y(n_8603)
);

HB1xp67_ASAP7_75t_L g8604 ( 
.A(n_8149),
.Y(n_8604)
);

BUFx6f_ASAP7_75t_L g8605 ( 
.A(n_8059),
.Y(n_8605)
);

INVx2_ASAP7_75t_L g8606 ( 
.A(n_7793),
.Y(n_8606)
);

NOR2xp33_ASAP7_75t_L g8607 ( 
.A(n_7953),
.B(n_4913),
.Y(n_8607)
);

NAND2x1p5_ASAP7_75t_L g8608 ( 
.A(n_7986),
.B(n_8164),
.Y(n_8608)
);

NAND2xp5_ASAP7_75t_L g8609 ( 
.A(n_7775),
.B(n_4914),
.Y(n_8609)
);

BUFx6f_ASAP7_75t_L g8610 ( 
.A(n_8060),
.Y(n_8610)
);

AOI22xp33_ASAP7_75t_L g8611 ( 
.A1(n_7797),
.A2(n_7802),
.B1(n_8143),
.B2(n_7661),
.Y(n_8611)
);

INVx2_ASAP7_75t_L g8612 ( 
.A(n_7667),
.Y(n_8612)
);

NOR2xp33_ASAP7_75t_L g8613 ( 
.A(n_7970),
.B(n_4916),
.Y(n_8613)
);

INVx2_ASAP7_75t_L g8614 ( 
.A(n_7821),
.Y(n_8614)
);

BUFx6f_ASAP7_75t_L g8615 ( 
.A(n_8061),
.Y(n_8615)
);

INVx3_ASAP7_75t_L g8616 ( 
.A(n_8067),
.Y(n_8616)
);

INVx1_ASAP7_75t_L g8617 ( 
.A(n_7822),
.Y(n_8617)
);

CKINVDCx5p33_ASAP7_75t_R g8618 ( 
.A(n_8197),
.Y(n_8618)
);

BUFx3_ASAP7_75t_L g8619 ( 
.A(n_8068),
.Y(n_8619)
);

INVx5_ASAP7_75t_L g8620 ( 
.A(n_8069),
.Y(n_8620)
);

INVx2_ASAP7_75t_L g8621 ( 
.A(n_7807),
.Y(n_8621)
);

NAND2xp33_ASAP7_75t_L g8622 ( 
.A(n_8181),
.B(n_4928),
.Y(n_8622)
);

INVx2_ASAP7_75t_L g8623 ( 
.A(n_8006),
.Y(n_8623)
);

INVx2_ASAP7_75t_L g8624 ( 
.A(n_8008),
.Y(n_8624)
);

NAND2xp5_ASAP7_75t_L g8625 ( 
.A(n_7758),
.B(n_4930),
.Y(n_8625)
);

NAND2xp5_ASAP7_75t_L g8626 ( 
.A(n_7715),
.B(n_4932),
.Y(n_8626)
);

AND2x2_ASAP7_75t_SL g8627 ( 
.A(n_8194),
.B(n_4886),
.Y(n_8627)
);

AND2x4_ASAP7_75t_L g8628 ( 
.A(n_8171),
.B(n_5273),
.Y(n_8628)
);

INVxp33_ASAP7_75t_L g8629 ( 
.A(n_8195),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_7799),
.Y(n_8630)
);

AND2x2_ASAP7_75t_L g8631 ( 
.A(n_7792),
.B(n_4934),
.Y(n_8631)
);

NAND2xp33_ASAP7_75t_L g8632 ( 
.A(n_8032),
.B(n_7943),
.Y(n_8632)
);

INVx1_ASAP7_75t_L g8633 ( 
.A(n_7965),
.Y(n_8633)
);

HB1xp67_ASAP7_75t_L g8634 ( 
.A(n_8173),
.Y(n_8634)
);

AND2x2_ASAP7_75t_L g8635 ( 
.A(n_8174),
.B(n_4935),
.Y(n_8635)
);

BUFx6f_ASAP7_75t_L g8636 ( 
.A(n_8071),
.Y(n_8636)
);

BUFx3_ASAP7_75t_L g8637 ( 
.A(n_8074),
.Y(n_8637)
);

AND2x2_ASAP7_75t_L g8638 ( 
.A(n_7686),
.B(n_4938),
.Y(n_8638)
);

INVx1_ASAP7_75t_L g8639 ( 
.A(n_7972),
.Y(n_8639)
);

INVx4_ASAP7_75t_L g8640 ( 
.A(n_8075),
.Y(n_8640)
);

BUFx6f_ASAP7_75t_L g8641 ( 
.A(n_8076),
.Y(n_8641)
);

BUFx10_ASAP7_75t_L g8642 ( 
.A(n_8139),
.Y(n_8642)
);

INVx2_ASAP7_75t_L g8643 ( 
.A(n_7951),
.Y(n_8643)
);

INVx1_ASAP7_75t_L g8644 ( 
.A(n_8009),
.Y(n_8644)
);

NAND2xp5_ASAP7_75t_L g8645 ( 
.A(n_8045),
.B(n_4942),
.Y(n_8645)
);

INVx1_ASAP7_75t_L g8646 ( 
.A(n_7996),
.Y(n_8646)
);

INVx1_ASAP7_75t_L g8647 ( 
.A(n_8003),
.Y(n_8647)
);

NAND2xp5_ASAP7_75t_SL g8648 ( 
.A(n_7725),
.B(n_4943),
.Y(n_8648)
);

BUFx6f_ASAP7_75t_L g8649 ( 
.A(n_8079),
.Y(n_8649)
);

AND2x2_ASAP7_75t_SL g8650 ( 
.A(n_7737),
.B(n_4900),
.Y(n_8650)
);

INVx3_ASAP7_75t_L g8651 ( 
.A(n_8088),
.Y(n_8651)
);

AND2x4_ASAP7_75t_L g8652 ( 
.A(n_8089),
.B(n_5276),
.Y(n_8652)
);

INVx1_ASAP7_75t_L g8653 ( 
.A(n_7801),
.Y(n_8653)
);

AND2x4_ASAP7_75t_L g8654 ( 
.A(n_8090),
.B(n_8092),
.Y(n_8654)
);

AND2x2_ASAP7_75t_L g8655 ( 
.A(n_8128),
.B(n_4949),
.Y(n_8655)
);

AOI22xp5_ASAP7_75t_L g8656 ( 
.A1(n_7894),
.A2(n_4957),
.B1(n_4958),
.B2(n_4952),
.Y(n_8656)
);

NAND2xp5_ASAP7_75t_SL g8657 ( 
.A(n_7732),
.B(n_4959),
.Y(n_8657)
);

BUFx10_ASAP7_75t_L g8658 ( 
.A(n_8200),
.Y(n_8658)
);

INVx1_ASAP7_75t_L g8659 ( 
.A(n_7812),
.Y(n_8659)
);

AND2x4_ASAP7_75t_L g8660 ( 
.A(n_8126),
.B(n_5278),
.Y(n_8660)
);

NAND3xp33_ASAP7_75t_L g8661 ( 
.A(n_8035),
.B(n_4962),
.C(n_4960),
.Y(n_8661)
);

INVx2_ASAP7_75t_L g8662 ( 
.A(n_7957),
.Y(n_8662)
);

INVxp67_ASAP7_75t_L g8663 ( 
.A(n_8052),
.Y(n_8663)
);

CKINVDCx5p33_ASAP7_75t_R g8664 ( 
.A(n_8202),
.Y(n_8664)
);

AND2x2_ASAP7_75t_SL g8665 ( 
.A(n_8080),
.B(n_4901),
.Y(n_8665)
);

INVx5_ASAP7_75t_L g8666 ( 
.A(n_8168),
.Y(n_8666)
);

INVx1_ASAP7_75t_L g8667 ( 
.A(n_7960),
.Y(n_8667)
);

INVx1_ASAP7_75t_L g8668 ( 
.A(n_7962),
.Y(n_8668)
);

INVx2_ASAP7_75t_L g8669 ( 
.A(n_7967),
.Y(n_8669)
);

CKINVDCx14_ASAP7_75t_R g8670 ( 
.A(n_7933),
.Y(n_8670)
);

HB1xp67_ASAP7_75t_L g8671 ( 
.A(n_8109),
.Y(n_8671)
);

NOR2xp33_ASAP7_75t_L g8672 ( 
.A(n_7980),
.B(n_4963),
.Y(n_8672)
);

INVx2_ASAP7_75t_L g8673 ( 
.A(n_7968),
.Y(n_8673)
);

NAND2xp5_ASAP7_75t_SL g8674 ( 
.A(n_8136),
.B(n_4965),
.Y(n_8674)
);

INVx4_ASAP7_75t_L g8675 ( 
.A(n_8112),
.Y(n_8675)
);

BUFx6f_ASAP7_75t_L g8676 ( 
.A(n_8113),
.Y(n_8676)
);

INVx2_ASAP7_75t_L g8677 ( 
.A(n_7973),
.Y(n_8677)
);

NAND2xp33_ASAP7_75t_R g8678 ( 
.A(n_8183),
.B(n_8185),
.Y(n_8678)
);

INVx1_ASAP7_75t_L g8679 ( 
.A(n_7979),
.Y(n_8679)
);

INVx1_ASAP7_75t_SL g8680 ( 
.A(n_8117),
.Y(n_8680)
);

BUFx3_ASAP7_75t_L g8681 ( 
.A(n_8118),
.Y(n_8681)
);

AND2x4_ASAP7_75t_L g8682 ( 
.A(n_8124),
.B(n_5280),
.Y(n_8682)
);

NAND2xp5_ASAP7_75t_L g8683 ( 
.A(n_7815),
.B(n_4967),
.Y(n_8683)
);

INVx1_ASAP7_75t_L g8684 ( 
.A(n_7998),
.Y(n_8684)
);

NAND2xp5_ASAP7_75t_SL g8685 ( 
.A(n_7756),
.B(n_4970),
.Y(n_8685)
);

INVx1_ASAP7_75t_L g8686 ( 
.A(n_7824),
.Y(n_8686)
);

INVx1_ASAP7_75t_L g8687 ( 
.A(n_7829),
.Y(n_8687)
);

OR2x2_ASAP7_75t_L g8688 ( 
.A(n_8050),
.B(n_4972),
.Y(n_8688)
);

NAND2xp5_ASAP7_75t_L g8689 ( 
.A(n_7984),
.B(n_4974),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_7860),
.Y(n_8690)
);

NAND2xp5_ASAP7_75t_SL g8691 ( 
.A(n_8186),
.B(n_4975),
.Y(n_8691)
);

INVx2_ASAP7_75t_L g8692 ( 
.A(n_7993),
.Y(n_8692)
);

INVx2_ASAP7_75t_L g8693 ( 
.A(n_7995),
.Y(n_8693)
);

AOI22xp5_ASAP7_75t_L g8694 ( 
.A1(n_8043),
.A2(n_4980),
.B1(n_4984),
.B2(n_4978),
.Y(n_8694)
);

INVx3_ASAP7_75t_L g8695 ( 
.A(n_8016),
.Y(n_8695)
);

INVx5_ASAP7_75t_L g8696 ( 
.A(n_8004),
.Y(n_8696)
);

NAND2xp5_ASAP7_75t_SL g8697 ( 
.A(n_8162),
.B(n_4987),
.Y(n_8697)
);

INVx3_ASAP7_75t_L g8698 ( 
.A(n_8063),
.Y(n_8698)
);

INVx4_ASAP7_75t_L g8699 ( 
.A(n_8015),
.Y(n_8699)
);

INVx2_ASAP7_75t_L g8700 ( 
.A(n_7982),
.Y(n_8700)
);

NAND2xp5_ASAP7_75t_SL g8701 ( 
.A(n_7654),
.B(n_4988),
.Y(n_8701)
);

BUFx6f_ASAP7_75t_L g8702 ( 
.A(n_7720),
.Y(n_8702)
);

AND2x4_ASAP7_75t_L g8703 ( 
.A(n_8132),
.B(n_5285),
.Y(n_8703)
);

INVx1_ASAP7_75t_L g8704 ( 
.A(n_7877),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_7987),
.Y(n_8705)
);

NAND2xp5_ASAP7_75t_SL g8706 ( 
.A(n_7976),
.B(n_7885),
.Y(n_8706)
);

INVx1_ASAP7_75t_L g8707 ( 
.A(n_7883),
.Y(n_8707)
);

NOR2xp33_ASAP7_75t_L g8708 ( 
.A(n_7893),
.B(n_4992),
.Y(n_8708)
);

BUFx3_ASAP7_75t_L g8709 ( 
.A(n_7941),
.Y(n_8709)
);

INVx2_ASAP7_75t_L g8710 ( 
.A(n_7989),
.Y(n_8710)
);

AND2x2_ASAP7_75t_L g8711 ( 
.A(n_7954),
.B(n_4998),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_7898),
.Y(n_8712)
);

INVx1_ASAP7_75t_L g8713 ( 
.A(n_7915),
.Y(n_8713)
);

INVx2_ASAP7_75t_L g8714 ( 
.A(n_7990),
.Y(n_8714)
);

BUFx3_ASAP7_75t_L g8715 ( 
.A(n_7944),
.Y(n_8715)
);

INVx2_ASAP7_75t_L g8716 ( 
.A(n_7666),
.Y(n_8716)
);

HB1xp67_ASAP7_75t_L g8717 ( 
.A(n_7770),
.Y(n_8717)
);

AOI22xp33_ASAP7_75t_L g8718 ( 
.A1(n_8155),
.A2(n_8017),
.B1(n_8025),
.B2(n_8000),
.Y(n_8718)
);

AOI21xp5_ASAP7_75t_L g8719 ( 
.A1(n_8551),
.A2(n_8632),
.B(n_8414),
.Y(n_8719)
);

BUFx3_ASAP7_75t_L g8720 ( 
.A(n_8253),
.Y(n_8720)
);

INVx2_ASAP7_75t_SL g8721 ( 
.A(n_8476),
.Y(n_8721)
);

NAND2xp5_ASAP7_75t_SL g8722 ( 
.A(n_8210),
.B(n_7675),
.Y(n_8722)
);

INVx2_ASAP7_75t_L g8723 ( 
.A(n_8231),
.Y(n_8723)
);

OAI22xp5_ASAP7_75t_L g8724 ( 
.A1(n_8558),
.A2(n_8024),
.B1(n_8107),
.B2(n_8091),
.Y(n_8724)
);

AOI21xp5_ASAP7_75t_L g8725 ( 
.A1(n_8486),
.A2(n_8029),
.B(n_8026),
.Y(n_8725)
);

OAI22x1_ASAP7_75t_SL g8726 ( 
.A1(n_8229),
.A2(n_5001),
.B1(n_5002),
.B2(n_5000),
.Y(n_8726)
);

NOR2xp33_ASAP7_75t_L g8727 ( 
.A(n_8430),
.B(n_7895),
.Y(n_8727)
);

OAI221xp5_ASAP7_75t_L g8728 ( 
.A1(n_8324),
.A2(n_7937),
.B1(n_8134),
.B2(n_8111),
.C(n_8121),
.Y(n_8728)
);

NAND2xp5_ASAP7_75t_L g8729 ( 
.A(n_8436),
.B(n_7947),
.Y(n_8729)
);

INVx8_ASAP7_75t_L g8730 ( 
.A(n_8214),
.Y(n_8730)
);

NAND2xp5_ASAP7_75t_L g8731 ( 
.A(n_8686),
.B(n_8070),
.Y(n_8731)
);

AND2x2_ASAP7_75t_L g8732 ( 
.A(n_8364),
.B(n_7966),
.Y(n_8732)
);

NAND2xp5_ASAP7_75t_L g8733 ( 
.A(n_8687),
.B(n_7896),
.Y(n_8733)
);

INVx1_ASAP7_75t_L g8734 ( 
.A(n_8209),
.Y(n_8734)
);

INVx2_ASAP7_75t_L g8735 ( 
.A(n_8249),
.Y(n_8735)
);

INVx2_ASAP7_75t_L g8736 ( 
.A(n_8254),
.Y(n_8736)
);

NAND2xp5_ASAP7_75t_SL g8737 ( 
.A(n_8627),
.B(n_8073),
.Y(n_8737)
);

NOR2xp33_ASAP7_75t_L g8738 ( 
.A(n_8336),
.B(n_7907),
.Y(n_8738)
);

NAND2xp5_ASAP7_75t_SL g8739 ( 
.A(n_8650),
.B(n_7718),
.Y(n_8739)
);

NAND3xp33_ASAP7_75t_L g8740 ( 
.A(n_8271),
.B(n_8159),
.C(n_8102),
.Y(n_8740)
);

OAI221xp5_ASAP7_75t_L g8741 ( 
.A1(n_8321),
.A2(n_8018),
.B1(n_8184),
.B2(n_7916),
.C(n_7924),
.Y(n_8741)
);

INVx1_ASAP7_75t_L g8742 ( 
.A(n_8211),
.Y(n_8742)
);

OAI22xp33_ASAP7_75t_L g8743 ( 
.A1(n_8415),
.A2(n_8148),
.B1(n_7923),
.B2(n_7808),
.Y(n_8743)
);

NAND2xp5_ASAP7_75t_L g8744 ( 
.A(n_8690),
.B(n_7791),
.Y(n_8744)
);

AOI22xp33_ASAP7_75t_L g8745 ( 
.A1(n_8223),
.A2(n_7964),
.B1(n_8028),
.B2(n_8182),
.Y(n_8745)
);

INVxp67_ASAP7_75t_L g8746 ( 
.A(n_8246),
.Y(n_8746)
);

NAND2xp5_ASAP7_75t_L g8747 ( 
.A(n_8704),
.B(n_7759),
.Y(n_8747)
);

INVxp67_ASAP7_75t_SL g8748 ( 
.A(n_8715),
.Y(n_8748)
);

NAND2xp5_ASAP7_75t_L g8749 ( 
.A(n_8707),
.B(n_7757),
.Y(n_8749)
);

NAND2xp5_ASAP7_75t_L g8750 ( 
.A(n_8712),
.B(n_8204),
.Y(n_8750)
);

NAND2xp5_ASAP7_75t_SL g8751 ( 
.A(n_8529),
.B(n_8114),
.Y(n_8751)
);

INVx1_ASAP7_75t_L g8752 ( 
.A(n_8219),
.Y(n_8752)
);

NOR2xp33_ASAP7_75t_L g8753 ( 
.A(n_8237),
.B(n_7884),
.Y(n_8753)
);

INVx2_ASAP7_75t_SL g8754 ( 
.A(n_8445),
.Y(n_8754)
);

NAND2xp5_ASAP7_75t_SL g8755 ( 
.A(n_8601),
.B(n_7696),
.Y(n_8755)
);

INVx2_ASAP7_75t_L g8756 ( 
.A(n_8261),
.Y(n_8756)
);

INVx2_ASAP7_75t_L g8757 ( 
.A(n_8274),
.Y(n_8757)
);

BUFx5_ASAP7_75t_L g8758 ( 
.A(n_8644),
.Y(n_8758)
);

NAND2xp5_ASAP7_75t_SL g8759 ( 
.A(n_8300),
.B(n_7981),
.Y(n_8759)
);

NOR2xp33_ASAP7_75t_L g8760 ( 
.A(n_8339),
.B(n_7889),
.Y(n_8760)
);

INVx2_ASAP7_75t_L g8761 ( 
.A(n_8277),
.Y(n_8761)
);

NAND2xp5_ASAP7_75t_SL g8762 ( 
.A(n_8446),
.B(n_7991),
.Y(n_8762)
);

NOR2xp33_ASAP7_75t_L g8763 ( 
.A(n_8216),
.B(n_8557),
.Y(n_8763)
);

AOI22xp5_ASAP7_75t_L g8764 ( 
.A1(n_8241),
.A2(n_8165),
.B1(n_8125),
.B2(n_8115),
.Y(n_8764)
);

INVx1_ASAP7_75t_L g8765 ( 
.A(n_8222),
.Y(n_8765)
);

NAND2xp5_ASAP7_75t_L g8766 ( 
.A(n_8713),
.B(n_8049),
.Y(n_8766)
);

INVx1_ASAP7_75t_L g8767 ( 
.A(n_8224),
.Y(n_8767)
);

AOI22xp5_ASAP7_75t_L g8768 ( 
.A1(n_8584),
.A2(n_8062),
.B1(n_8086),
.B2(n_8077),
.Y(n_8768)
);

NAND2xp5_ASAP7_75t_L g8769 ( 
.A(n_8684),
.B(n_8653),
.Y(n_8769)
);

NAND2xp5_ASAP7_75t_SL g8770 ( 
.A(n_8509),
.B(n_8157),
.Y(n_8770)
);

INVx1_ASAP7_75t_L g8771 ( 
.A(n_8225),
.Y(n_8771)
);

INVx1_ASAP7_75t_L g8772 ( 
.A(n_8228),
.Y(n_8772)
);

NAND2xp5_ASAP7_75t_L g8773 ( 
.A(n_8659),
.B(n_8101),
.Y(n_8773)
);

NAND2xp5_ASAP7_75t_SL g8774 ( 
.A(n_8702),
.B(n_8105),
.Y(n_8774)
);

NAND2xp33_ASAP7_75t_L g8775 ( 
.A(n_8383),
.B(n_8251),
.Y(n_8775)
);

INVx2_ASAP7_75t_L g8776 ( 
.A(n_8279),
.Y(n_8776)
);

INVx1_ASAP7_75t_L g8777 ( 
.A(n_8233),
.Y(n_8777)
);

CKINVDCx5p33_ASAP7_75t_R g8778 ( 
.A(n_8310),
.Y(n_8778)
);

OAI22xp33_ASAP7_75t_L g8779 ( 
.A1(n_8385),
.A2(n_5005),
.B1(n_5009),
.B2(n_5004),
.Y(n_8779)
);

NAND2xp5_ASAP7_75t_L g8780 ( 
.A(n_8276),
.B(n_5011),
.Y(n_8780)
);

INVx2_ASAP7_75t_L g8781 ( 
.A(n_8284),
.Y(n_8781)
);

NAND2xp5_ASAP7_75t_L g8782 ( 
.A(n_8289),
.B(n_5012),
.Y(n_8782)
);

NAND2xp5_ASAP7_75t_L g8783 ( 
.A(n_8630),
.B(n_5013),
.Y(n_8783)
);

AOI22xp33_ASAP7_75t_L g8784 ( 
.A1(n_8236),
.A2(n_8014),
.B1(n_8021),
.B2(n_8011),
.Y(n_8784)
);

NOR2xp33_ASAP7_75t_L g8785 ( 
.A(n_8273),
.B(n_5015),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_8244),
.Y(n_8786)
);

NOR2xp33_ASAP7_75t_L g8787 ( 
.A(n_8212),
.B(n_8252),
.Y(n_8787)
);

NAND2xp5_ASAP7_75t_SL g8788 ( 
.A(n_8702),
.B(n_8055),
.Y(n_8788)
);

NAND2xp5_ASAP7_75t_L g8789 ( 
.A(n_8537),
.B(n_5017),
.Y(n_8789)
);

NAND2xp5_ASAP7_75t_L g8790 ( 
.A(n_8315),
.B(n_5022),
.Y(n_8790)
);

INVx1_ASAP7_75t_L g8791 ( 
.A(n_8256),
.Y(n_8791)
);

NAND2xp5_ASAP7_75t_L g8792 ( 
.A(n_8376),
.B(n_5023),
.Y(n_8792)
);

NAND2xp5_ASAP7_75t_L g8793 ( 
.A(n_8403),
.B(n_5025),
.Y(n_8793)
);

NAND2xp5_ASAP7_75t_L g8794 ( 
.A(n_8329),
.B(n_5028),
.Y(n_8794)
);

INVx2_ASAP7_75t_L g8795 ( 
.A(n_8292),
.Y(n_8795)
);

NAND2xp5_ASAP7_75t_L g8796 ( 
.A(n_8655),
.B(n_5030),
.Y(n_8796)
);

AOI22xp5_ASAP7_75t_L g8797 ( 
.A1(n_8242),
.A2(n_5034),
.B1(n_5035),
.B2(n_5032),
.Y(n_8797)
);

NAND2xp5_ASAP7_75t_L g8798 ( 
.A(n_8462),
.B(n_5036),
.Y(n_8798)
);

NAND2xp5_ASAP7_75t_SL g8799 ( 
.A(n_8445),
.B(n_8478),
.Y(n_8799)
);

NAND2xp5_ASAP7_75t_SL g8800 ( 
.A(n_8478),
.B(n_5040),
.Y(n_8800)
);

NAND2xp5_ASAP7_75t_L g8801 ( 
.A(n_8334),
.B(n_5041),
.Y(n_8801)
);

INVx2_ASAP7_75t_SL g8802 ( 
.A(n_8253),
.Y(n_8802)
);

INVx2_ASAP7_75t_L g8803 ( 
.A(n_8293),
.Y(n_8803)
);

NAND2xp5_ASAP7_75t_SL g8804 ( 
.A(n_8526),
.B(n_5042),
.Y(n_8804)
);

INVx1_ASAP7_75t_L g8805 ( 
.A(n_8269),
.Y(n_8805)
);

AND2x6_ASAP7_75t_SL g8806 ( 
.A(n_8248),
.B(n_5291),
.Y(n_8806)
);

NAND2xp5_ASAP7_75t_L g8807 ( 
.A(n_8369),
.B(n_5048),
.Y(n_8807)
);

NAND3xp33_ASAP7_75t_L g8808 ( 
.A(n_8631),
.B(n_5050),
.C(n_5049),
.Y(n_8808)
);

OR2x2_ASAP7_75t_L g8809 ( 
.A(n_8498),
.B(n_5296),
.Y(n_8809)
);

INVx1_ASAP7_75t_L g8810 ( 
.A(n_8278),
.Y(n_8810)
);

NAND2xp5_ASAP7_75t_L g8811 ( 
.A(n_8663),
.B(n_5052),
.Y(n_8811)
);

BUFx3_ASAP7_75t_L g8812 ( 
.A(n_8257),
.Y(n_8812)
);

NAND2xp5_ASAP7_75t_L g8813 ( 
.A(n_8437),
.B(n_5055),
.Y(n_8813)
);

NAND2xp5_ASAP7_75t_SL g8814 ( 
.A(n_8526),
.B(n_5057),
.Y(n_8814)
);

NAND2xp5_ASAP7_75t_SL g8815 ( 
.A(n_8527),
.B(n_5061),
.Y(n_8815)
);

NOR2xp33_ASAP7_75t_L g8816 ( 
.A(n_8288),
.B(n_5063),
.Y(n_8816)
);

NAND2xp5_ASAP7_75t_SL g8817 ( 
.A(n_8527),
.B(n_5064),
.Y(n_8817)
);

NAND2xp5_ASAP7_75t_SL g8818 ( 
.A(n_8570),
.B(n_5065),
.Y(n_8818)
);

NAND2xp5_ASAP7_75t_L g8819 ( 
.A(n_8483),
.B(n_5066),
.Y(n_8819)
);

INVx8_ASAP7_75t_L g8820 ( 
.A(n_8383),
.Y(n_8820)
);

NAND2xp5_ASAP7_75t_SL g8821 ( 
.A(n_8570),
.B(n_5067),
.Y(n_8821)
);

NOR2xp67_ASAP7_75t_L g8822 ( 
.A(n_8309),
.B(n_3),
.Y(n_8822)
);

AND2x4_ASAP7_75t_L g8823 ( 
.A(n_8355),
.B(n_5297),
.Y(n_8823)
);

INVx1_ASAP7_75t_L g8824 ( 
.A(n_8283),
.Y(n_8824)
);

INVx2_ASAP7_75t_SL g8825 ( 
.A(n_8257),
.Y(n_8825)
);

INVxp67_ASAP7_75t_L g8826 ( 
.A(n_8503),
.Y(n_8826)
);

NOR2xp33_ASAP7_75t_L g8827 ( 
.A(n_8394),
.B(n_5069),
.Y(n_8827)
);

INVx2_ASAP7_75t_L g8828 ( 
.A(n_8297),
.Y(n_8828)
);

AOI22xp33_ASAP7_75t_L g8829 ( 
.A1(n_8227),
.A2(n_5074),
.B1(n_5077),
.B2(n_5070),
.Y(n_8829)
);

INVxp67_ASAP7_75t_SL g8830 ( 
.A(n_8604),
.Y(n_8830)
);

INVx2_ASAP7_75t_L g8831 ( 
.A(n_8299),
.Y(n_8831)
);

INVx2_ASAP7_75t_SL g8832 ( 
.A(n_8272),
.Y(n_8832)
);

INVx2_ASAP7_75t_SL g8833 ( 
.A(n_8272),
.Y(n_8833)
);

AND2x4_ASAP7_75t_SL g8834 ( 
.A(n_8240),
.B(n_5302),
.Y(n_8834)
);

INVx2_ASAP7_75t_L g8835 ( 
.A(n_8307),
.Y(n_8835)
);

CKINVDCx5p33_ASAP7_75t_R g8836 ( 
.A(n_8286),
.Y(n_8836)
);

INVx2_ASAP7_75t_SL g8837 ( 
.A(n_8260),
.Y(n_8837)
);

AOI22xp33_ASAP7_75t_SL g8838 ( 
.A1(n_8357),
.A2(n_5305),
.B1(n_5306),
.B2(n_5303),
.Y(n_8838)
);

NAND2xp5_ASAP7_75t_L g8839 ( 
.A(n_8497),
.B(n_5078),
.Y(n_8839)
);

NAND2xp5_ASAP7_75t_L g8840 ( 
.A(n_8543),
.B(n_5079),
.Y(n_8840)
);

O2A1O1Ixp33_ASAP7_75t_L g8841 ( 
.A1(n_8522),
.A2(n_5318),
.B(n_5320),
.C(n_5310),
.Y(n_8841)
);

INVx2_ASAP7_75t_L g8842 ( 
.A(n_8318),
.Y(n_8842)
);

NAND2xp5_ASAP7_75t_L g8843 ( 
.A(n_8546),
.B(n_5080),
.Y(n_8843)
);

INVx1_ASAP7_75t_L g8844 ( 
.A(n_8287),
.Y(n_8844)
);

INVx2_ASAP7_75t_L g8845 ( 
.A(n_8331),
.Y(n_8845)
);

INVx2_ASAP7_75t_SL g8846 ( 
.A(n_8217),
.Y(n_8846)
);

NAND2xp5_ASAP7_75t_L g8847 ( 
.A(n_8511),
.B(n_5083),
.Y(n_8847)
);

BUFx6f_ASAP7_75t_L g8848 ( 
.A(n_8217),
.Y(n_8848)
);

OAI22xp33_ASAP7_75t_L g8849 ( 
.A1(n_8255),
.A2(n_5087),
.B1(n_5090),
.B2(n_5085),
.Y(n_8849)
);

NOR2xp33_ASAP7_75t_L g8850 ( 
.A(n_8406),
.B(n_5091),
.Y(n_8850)
);

NAND2xp5_ASAP7_75t_L g8851 ( 
.A(n_8634),
.B(n_5092),
.Y(n_8851)
);

AND2x2_ASAP7_75t_L g8852 ( 
.A(n_8417),
.B(n_5094),
.Y(n_8852)
);

NAND2xp5_ASAP7_75t_SL g8853 ( 
.A(n_8258),
.B(n_5098),
.Y(n_8853)
);

NAND2xp5_ASAP7_75t_L g8854 ( 
.A(n_8665),
.B(n_5100),
.Y(n_8854)
);

INVx1_ASAP7_75t_L g8855 ( 
.A(n_8291),
.Y(n_8855)
);

CKINVDCx5p33_ASAP7_75t_R g8856 ( 
.A(n_8259),
.Y(n_8856)
);

OR2x2_ASAP7_75t_L g8857 ( 
.A(n_8488),
.B(n_5324),
.Y(n_8857)
);

INVx4_ASAP7_75t_L g8858 ( 
.A(n_8263),
.Y(n_8858)
);

NAND2xp5_ASAP7_75t_L g8859 ( 
.A(n_8431),
.B(n_5107),
.Y(n_8859)
);

INVx2_ASAP7_75t_SL g8860 ( 
.A(n_8230),
.Y(n_8860)
);

INVx2_ASAP7_75t_L g8861 ( 
.A(n_8335),
.Y(n_8861)
);

BUFx6f_ASAP7_75t_L g8862 ( 
.A(n_8230),
.Y(n_8862)
);

AOI22xp33_ASAP7_75t_L g8863 ( 
.A1(n_8593),
.A2(n_5112),
.B1(n_5113),
.B2(n_5110),
.Y(n_8863)
);

NAND2xp5_ASAP7_75t_L g8864 ( 
.A(n_8464),
.B(n_5114),
.Y(n_8864)
);

INVx2_ASAP7_75t_L g8865 ( 
.A(n_8346),
.Y(n_8865)
);

NAND2xp5_ASAP7_75t_SL g8866 ( 
.A(n_8309),
.B(n_5115),
.Y(n_8866)
);

CKINVDCx5p33_ASAP7_75t_R g8867 ( 
.A(n_8439),
.Y(n_8867)
);

AOI22xp5_ASAP7_75t_L g8868 ( 
.A1(n_8622),
.A2(n_8711),
.B1(n_8448),
.B2(n_8708),
.Y(n_8868)
);

NAND2xp5_ASAP7_75t_L g8869 ( 
.A(n_8459),
.B(n_5117),
.Y(n_8869)
);

INVx2_ASAP7_75t_L g8870 ( 
.A(n_8347),
.Y(n_8870)
);

INVx1_ASAP7_75t_L g8871 ( 
.A(n_8295),
.Y(n_8871)
);

NOR2xp33_ASAP7_75t_L g8872 ( 
.A(n_8312),
.B(n_5118),
.Y(n_8872)
);

NAND2xp5_ASAP7_75t_L g8873 ( 
.A(n_8461),
.B(n_8398),
.Y(n_8873)
);

INVx1_ASAP7_75t_L g8874 ( 
.A(n_8298),
.Y(n_8874)
);

INVx1_ASAP7_75t_L g8875 ( 
.A(n_8302),
.Y(n_8875)
);

NOR2xp33_ASAP7_75t_L g8876 ( 
.A(n_8371),
.B(n_5122),
.Y(n_8876)
);

NAND2xp5_ASAP7_75t_L g8877 ( 
.A(n_8418),
.B(n_5123),
.Y(n_8877)
);

AOI22xp33_ASAP7_75t_L g8878 ( 
.A1(n_8652),
.A2(n_5126),
.B1(n_5130),
.B2(n_5125),
.Y(n_8878)
);

NAND2x1p5_ASAP7_75t_L g8879 ( 
.A(n_8267),
.B(n_5326),
.Y(n_8879)
);

NAND2xp5_ASAP7_75t_SL g8880 ( 
.A(n_8718),
.B(n_5131),
.Y(n_8880)
);

INVx2_ASAP7_75t_L g8881 ( 
.A(n_8354),
.Y(n_8881)
);

OAI22xp5_ASAP7_75t_L g8882 ( 
.A1(n_8441),
.A2(n_5133),
.B1(n_5135),
.B2(n_5132),
.Y(n_8882)
);

INVx1_ASAP7_75t_L g8883 ( 
.A(n_8303),
.Y(n_8883)
);

AOI22xp5_ASAP7_75t_L g8884 ( 
.A1(n_8265),
.A2(n_5138),
.B1(n_5141),
.B2(n_5137),
.Y(n_8884)
);

NAND2xp5_ASAP7_75t_L g8885 ( 
.A(n_8232),
.B(n_8304),
.Y(n_8885)
);

NOR2xp33_ASAP7_75t_L g8886 ( 
.A(n_8629),
.B(n_5145),
.Y(n_8886)
);

NAND2xp5_ASAP7_75t_L g8887 ( 
.A(n_8317),
.B(n_5148),
.Y(n_8887)
);

OR2x2_ASAP7_75t_L g8888 ( 
.A(n_8521),
.B(n_5329),
.Y(n_8888)
);

NAND2xp5_ASAP7_75t_L g8889 ( 
.A(n_8322),
.B(n_8323),
.Y(n_8889)
);

HB1xp67_ASAP7_75t_L g8890 ( 
.A(n_8671),
.Y(n_8890)
);

INVx1_ASAP7_75t_L g8891 ( 
.A(n_8325),
.Y(n_8891)
);

OR2x2_ASAP7_75t_L g8892 ( 
.A(n_8456),
.B(n_5331),
.Y(n_8892)
);

NAND2xp5_ASAP7_75t_L g8893 ( 
.A(n_8350),
.B(n_5149),
.Y(n_8893)
);

NAND2xp5_ASAP7_75t_L g8894 ( 
.A(n_8351),
.B(n_8356),
.Y(n_8894)
);

INVx1_ASAP7_75t_L g8895 ( 
.A(n_8358),
.Y(n_8895)
);

INVx1_ASAP7_75t_L g8896 ( 
.A(n_8365),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_8367),
.Y(n_8897)
);

NAND2xp5_ASAP7_75t_L g8898 ( 
.A(n_8372),
.B(n_5151),
.Y(n_8898)
);

BUFx3_ASAP7_75t_L g8899 ( 
.A(n_8314),
.Y(n_8899)
);

AOI22xp5_ASAP7_75t_L g8900 ( 
.A1(n_8265),
.A2(n_5154),
.B1(n_5155),
.B2(n_5153),
.Y(n_8900)
);

NOR2xp33_ASAP7_75t_L g8901 ( 
.A(n_8576),
.B(n_5159),
.Y(n_8901)
);

INVx2_ASAP7_75t_L g8902 ( 
.A(n_8361),
.Y(n_8902)
);

NAND2xp5_ASAP7_75t_L g8903 ( 
.A(n_8373),
.B(n_5160),
.Y(n_8903)
);

OAI22xp5_ASAP7_75t_L g8904 ( 
.A1(n_8327),
.A2(n_5162),
.B1(n_5164),
.B2(n_5161),
.Y(n_8904)
);

NAND2xp5_ASAP7_75t_L g8905 ( 
.A(n_8374),
.B(n_5166),
.Y(n_8905)
);

NAND2xp5_ASAP7_75t_L g8906 ( 
.A(n_8377),
.B(n_5169),
.Y(n_8906)
);

NOR2xp33_ASAP7_75t_L g8907 ( 
.A(n_8332),
.B(n_5171),
.Y(n_8907)
);

AOI22xp33_ASAP7_75t_L g8908 ( 
.A1(n_8682),
.A2(n_5176),
.B1(n_5179),
.B2(n_5173),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_8384),
.Y(n_8909)
);

NAND2xp33_ASAP7_75t_L g8910 ( 
.A(n_8618),
.B(n_5180),
.Y(n_8910)
);

INVx1_ASAP7_75t_L g8911 ( 
.A(n_8387),
.Y(n_8911)
);

INVx1_ASAP7_75t_L g8912 ( 
.A(n_8389),
.Y(n_8912)
);

AOI22xp5_ASAP7_75t_L g8913 ( 
.A1(n_8281),
.A2(n_5183),
.B1(n_5185),
.B2(n_5181),
.Y(n_8913)
);

INVx4_ASAP7_75t_L g8914 ( 
.A(n_8238),
.Y(n_8914)
);

NAND2xp5_ASAP7_75t_SL g8915 ( 
.A(n_8539),
.B(n_5186),
.Y(n_8915)
);

OR2x2_ASAP7_75t_L g8916 ( 
.A(n_8492),
.B(n_5334),
.Y(n_8916)
);

NAND2xp5_ASAP7_75t_SL g8917 ( 
.A(n_8548),
.B(n_5187),
.Y(n_8917)
);

NAND2xp5_ASAP7_75t_SL g8918 ( 
.A(n_8664),
.B(n_5190),
.Y(n_8918)
);

NOR2xp33_ASAP7_75t_L g8919 ( 
.A(n_8709),
.B(n_5191),
.Y(n_8919)
);

INVx2_ASAP7_75t_L g8920 ( 
.A(n_8363),
.Y(n_8920)
);

NAND2xp5_ASAP7_75t_L g8921 ( 
.A(n_8390),
.B(n_5193),
.Y(n_8921)
);

INVx2_ASAP7_75t_L g8922 ( 
.A(n_8368),
.Y(n_8922)
);

INVx2_ASAP7_75t_SL g8923 ( 
.A(n_8419),
.Y(n_8923)
);

OAI22xp5_ASAP7_75t_L g8924 ( 
.A1(n_8343),
.A2(n_5200),
.B1(n_5201),
.B2(n_5195),
.Y(n_8924)
);

NAND2xp5_ASAP7_75t_L g8925 ( 
.A(n_8396),
.B(n_5204),
.Y(n_8925)
);

NAND2xp5_ASAP7_75t_L g8926 ( 
.A(n_8400),
.B(n_5205),
.Y(n_8926)
);

INVx1_ASAP7_75t_L g8927 ( 
.A(n_8401),
.Y(n_8927)
);

NAND2xp5_ASAP7_75t_SL g8928 ( 
.A(n_8450),
.B(n_8226),
.Y(n_8928)
);

NAND2xp5_ASAP7_75t_L g8929 ( 
.A(n_8411),
.B(n_5208),
.Y(n_8929)
);

AOI22xp5_ASAP7_75t_SL g8930 ( 
.A1(n_8281),
.A2(n_5211),
.B1(n_5212),
.B2(n_5210),
.Y(n_8930)
);

INVx1_ASAP7_75t_L g8931 ( 
.A(n_8420),
.Y(n_8931)
);

NAND2xp5_ASAP7_75t_SL g8932 ( 
.A(n_8696),
.B(n_5215),
.Y(n_8932)
);

NAND2xp5_ASAP7_75t_L g8933 ( 
.A(n_8424),
.B(n_5216),
.Y(n_8933)
);

INVx1_ASAP7_75t_L g8934 ( 
.A(n_8425),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_L g8935 ( 
.A(n_8444),
.B(n_5219),
.Y(n_8935)
);

NAND2xp5_ASAP7_75t_L g8936 ( 
.A(n_8447),
.B(n_8451),
.Y(n_8936)
);

INVx2_ASAP7_75t_L g8937 ( 
.A(n_8391),
.Y(n_8937)
);

INVx2_ASAP7_75t_SL g8938 ( 
.A(n_8426),
.Y(n_8938)
);

AOI22xp33_ASAP7_75t_L g8939 ( 
.A1(n_8362),
.A2(n_5224),
.B1(n_5226),
.B2(n_5221),
.Y(n_8939)
);

BUFx6f_ASAP7_75t_L g8940 ( 
.A(n_8282),
.Y(n_8940)
);

INVx1_ASAP7_75t_L g8941 ( 
.A(n_8452),
.Y(n_8941)
);

NOR3xp33_ASAP7_75t_L g8942 ( 
.A(n_8534),
.B(n_5338),
.C(n_5336),
.Y(n_8942)
);

NOR2xp33_ASAP7_75t_L g8943 ( 
.A(n_8427),
.B(n_5227),
.Y(n_8943)
);

NAND2xp5_ASAP7_75t_L g8944 ( 
.A(n_8465),
.B(n_5228),
.Y(n_8944)
);

OAI22xp33_ASAP7_75t_L g8945 ( 
.A1(n_8370),
.A2(n_8567),
.B1(n_8268),
.B2(n_8280),
.Y(n_8945)
);

NAND2xp5_ASAP7_75t_SL g8946 ( 
.A(n_8696),
.B(n_5229),
.Y(n_8946)
);

INVx1_ASAP7_75t_L g8947 ( 
.A(n_8466),
.Y(n_8947)
);

NAND2xp33_ASAP7_75t_L g8948 ( 
.A(n_8208),
.B(n_5234),
.Y(n_8948)
);

NAND2xp5_ASAP7_75t_SL g8949 ( 
.A(n_8282),
.B(n_5235),
.Y(n_8949)
);

INVx2_ASAP7_75t_SL g8950 ( 
.A(n_8426),
.Y(n_8950)
);

OR2x6_ASAP7_75t_L g8951 ( 
.A(n_8235),
.B(n_4907),
.Y(n_8951)
);

INVx1_ASAP7_75t_L g8952 ( 
.A(n_8472),
.Y(n_8952)
);

INVx2_ASAP7_75t_L g8953 ( 
.A(n_8393),
.Y(n_8953)
);

NAND2xp33_ASAP7_75t_L g8954 ( 
.A(n_8342),
.B(n_5237),
.Y(n_8954)
);

O2A1O1Ixp33_ASAP7_75t_L g8955 ( 
.A1(n_8573),
.A2(n_5350),
.B(n_5351),
.C(n_5348),
.Y(n_8955)
);

INVx1_ASAP7_75t_L g8956 ( 
.A(n_8473),
.Y(n_8956)
);

NOR2xp33_ASAP7_75t_L g8957 ( 
.A(n_8421),
.B(n_5239),
.Y(n_8957)
);

A2O1A1Ixp33_ASAP7_75t_L g8958 ( 
.A1(n_8563),
.A2(n_5358),
.B(n_5359),
.C(n_5356),
.Y(n_8958)
);

NOR2xp33_ASAP7_75t_L g8959 ( 
.A(n_8626),
.B(n_5241),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_8474),
.Y(n_8960)
);

INVx2_ASAP7_75t_L g8961 ( 
.A(n_8402),
.Y(n_8961)
);

INVx1_ASAP7_75t_L g8962 ( 
.A(n_8482),
.Y(n_8962)
);

INVxp67_ASAP7_75t_L g8963 ( 
.A(n_8678),
.Y(n_8963)
);

INVx1_ASAP7_75t_L g8964 ( 
.A(n_8487),
.Y(n_8964)
);

AND2x2_ASAP7_75t_L g8965 ( 
.A(n_8635),
.B(n_5243),
.Y(n_8965)
);

NAND2xp5_ASAP7_75t_SL g8966 ( 
.A(n_8296),
.B(n_5244),
.Y(n_8966)
);

INVxp67_ASAP7_75t_SL g8967 ( 
.A(n_8504),
.Y(n_8967)
);

NOR2xp33_ASAP7_75t_L g8968 ( 
.A(n_8243),
.B(n_5247),
.Y(n_8968)
);

NAND2xp5_ASAP7_75t_L g8969 ( 
.A(n_8493),
.B(n_8494),
.Y(n_8969)
);

AOI22xp5_ASAP7_75t_L g8970 ( 
.A1(n_8305),
.A2(n_5251),
.B1(n_5255),
.B2(n_5249),
.Y(n_8970)
);

NAND2xp5_ASAP7_75t_L g8971 ( 
.A(n_8495),
.B(n_5257),
.Y(n_8971)
);

NAND2xp5_ASAP7_75t_L g8972 ( 
.A(n_8501),
.B(n_5258),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_8507),
.Y(n_8973)
);

NAND2xp5_ASAP7_75t_L g8974 ( 
.A(n_8245),
.B(n_5265),
.Y(n_8974)
);

NAND2xp5_ASAP7_75t_L g8975 ( 
.A(n_8583),
.B(n_5269),
.Y(n_8975)
);

NAND2xp5_ASAP7_75t_SL g8976 ( 
.A(n_8296),
.B(n_5270),
.Y(n_8976)
);

NAND2xp33_ASAP7_75t_SL g8977 ( 
.A(n_8395),
.B(n_5277),
.Y(n_8977)
);

INVx2_ASAP7_75t_SL g8978 ( 
.A(n_8320),
.Y(n_8978)
);

AOI22xp5_ASAP7_75t_L g8979 ( 
.A1(n_8305),
.A2(n_5282),
.B1(n_5284),
.B2(n_5279),
.Y(n_8979)
);

INVx1_ASAP7_75t_L g8980 ( 
.A(n_8512),
.Y(n_8980)
);

NOR2xp33_ASAP7_75t_L g8981 ( 
.A(n_8266),
.B(n_5287),
.Y(n_8981)
);

NAND2xp5_ASAP7_75t_L g8982 ( 
.A(n_8514),
.B(n_5290),
.Y(n_8982)
);

AOI22xp5_ASAP7_75t_L g8983 ( 
.A1(n_8308),
.A2(n_5295),
.B1(n_5300),
.B2(n_5292),
.Y(n_8983)
);

NAND2xp5_ASAP7_75t_SL g8984 ( 
.A(n_8320),
.B(n_5301),
.Y(n_8984)
);

AND2x2_ASAP7_75t_L g8985 ( 
.A(n_8344),
.B(n_5304),
.Y(n_8985)
);

NAND2xp5_ASAP7_75t_L g8986 ( 
.A(n_8515),
.B(n_5308),
.Y(n_8986)
);

O2A1O1Ixp5_ASAP7_75t_L g8987 ( 
.A1(n_8706),
.A2(n_5367),
.B(n_5375),
.C(n_5365),
.Y(n_8987)
);

INVx2_ASAP7_75t_L g8988 ( 
.A(n_8405),
.Y(n_8988)
);

NAND2xp5_ASAP7_75t_L g8989 ( 
.A(n_8535),
.B(n_5311),
.Y(n_8989)
);

INVx1_ASAP7_75t_L g8990 ( 
.A(n_8536),
.Y(n_8990)
);

O2A1O1Ixp33_ASAP7_75t_L g8991 ( 
.A1(n_8513),
.A2(n_5402),
.B(n_5403),
.C(n_5390),
.Y(n_8991)
);

NAND2xp5_ASAP7_75t_L g8992 ( 
.A(n_8689),
.B(n_5314),
.Y(n_8992)
);

INVx3_ASAP7_75t_L g8993 ( 
.A(n_8328),
.Y(n_8993)
);

NAND2xp5_ASAP7_75t_L g8994 ( 
.A(n_8585),
.B(n_5315),
.Y(n_8994)
);

BUFx8_ASAP7_75t_L g8995 ( 
.A(n_8221),
.Y(n_8995)
);

AND2x6_ASAP7_75t_L g8996 ( 
.A(n_8646),
.B(n_5406),
.Y(n_8996)
);

INVx2_ASAP7_75t_L g8997 ( 
.A(n_8428),
.Y(n_8997)
);

AOI22xp33_ASAP7_75t_L g8998 ( 
.A1(n_8703),
.A2(n_8475),
.B1(n_8660),
.B2(n_8408),
.Y(n_8998)
);

NAND2xp5_ASAP7_75t_L g8999 ( 
.A(n_8598),
.B(n_5316),
.Y(n_8999)
);

INVx3_ASAP7_75t_L g9000 ( 
.A(n_8328),
.Y(n_9000)
);

NAND2x1_ASAP7_75t_L g9001 ( 
.A(n_8698),
.B(n_5407),
.Y(n_9001)
);

O2A1O1Ixp33_ASAP7_75t_L g9002 ( 
.A1(n_8609),
.A2(n_5409),
.B(n_5413),
.C(n_5408),
.Y(n_9002)
);

NAND2xp5_ASAP7_75t_SL g9003 ( 
.A(n_8338),
.B(n_5317),
.Y(n_9003)
);

O2A1O1Ixp33_ASAP7_75t_L g9004 ( 
.A1(n_8645),
.A2(n_5431),
.B(n_5440),
.C(n_5429),
.Y(n_9004)
);

NOR2xp33_ASAP7_75t_L g9005 ( 
.A(n_8311),
.B(n_5319),
.Y(n_9005)
);

NAND2xp5_ASAP7_75t_L g9006 ( 
.A(n_8568),
.B(n_5321),
.Y(n_9006)
);

NAND2xp5_ASAP7_75t_L g9007 ( 
.A(n_8471),
.B(n_5323),
.Y(n_9007)
);

HB1xp67_ASAP7_75t_L g9008 ( 
.A(n_8338),
.Y(n_9008)
);

NAND2xp5_ASAP7_75t_L g9009 ( 
.A(n_8625),
.B(n_5325),
.Y(n_9009)
);

NAND2xp5_ASAP7_75t_L g9010 ( 
.A(n_8683),
.B(n_5327),
.Y(n_9010)
);

AOI22xp33_ASAP7_75t_L g9011 ( 
.A1(n_8330),
.A2(n_5332),
.B1(n_5335),
.B2(n_5330),
.Y(n_9011)
);

NAND2xp5_ASAP7_75t_SL g9012 ( 
.A(n_8340),
.B(n_5339),
.Y(n_9012)
);

INVx2_ASAP7_75t_L g9013 ( 
.A(n_8429),
.Y(n_9013)
);

INVxp67_ASAP7_75t_L g9014 ( 
.A(n_8340),
.Y(n_9014)
);

INVx2_ASAP7_75t_L g9015 ( 
.A(n_8453),
.Y(n_9015)
);

NAND2xp5_ASAP7_75t_L g9016 ( 
.A(n_8647),
.B(n_5340),
.Y(n_9016)
);

INVx2_ASAP7_75t_L g9017 ( 
.A(n_8218),
.Y(n_9017)
);

INVx1_ASAP7_75t_L g9018 ( 
.A(n_8633),
.Y(n_9018)
);

INVx1_ASAP7_75t_L g9019 ( 
.A(n_8639),
.Y(n_9019)
);

NAND2xp5_ASAP7_75t_L g9020 ( 
.A(n_8375),
.B(n_5341),
.Y(n_9020)
);

AND2x6_ASAP7_75t_SL g9021 ( 
.A(n_8316),
.B(n_5445),
.Y(n_9021)
);

INVx2_ASAP7_75t_SL g9022 ( 
.A(n_8348),
.Y(n_9022)
);

BUFx3_ASAP7_75t_L g9023 ( 
.A(n_8313),
.Y(n_9023)
);

NAND2xp5_ASAP7_75t_L g9024 ( 
.A(n_8590),
.B(n_5342),
.Y(n_9024)
);

INVxp67_ASAP7_75t_L g9025 ( 
.A(n_8348),
.Y(n_9025)
);

NAND2xp5_ASAP7_75t_SL g9026 ( 
.A(n_8359),
.B(n_5343),
.Y(n_9026)
);

OAI22xp33_ASAP7_75t_L g9027 ( 
.A1(n_8319),
.A2(n_5347),
.B1(n_5349),
.B2(n_5344),
.Y(n_9027)
);

CKINVDCx5p33_ASAP7_75t_R g9028 ( 
.A(n_8353),
.Y(n_9028)
);

INVx1_ASAP7_75t_L g9029 ( 
.A(n_8623),
.Y(n_9029)
);

OR2x2_ASAP7_75t_L g9030 ( 
.A(n_8524),
.B(n_8423),
.Y(n_9030)
);

OAI221xp5_ASAP7_75t_L g9031 ( 
.A1(n_8531),
.A2(n_5455),
.B1(n_5470),
.B2(n_5453),
.C(n_5448),
.Y(n_9031)
);

NAND2xp5_ASAP7_75t_L g9032 ( 
.A(n_8392),
.B(n_8381),
.Y(n_9032)
);

NAND2xp5_ASAP7_75t_L g9033 ( 
.A(n_8250),
.B(n_5352),
.Y(n_9033)
);

AND2x2_ASAP7_75t_SL g9034 ( 
.A(n_8220),
.B(n_4953),
.Y(n_9034)
);

AOI22xp33_ASAP7_75t_L g9035 ( 
.A1(n_8345),
.A2(n_5354),
.B1(n_5357),
.B2(n_5353),
.Y(n_9035)
);

NAND2xp5_ASAP7_75t_SL g9036 ( 
.A(n_8359),
.B(n_5360),
.Y(n_9036)
);

OR2x2_ASAP7_75t_L g9037 ( 
.A(n_8510),
.B(n_5483),
.Y(n_9037)
);

NAND2xp5_ASAP7_75t_L g9038 ( 
.A(n_8409),
.B(n_8308),
.Y(n_9038)
);

INVx2_ASAP7_75t_L g9039 ( 
.A(n_8455),
.Y(n_9039)
);

NAND2xp5_ASAP7_75t_L g9040 ( 
.A(n_8409),
.B(n_5361),
.Y(n_9040)
);

NAND2xp5_ASAP7_75t_L g9041 ( 
.A(n_8688),
.B(n_5362),
.Y(n_9041)
);

NAND2xp5_ASAP7_75t_L g9042 ( 
.A(n_8589),
.B(n_5364),
.Y(n_9042)
);

AND2x6_ASAP7_75t_L g9043 ( 
.A(n_8624),
.B(n_5484),
.Y(n_9043)
);

OAI22xp5_ASAP7_75t_L g9044 ( 
.A1(n_8661),
.A2(n_5369),
.B1(n_5371),
.B2(n_5366),
.Y(n_9044)
);

NOR2xp33_ASAP7_75t_L g9045 ( 
.A(n_8572),
.B(n_5372),
.Y(n_9045)
);

NAND2xp5_ASAP7_75t_L g9046 ( 
.A(n_8628),
.B(n_5373),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_8538),
.Y(n_9047)
);

BUFx6f_ASAP7_75t_SL g9048 ( 
.A(n_8221),
.Y(n_9048)
);

INVx2_ASAP7_75t_L g9049 ( 
.A(n_8467),
.Y(n_9049)
);

NOR2xp33_ASAP7_75t_L g9050 ( 
.A(n_8549),
.B(n_5374),
.Y(n_9050)
);

INVx2_ASAP7_75t_L g9051 ( 
.A(n_8499),
.Y(n_9051)
);

AOI21xp5_ASAP7_75t_L g9052 ( 
.A1(n_8594),
.A2(n_5499),
.B(n_5492),
.Y(n_9052)
);

NAND2x1p5_ASAP7_75t_L g9053 ( 
.A(n_8407),
.B(n_5502),
.Y(n_9053)
);

INVx8_ASAP7_75t_L g9054 ( 
.A(n_8412),
.Y(n_9054)
);

NOR2xp67_ASAP7_75t_L g9055 ( 
.A(n_8326),
.B(n_3),
.Y(n_9055)
);

NOR2xp33_ASAP7_75t_L g9056 ( 
.A(n_8672),
.B(n_5376),
.Y(n_9056)
);

INVx1_ASAP7_75t_L g9057 ( 
.A(n_8541),
.Y(n_9057)
);

NAND2xp33_ASAP7_75t_L g9058 ( 
.A(n_8516),
.B(n_5377),
.Y(n_9058)
);

INVx2_ASAP7_75t_L g9059 ( 
.A(n_8502),
.Y(n_9059)
);

AND2x4_ASAP7_75t_L g9060 ( 
.A(n_8352),
.B(n_5508),
.Y(n_9060)
);

NOR2xp67_ASAP7_75t_L g9061 ( 
.A(n_8349),
.B(n_4),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_8545),
.Y(n_9062)
);

INVx1_ASAP7_75t_L g9063 ( 
.A(n_8550),
.Y(n_9063)
);

INVx2_ASAP7_75t_L g9064 ( 
.A(n_8508),
.Y(n_9064)
);

INVx3_ASAP7_75t_L g9065 ( 
.A(n_8360),
.Y(n_9065)
);

NOR2xp33_ASAP7_75t_L g9066 ( 
.A(n_8569),
.B(n_5378),
.Y(n_9066)
);

INVx2_ASAP7_75t_SL g9067 ( 
.A(n_8360),
.Y(n_9067)
);

INVx2_ASAP7_75t_L g9068 ( 
.A(n_8517),
.Y(n_9068)
);

INVx1_ASAP7_75t_L g9069 ( 
.A(n_8554),
.Y(n_9069)
);

OAI22xp5_ASAP7_75t_L g9070 ( 
.A1(n_8434),
.A2(n_5381),
.B1(n_5382),
.B2(n_5379),
.Y(n_9070)
);

AOI21xp5_ASAP7_75t_L g9071 ( 
.A1(n_8648),
.A2(n_5514),
.B(n_5512),
.Y(n_9071)
);

OR2x6_ASAP7_75t_L g9072 ( 
.A(n_8433),
.B(n_4981),
.Y(n_9072)
);

INVx2_ASAP7_75t_L g9073 ( 
.A(n_8523),
.Y(n_9073)
);

NOR2xp33_ASAP7_75t_L g9074 ( 
.A(n_8301),
.B(n_5384),
.Y(n_9074)
);

AND2x2_ASAP7_75t_L g9075 ( 
.A(n_8638),
.B(n_5387),
.Y(n_9075)
);

INVx2_ASAP7_75t_L g9076 ( 
.A(n_8525),
.Y(n_9076)
);

INVx2_ASAP7_75t_L g9077 ( 
.A(n_8528),
.Y(n_9077)
);

INVx1_ASAP7_75t_L g9078 ( 
.A(n_8555),
.Y(n_9078)
);

AND2x4_ASAP7_75t_L g9079 ( 
.A(n_8234),
.B(n_5515),
.Y(n_9079)
);

AND2x2_ASAP7_75t_SL g9080 ( 
.A(n_8239),
.B(n_4986),
.Y(n_9080)
);

AND2x2_ASAP7_75t_L g9081 ( 
.A(n_8479),
.B(n_5391),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_8559),
.Y(n_9082)
);

O2A1O1Ixp5_ASAP7_75t_L g9083 ( 
.A1(n_8674),
.A2(n_5522),
.B(n_5526),
.C(n_5516),
.Y(n_9083)
);

NAND2xp5_ASAP7_75t_SL g9084 ( 
.A(n_8378),
.B(n_5393),
.Y(n_9084)
);

INVx1_ASAP7_75t_L g9085 ( 
.A(n_8560),
.Y(n_9085)
);

OR2x2_ASAP7_75t_L g9086 ( 
.A(n_8440),
.B(n_5529),
.Y(n_9086)
);

NAND2xp5_ASAP7_75t_L g9087 ( 
.A(n_8422),
.B(n_5396),
.Y(n_9087)
);

NAND2xp5_ASAP7_75t_SL g9088 ( 
.A(n_8378),
.B(n_5397),
.Y(n_9088)
);

NAND2xp5_ASAP7_75t_SL g9089 ( 
.A(n_8388),
.B(n_5398),
.Y(n_9089)
);

NOR2xp33_ASAP7_75t_L g9090 ( 
.A(n_8306),
.B(n_8670),
.Y(n_9090)
);

INVx1_ASAP7_75t_L g9091 ( 
.A(n_8561),
.Y(n_9091)
);

NAND2xp5_ASAP7_75t_L g9092 ( 
.A(n_8416),
.B(n_5399),
.Y(n_9092)
);

INVx1_ASAP7_75t_L g9093 ( 
.A(n_8562),
.Y(n_9093)
);

OAI22xp5_ASAP7_75t_L g9094 ( 
.A1(n_8470),
.A2(n_5401),
.B1(n_5404),
.B2(n_5400),
.Y(n_9094)
);

NOR2xp33_ASAP7_75t_L g9095 ( 
.A(n_8270),
.B(n_5405),
.Y(n_9095)
);

INVx2_ASAP7_75t_L g9096 ( 
.A(n_8530),
.Y(n_9096)
);

NAND2xp5_ASAP7_75t_L g9097 ( 
.A(n_8435),
.B(n_5410),
.Y(n_9097)
);

INVxp33_ASAP7_75t_SL g9098 ( 
.A(n_8404),
.Y(n_9098)
);

NOR2xp33_ASAP7_75t_L g9099 ( 
.A(n_8388),
.B(n_5411),
.Y(n_9099)
);

INVx1_ASAP7_75t_L g9100 ( 
.A(n_8564),
.Y(n_9100)
);

NAND2xp5_ASAP7_75t_L g9101 ( 
.A(n_8620),
.B(n_5412),
.Y(n_9101)
);

NAND2xp5_ASAP7_75t_L g9102 ( 
.A(n_8620),
.B(n_8680),
.Y(n_9102)
);

A2O1A1Ixp33_ASAP7_75t_L g9103 ( 
.A1(n_8607),
.A2(n_5537),
.B(n_5533),
.C(n_5103),
.Y(n_9103)
);

BUFx8_ASAP7_75t_L g9104 ( 
.A(n_8469),
.Y(n_9104)
);

INVx2_ASAP7_75t_L g9105 ( 
.A(n_8533),
.Y(n_9105)
);

XOR2xp5_ASAP7_75t_L g9106 ( 
.A(n_8294),
.B(n_5414),
.Y(n_9106)
);

INVx3_ASAP7_75t_L g9107 ( 
.A(n_8443),
.Y(n_9107)
);

INVx1_ASAP7_75t_L g9108 ( 
.A(n_8579),
.Y(n_9108)
);

AND2x2_ASAP7_75t_L g9109 ( 
.A(n_8480),
.B(n_5415),
.Y(n_9109)
);

NAND2xp5_ASAP7_75t_L g9110 ( 
.A(n_8443),
.B(n_5416),
.Y(n_9110)
);

NAND2xp5_ASAP7_75t_L g9111 ( 
.A(n_8692),
.B(n_5417),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_8581),
.Y(n_9112)
);

INVx1_ASAP7_75t_L g9113 ( 
.A(n_8597),
.Y(n_9113)
);

NAND2xp5_ASAP7_75t_L g9114 ( 
.A(n_8602),
.B(n_8617),
.Y(n_9114)
);

AOI22xp33_ASAP7_75t_L g9115 ( 
.A1(n_8586),
.A2(n_5423),
.B1(n_5424),
.B2(n_5418),
.Y(n_9115)
);

NOR2xp33_ASAP7_75t_L g9116 ( 
.A(n_8285),
.B(n_5425),
.Y(n_9116)
);

NAND2xp5_ASAP7_75t_SL g9117 ( 
.A(n_8666),
.B(n_5426),
.Y(n_9117)
);

BUFx2_ASAP7_75t_L g9118 ( 
.A(n_8463),
.Y(n_9118)
);

AND2x2_ASAP7_75t_L g9119 ( 
.A(n_8442),
.B(n_5430),
.Y(n_9119)
);

INVxp67_ASAP7_75t_SL g9120 ( 
.A(n_8491),
.Y(n_9120)
);

NAND3xp33_ASAP7_75t_L g9121 ( 
.A(n_8656),
.B(n_5433),
.C(n_5432),
.Y(n_9121)
);

BUFx6f_ASAP7_75t_L g9122 ( 
.A(n_8496),
.Y(n_9122)
);

AO221x1_ASAP7_75t_L g9123 ( 
.A1(n_8380),
.A2(n_5129),
.B1(n_5134),
.B2(n_5109),
.C(n_5081),
.Y(n_9123)
);

NAND2xp5_ASAP7_75t_SL g9124 ( 
.A(n_8666),
.B(n_5434),
.Y(n_9124)
);

INVx2_ASAP7_75t_SL g9125 ( 
.A(n_8412),
.Y(n_9125)
);

INVx8_ASAP7_75t_L g9126 ( 
.A(n_8469),
.Y(n_9126)
);

NAND2xp5_ASAP7_75t_SL g9127 ( 
.A(n_8676),
.B(n_5435),
.Y(n_9127)
);

NAND2xp5_ASAP7_75t_L g9128 ( 
.A(n_8667),
.B(n_5436),
.Y(n_9128)
);

INVx1_ASAP7_75t_L g9129 ( 
.A(n_8668),
.Y(n_9129)
);

OAI22xp5_ASAP7_75t_L g9130 ( 
.A1(n_8477),
.A2(n_5439),
.B1(n_5442),
.B2(n_5437),
.Y(n_9130)
);

NOR2xp33_ASAP7_75t_L g9131 ( 
.A(n_8613),
.B(n_5443),
.Y(n_9131)
);

INVx2_ASAP7_75t_SL g9132 ( 
.A(n_8532),
.Y(n_9132)
);

NAND2xp5_ASAP7_75t_L g9133 ( 
.A(n_8679),
.B(n_8484),
.Y(n_9133)
);

INVxp67_ASAP7_75t_SL g9134 ( 
.A(n_8520),
.Y(n_9134)
);

INVx2_ASAP7_75t_L g9135 ( 
.A(n_8547),
.Y(n_9135)
);

INVx3_ASAP7_75t_L g9136 ( 
.A(n_8410),
.Y(n_9136)
);

INVx1_ASAP7_75t_L g9137 ( 
.A(n_8552),
.Y(n_9137)
);

INVx3_ASAP7_75t_L g9138 ( 
.A(n_8432),
.Y(n_9138)
);

NAND2xp5_ASAP7_75t_SL g9139 ( 
.A(n_8676),
.B(n_5446),
.Y(n_9139)
);

NAND2xp5_ASAP7_75t_SL g9140 ( 
.A(n_8519),
.B(n_5447),
.Y(n_9140)
);

INVx1_ASAP7_75t_L g9141 ( 
.A(n_8556),
.Y(n_9141)
);

AO221x1_ASAP7_75t_L g9142 ( 
.A1(n_8379),
.A2(n_5163),
.B1(n_5167),
.B2(n_5140),
.C(n_5139),
.Y(n_9142)
);

BUFx6f_ASAP7_75t_L g9143 ( 
.A(n_8496),
.Y(n_9143)
);

AND2x2_ASAP7_75t_L g9144 ( 
.A(n_8366),
.B(n_5449),
.Y(n_9144)
);

AND2x2_ASAP7_75t_L g9145 ( 
.A(n_8397),
.B(n_5450),
.Y(n_9145)
);

NOR2xp33_ASAP7_75t_L g9146 ( 
.A(n_8553),
.B(n_8695),
.Y(n_9146)
);

NOR2xp33_ASAP7_75t_L g9147 ( 
.A(n_8213),
.B(n_5451),
.Y(n_9147)
);

INVx2_ASAP7_75t_L g9148 ( 
.A(n_8580),
.Y(n_9148)
);

NAND2xp5_ASAP7_75t_L g9149 ( 
.A(n_8654),
.B(n_5452),
.Y(n_9149)
);

NAND2xp5_ASAP7_75t_L g9150 ( 
.A(n_8544),
.B(n_5454),
.Y(n_9150)
);

INVx2_ASAP7_75t_SL g9151 ( 
.A(n_8578),
.Y(n_9151)
);

INVx2_ASAP7_75t_L g9152 ( 
.A(n_8582),
.Y(n_9152)
);

INVx2_ASAP7_75t_L g9153 ( 
.A(n_8592),
.Y(n_9153)
);

NOR2xp33_ASAP7_75t_L g9154 ( 
.A(n_8681),
.B(n_5456),
.Y(n_9154)
);

NOR2xp33_ASAP7_75t_L g9155 ( 
.A(n_8399),
.B(n_5458),
.Y(n_9155)
);

INVx2_ASAP7_75t_L g9156 ( 
.A(n_8595),
.Y(n_9156)
);

NAND2xp5_ASAP7_75t_SL g9157 ( 
.A(n_8519),
.B(n_5459),
.Y(n_9157)
);

NAND2xp5_ASAP7_75t_SL g9158 ( 
.A(n_8565),
.B(n_5461),
.Y(n_9158)
);

AOI22xp5_ASAP7_75t_L g9159 ( 
.A1(n_8457),
.A2(n_5465),
.B1(n_5466),
.B2(n_5463),
.Y(n_9159)
);

AOI22xp33_ASAP7_75t_L g9160 ( 
.A1(n_8438),
.A2(n_5471),
.B1(n_5473),
.B2(n_5469),
.Y(n_9160)
);

INVx2_ASAP7_75t_SL g9161 ( 
.A(n_8591),
.Y(n_9161)
);

NOR2xp33_ASAP7_75t_L g9162 ( 
.A(n_8468),
.B(n_5474),
.Y(n_9162)
);

AND2x2_ASAP7_75t_L g9163 ( 
.A(n_8694),
.B(n_5475),
.Y(n_9163)
);

NAND2xp5_ASAP7_75t_SL g9164 ( 
.A(n_8565),
.B(n_8596),
.Y(n_9164)
);

AND2x2_ASAP7_75t_L g9165 ( 
.A(n_8619),
.B(n_5476),
.Y(n_9165)
);

INVx2_ASAP7_75t_L g9166 ( 
.A(n_8600),
.Y(n_9166)
);

NAND2xp5_ASAP7_75t_SL g9167 ( 
.A(n_8596),
.B(n_5477),
.Y(n_9167)
);

AOI22xp33_ASAP7_75t_L g9168 ( 
.A1(n_8606),
.A2(n_5480),
.B1(n_5486),
.B2(n_5479),
.Y(n_9168)
);

CKINVDCx14_ASAP7_75t_R g9169 ( 
.A(n_8642),
.Y(n_9169)
);

NAND2xp5_ASAP7_75t_L g9170 ( 
.A(n_8637),
.B(n_5487),
.Y(n_9170)
);

INVxp67_ASAP7_75t_L g9171 ( 
.A(n_8599),
.Y(n_9171)
);

AOI22xp5_ASAP7_75t_L g9172 ( 
.A1(n_8518),
.A2(n_8481),
.B1(n_8215),
.B2(n_8490),
.Y(n_9172)
);

NOR2xp67_ASAP7_75t_L g9173 ( 
.A(n_8454),
.B(n_4),
.Y(n_9173)
);

AOI22xp33_ASAP7_75t_L g9174 ( 
.A1(n_8612),
.A2(n_5489),
.B1(n_5491),
.B2(n_5488),
.Y(n_9174)
);

CKINVDCx5p33_ASAP7_75t_R g9175 ( 
.A(n_8290),
.Y(n_9175)
);

A2O1A1Ixp33_ASAP7_75t_L g9176 ( 
.A1(n_8500),
.A2(n_8542),
.B(n_8657),
.C(n_8697),
.Y(n_9176)
);

INVx2_ASAP7_75t_L g9177 ( 
.A(n_8614),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_8621),
.Y(n_9178)
);

NAND2xp5_ASAP7_75t_L g9179 ( 
.A(n_8643),
.B(n_5493),
.Y(n_9179)
);

INVx1_ASAP7_75t_L g9180 ( 
.A(n_8662),
.Y(n_9180)
);

NOR3xp33_ASAP7_75t_L g9181 ( 
.A(n_8685),
.B(n_5174),
.C(n_5168),
.Y(n_9181)
);

INVx2_ASAP7_75t_L g9182 ( 
.A(n_8669),
.Y(n_9182)
);

INVx4_ASAP7_75t_L g9183 ( 
.A(n_8382),
.Y(n_9183)
);

NOR2xp33_ASAP7_75t_L g9184 ( 
.A(n_8485),
.B(n_5495),
.Y(n_9184)
);

NAND2xp5_ASAP7_75t_SL g9185 ( 
.A(n_8599),
.B(n_5505),
.Y(n_9185)
);

NAND2xp5_ASAP7_75t_L g9186 ( 
.A(n_8673),
.B(n_5507),
.Y(n_9186)
);

NAND2xp5_ASAP7_75t_SL g9187 ( 
.A(n_8605),
.B(n_5509),
.Y(n_9187)
);

NOR2xp33_ASAP7_75t_L g9188 ( 
.A(n_8691),
.B(n_5192),
.Y(n_9188)
);

A2O1A1Ixp33_ASAP7_75t_L g9189 ( 
.A1(n_8489),
.A2(n_5242),
.B(n_5246),
.C(n_5202),
.Y(n_9189)
);

O2A1O1Ixp33_ASAP7_75t_L g9190 ( 
.A1(n_8701),
.A2(n_5370),
.B(n_5385),
.C(n_5253),
.Y(n_9190)
);

NAND2xp5_ASAP7_75t_SL g9191 ( 
.A(n_8605),
.B(n_5394),
.Y(n_9191)
);

INVx1_ASAP7_75t_L g9192 ( 
.A(n_8677),
.Y(n_9192)
);

AND2x2_ASAP7_75t_L g9193 ( 
.A(n_8603),
.B(n_5395),
.Y(n_9193)
);

INVx1_ASAP7_75t_L g9194 ( 
.A(n_8693),
.Y(n_9194)
);

NAND2xp5_ASAP7_75t_SL g9195 ( 
.A(n_8610),
.B(n_5419),
.Y(n_9195)
);

NAND2xp5_ASAP7_75t_L g9196 ( 
.A(n_8611),
.B(n_5420),
.Y(n_9196)
);

AND2x2_ASAP7_75t_L g9197 ( 
.A(n_8540),
.B(n_5428),
.Y(n_9197)
);

NAND3xp33_ASAP7_75t_L g9198 ( 
.A(n_8699),
.B(n_5441),
.C(n_5438),
.Y(n_9198)
);

INVx1_ASAP7_75t_L g9199 ( 
.A(n_8700),
.Y(n_9199)
);

INVx2_ASAP7_75t_L g9200 ( 
.A(n_8705),
.Y(n_9200)
);

NAND2xp33_ASAP7_75t_L g9201 ( 
.A(n_8458),
.B(n_5478),
.Y(n_9201)
);

NAND2xp5_ASAP7_75t_L g9202 ( 
.A(n_8506),
.B(n_5506),
.Y(n_9202)
);

OR2x2_ASAP7_75t_L g9203 ( 
.A(n_8566),
.B(n_5517),
.Y(n_9203)
);

INVx2_ASAP7_75t_SL g9204 ( 
.A(n_8610),
.Y(n_9204)
);

NAND2xp5_ASAP7_75t_L g9205 ( 
.A(n_8574),
.B(n_5523),
.Y(n_9205)
);

INVx2_ASAP7_75t_L g9206 ( 
.A(n_8710),
.Y(n_9206)
);

AOI22xp33_ASAP7_75t_L g9207 ( 
.A1(n_8518),
.A2(n_5545),
.B1(n_5524),
.B2(n_6),
.Y(n_9207)
);

AOI22xp5_ASAP7_75t_L g9208 ( 
.A1(n_8275),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_9208)
);

NAND2xp5_ASAP7_75t_L g9209 ( 
.A(n_8571),
.B(n_5),
.Y(n_9209)
);

NAND2xp5_ASAP7_75t_L g9210 ( 
.A(n_8575),
.B(n_6),
.Y(n_9210)
);

AOI22xp33_ASAP7_75t_SL g9211 ( 
.A1(n_8717),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_9211)
);

INVxp67_ASAP7_75t_L g9212 ( 
.A(n_8615),
.Y(n_9212)
);

NAND2xp5_ASAP7_75t_L g9213 ( 
.A(n_8616),
.B(n_7),
.Y(n_9213)
);

NAND2xp5_ASAP7_75t_L g9214 ( 
.A(n_8651),
.B(n_7),
.Y(n_9214)
);

INVx1_ASAP7_75t_L g9215 ( 
.A(n_8714),
.Y(n_9215)
);

NAND2xp5_ASAP7_75t_SL g9216 ( 
.A(n_8615),
.B(n_123),
.Y(n_9216)
);

NAND2xp5_ASAP7_75t_L g9217 ( 
.A(n_8636),
.B(n_8),
.Y(n_9217)
);

INVx2_ASAP7_75t_L g9218 ( 
.A(n_8636),
.Y(n_9218)
);

INVxp67_ASAP7_75t_L g9219 ( 
.A(n_8641),
.Y(n_9219)
);

NAND2xp5_ASAP7_75t_L g9220 ( 
.A(n_8641),
.B(n_8),
.Y(n_9220)
);

NAND2xp5_ASAP7_75t_L g9221 ( 
.A(n_8649),
.B(n_8577),
.Y(n_9221)
);

AOI22xp33_ASAP7_75t_L g9222 ( 
.A1(n_8460),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_9222)
);

AOI22xp5_ASAP7_75t_L g9223 ( 
.A1(n_8449),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_9223)
);

AOI21xp5_ASAP7_75t_L g9224 ( 
.A1(n_8716),
.A2(n_124),
.B(n_123),
.Y(n_9224)
);

NAND2xp5_ASAP7_75t_L g9225 ( 
.A(n_8649),
.B(n_11),
.Y(n_9225)
);

INVx1_ASAP7_75t_L g9226 ( 
.A(n_8608),
.Y(n_9226)
);

INVx2_ASAP7_75t_L g9227 ( 
.A(n_8587),
.Y(n_9227)
);

NAND3xp33_ASAP7_75t_L g9228 ( 
.A(n_8505),
.B(n_12),
.C(n_13),
.Y(n_9228)
);

NAND2xp5_ASAP7_75t_L g9229 ( 
.A(n_8588),
.B(n_13),
.Y(n_9229)
);

AO22x2_ASAP7_75t_L g9230 ( 
.A1(n_8333),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_9230)
);

INVx2_ASAP7_75t_L g9231 ( 
.A(n_8640),
.Y(n_9231)
);

NOR2xp67_ASAP7_75t_L g9232 ( 
.A(n_8675),
.B(n_14),
.Y(n_9232)
);

INVx1_ASAP7_75t_L g9233 ( 
.A(n_8658),
.Y(n_9233)
);

INVx2_ASAP7_75t_L g9234 ( 
.A(n_8337),
.Y(n_9234)
);

INVx2_ASAP7_75t_L g9235 ( 
.A(n_8341),
.Y(n_9235)
);

AOI22xp33_ASAP7_75t_L g9236 ( 
.A1(n_8386),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_9236)
);

NAND2xp5_ASAP7_75t_L g9237 ( 
.A(n_8729),
.B(n_8247),
.Y(n_9237)
);

AND2x2_ASAP7_75t_L g9238 ( 
.A(n_8732),
.B(n_8413),
.Y(n_9238)
);

NAND2xp5_ASAP7_75t_SL g9239 ( 
.A(n_9034),
.B(n_8262),
.Y(n_9239)
);

INVxp67_ASAP7_75t_L g9240 ( 
.A(n_8787),
.Y(n_9240)
);

INVx2_ASAP7_75t_L g9241 ( 
.A(n_8723),
.Y(n_9241)
);

HB1xp67_ASAP7_75t_L g9242 ( 
.A(n_8830),
.Y(n_9242)
);

INVx3_ASAP7_75t_L g9243 ( 
.A(n_8820),
.Y(n_9243)
);

HB1xp67_ASAP7_75t_L g9244 ( 
.A(n_8826),
.Y(n_9244)
);

BUFx3_ASAP7_75t_L g9245 ( 
.A(n_9054),
.Y(n_9245)
);

AND2x4_ASAP7_75t_L g9246 ( 
.A(n_8899),
.B(n_8264),
.Y(n_9246)
);

INVx1_ASAP7_75t_L g9247 ( 
.A(n_8889),
.Y(n_9247)
);

HB1xp67_ASAP7_75t_L g9248 ( 
.A(n_8890),
.Y(n_9248)
);

HB1xp67_ASAP7_75t_L g9249 ( 
.A(n_8746),
.Y(n_9249)
);

AND2x2_ASAP7_75t_L g9250 ( 
.A(n_8965),
.B(n_124),
.Y(n_9250)
);

NOR2xp67_ASAP7_75t_L g9251 ( 
.A(n_9090),
.B(n_16),
.Y(n_9251)
);

INVx1_ASAP7_75t_SL g9252 ( 
.A(n_9098),
.Y(n_9252)
);

AND2x2_ASAP7_75t_L g9253 ( 
.A(n_8985),
.B(n_9075),
.Y(n_9253)
);

HB1xp67_ASAP7_75t_L g9254 ( 
.A(n_8894),
.Y(n_9254)
);

INVx2_ASAP7_75t_L g9255 ( 
.A(n_8735),
.Y(n_9255)
);

INVx2_ASAP7_75t_SL g9256 ( 
.A(n_8820),
.Y(n_9256)
);

HB1xp67_ASAP7_75t_L g9257 ( 
.A(n_8936),
.Y(n_9257)
);

OAI21xp5_ASAP7_75t_L g9258 ( 
.A1(n_9131),
.A2(n_9056),
.B(n_8957),
.Y(n_9258)
);

NAND2xp5_ASAP7_75t_L g9259 ( 
.A(n_8769),
.B(n_17),
.Y(n_9259)
);

NAND2xp5_ASAP7_75t_SL g9260 ( 
.A(n_8719),
.B(n_125),
.Y(n_9260)
);

INVx1_ASAP7_75t_SL g9261 ( 
.A(n_9118),
.Y(n_9261)
);

INVx2_ASAP7_75t_L g9262 ( 
.A(n_8736),
.Y(n_9262)
);

NAND2xp5_ASAP7_75t_L g9263 ( 
.A(n_8724),
.B(n_17),
.Y(n_9263)
);

AND2x2_ASAP7_75t_L g9264 ( 
.A(n_8873),
.B(n_9080),
.Y(n_9264)
);

INVx2_ASAP7_75t_L g9265 ( 
.A(n_8756),
.Y(n_9265)
);

AND2x6_ASAP7_75t_L g9266 ( 
.A(n_9226),
.B(n_18),
.Y(n_9266)
);

INVx3_ASAP7_75t_L g9267 ( 
.A(n_8848),
.Y(n_9267)
);

NAND2xp5_ASAP7_75t_SL g9268 ( 
.A(n_8868),
.B(n_125),
.Y(n_9268)
);

INVx4_ASAP7_75t_L g9269 ( 
.A(n_9175),
.Y(n_9269)
);

AND2x4_ASAP7_75t_L g9270 ( 
.A(n_8923),
.B(n_126),
.Y(n_9270)
);

INVx2_ASAP7_75t_SL g9271 ( 
.A(n_9054),
.Y(n_9271)
);

AND2x2_ASAP7_75t_L g9272 ( 
.A(n_8852),
.B(n_8763),
.Y(n_9272)
);

INVx1_ASAP7_75t_L g9273 ( 
.A(n_8969),
.Y(n_9273)
);

AND2x2_ASAP7_75t_L g9274 ( 
.A(n_9165),
.B(n_126),
.Y(n_9274)
);

OAI21xp5_ASAP7_75t_L g9275 ( 
.A1(n_8968),
.A2(n_18),
.B(n_19),
.Y(n_9275)
);

INVx1_ASAP7_75t_L g9276 ( 
.A(n_8734),
.Y(n_9276)
);

AND2x2_ASAP7_75t_L g9277 ( 
.A(n_9193),
.B(n_127),
.Y(n_9277)
);

INVx1_ASAP7_75t_L g9278 ( 
.A(n_8742),
.Y(n_9278)
);

AND2x2_ASAP7_75t_SL g9279 ( 
.A(n_8775),
.B(n_18),
.Y(n_9279)
);

INVx1_ASAP7_75t_L g9280 ( 
.A(n_8752),
.Y(n_9280)
);

INVx3_ASAP7_75t_L g9281 ( 
.A(n_8848),
.Y(n_9281)
);

INVx1_ASAP7_75t_L g9282 ( 
.A(n_8765),
.Y(n_9282)
);

INVx3_ASAP7_75t_L g9283 ( 
.A(n_8862),
.Y(n_9283)
);

INVx1_ASAP7_75t_SL g9284 ( 
.A(n_8862),
.Y(n_9284)
);

AND2x2_ASAP7_75t_L g9285 ( 
.A(n_9230),
.B(n_127),
.Y(n_9285)
);

HB1xp67_ASAP7_75t_L g9286 ( 
.A(n_8767),
.Y(n_9286)
);

BUFx6f_ASAP7_75t_L g9287 ( 
.A(n_9023),
.Y(n_9287)
);

NAND2x1p5_ASAP7_75t_L g9288 ( 
.A(n_8799),
.B(n_128),
.Y(n_9288)
);

AND2x2_ASAP7_75t_L g9289 ( 
.A(n_9230),
.B(n_128),
.Y(n_9289)
);

HB1xp67_ASAP7_75t_L g9290 ( 
.A(n_8771),
.Y(n_9290)
);

INVx2_ASAP7_75t_L g9291 ( 
.A(n_8757),
.Y(n_9291)
);

INVx2_ASAP7_75t_L g9292 ( 
.A(n_8761),
.Y(n_9292)
);

AND2x2_ASAP7_75t_L g9293 ( 
.A(n_8738),
.B(n_129),
.Y(n_9293)
);

AND2x2_ASAP7_75t_L g9294 ( 
.A(n_9197),
.B(n_129),
.Y(n_9294)
);

HB1xp67_ASAP7_75t_L g9295 ( 
.A(n_8772),
.Y(n_9295)
);

AND2x2_ASAP7_75t_SL g9296 ( 
.A(n_8829),
.B(n_19),
.Y(n_9296)
);

INVx1_ASAP7_75t_L g9297 ( 
.A(n_8777),
.Y(n_9297)
);

NAND2xp5_ASAP7_75t_L g9298 ( 
.A(n_8996),
.B(n_20),
.Y(n_9298)
);

INVx2_ASAP7_75t_L g9299 ( 
.A(n_8776),
.Y(n_9299)
);

AND2x4_ASAP7_75t_L g9300 ( 
.A(n_8720),
.B(n_130),
.Y(n_9300)
);

INVx1_ASAP7_75t_L g9301 ( 
.A(n_8786),
.Y(n_9301)
);

INVx1_ASAP7_75t_L g9302 ( 
.A(n_8791),
.Y(n_9302)
);

INVx3_ASAP7_75t_L g9303 ( 
.A(n_8940),
.Y(n_9303)
);

INVx1_ASAP7_75t_L g9304 ( 
.A(n_8805),
.Y(n_9304)
);

INVx2_ASAP7_75t_L g9305 ( 
.A(n_8781),
.Y(n_9305)
);

AND2x2_ASAP7_75t_L g9306 ( 
.A(n_8857),
.B(n_130),
.Y(n_9306)
);

BUFx6f_ASAP7_75t_L g9307 ( 
.A(n_9122),
.Y(n_9307)
);

INVx2_ASAP7_75t_L g9308 ( 
.A(n_8795),
.Y(n_9308)
);

OR2x6_ASAP7_75t_L g9309 ( 
.A(n_8730),
.B(n_9126),
.Y(n_9309)
);

INVx2_ASAP7_75t_L g9310 ( 
.A(n_8803),
.Y(n_9310)
);

NAND2xp5_ASAP7_75t_L g9311 ( 
.A(n_8996),
.B(n_20),
.Y(n_9311)
);

AND2x2_ASAP7_75t_L g9312 ( 
.A(n_9037),
.B(n_131),
.Y(n_9312)
);

AND2x2_ASAP7_75t_L g9313 ( 
.A(n_8727),
.B(n_131),
.Y(n_9313)
);

AND2x2_ASAP7_75t_L g9314 ( 
.A(n_8885),
.B(n_132),
.Y(n_9314)
);

AND2x2_ASAP7_75t_L g9315 ( 
.A(n_8930),
.B(n_133),
.Y(n_9315)
);

NOR2xp33_ASAP7_75t_L g9316 ( 
.A(n_8943),
.B(n_133),
.Y(n_9316)
);

AND2x4_ASAP7_75t_L g9317 ( 
.A(n_8812),
.B(n_134),
.Y(n_9317)
);

BUFx3_ASAP7_75t_L g9318 ( 
.A(n_8730),
.Y(n_9318)
);

AND2x2_ASAP7_75t_L g9319 ( 
.A(n_8919),
.B(n_9030),
.Y(n_9319)
);

INVx2_ASAP7_75t_SL g9320 ( 
.A(n_8940),
.Y(n_9320)
);

AND2x2_ASAP7_75t_L g9321 ( 
.A(n_9163),
.B(n_134),
.Y(n_9321)
);

AND2x4_ASAP7_75t_L g9322 ( 
.A(n_8754),
.B(n_135),
.Y(n_9322)
);

AND2x2_ASAP7_75t_L g9323 ( 
.A(n_9081),
.B(n_135),
.Y(n_9323)
);

AND2x2_ASAP7_75t_L g9324 ( 
.A(n_9109),
.B(n_136),
.Y(n_9324)
);

INVx2_ASAP7_75t_L g9325 ( 
.A(n_8828),
.Y(n_9325)
);

AND2x2_ASAP7_75t_L g9326 ( 
.A(n_8998),
.B(n_136),
.Y(n_9326)
);

OAI21xp5_ASAP7_75t_L g9327 ( 
.A1(n_9050),
.A2(n_20),
.B(n_21),
.Y(n_9327)
);

AND2x2_ASAP7_75t_L g9328 ( 
.A(n_9008),
.B(n_137),
.Y(n_9328)
);

NAND2xp5_ASAP7_75t_SL g9329 ( 
.A(n_8740),
.B(n_137),
.Y(n_9329)
);

AND2x6_ASAP7_75t_L g9330 ( 
.A(n_8810),
.B(n_21),
.Y(n_9330)
);

BUFx6f_ASAP7_75t_L g9331 ( 
.A(n_9122),
.Y(n_9331)
);

NAND2xp5_ASAP7_75t_L g9332 ( 
.A(n_8996),
.B(n_21),
.Y(n_9332)
);

INVx2_ASAP7_75t_L g9333 ( 
.A(n_8831),
.Y(n_9333)
);

BUFx6f_ASAP7_75t_L g9334 ( 
.A(n_9143),
.Y(n_9334)
);

INVx1_ASAP7_75t_L g9335 ( 
.A(n_8824),
.Y(n_9335)
);

INVx2_ASAP7_75t_L g9336 ( 
.A(n_8835),
.Y(n_9336)
);

INVx1_ASAP7_75t_L g9337 ( 
.A(n_8844),
.Y(n_9337)
);

INVx2_ASAP7_75t_L g9338 ( 
.A(n_8842),
.Y(n_9338)
);

INVx2_ASAP7_75t_L g9339 ( 
.A(n_8845),
.Y(n_9339)
);

BUFx3_ASAP7_75t_L g9340 ( 
.A(n_9143),
.Y(n_9340)
);

BUFx8_ASAP7_75t_L g9341 ( 
.A(n_9048),
.Y(n_9341)
);

INVx2_ASAP7_75t_SL g9342 ( 
.A(n_8993),
.Y(n_9342)
);

NAND2xp5_ASAP7_75t_SL g9343 ( 
.A(n_8758),
.B(n_138),
.Y(n_9343)
);

AND2x2_ASAP7_75t_L g9344 ( 
.A(n_8748),
.B(n_138),
.Y(n_9344)
);

INVx2_ASAP7_75t_L g9345 ( 
.A(n_8861),
.Y(n_9345)
);

BUFx3_ASAP7_75t_L g9346 ( 
.A(n_8995),
.Y(n_9346)
);

NAND2xp5_ASAP7_75t_SL g9347 ( 
.A(n_8758),
.B(n_8743),
.Y(n_9347)
);

INVx8_ASAP7_75t_L g9348 ( 
.A(n_9126),
.Y(n_9348)
);

AND2x6_ASAP7_75t_L g9349 ( 
.A(n_8855),
.B(n_22),
.Y(n_9349)
);

NOR2xp33_ASAP7_75t_L g9350 ( 
.A(n_8836),
.B(n_139),
.Y(n_9350)
);

NAND2xp5_ASAP7_75t_L g9351 ( 
.A(n_8963),
.B(n_22),
.Y(n_9351)
);

AND2x2_ASAP7_75t_L g9352 ( 
.A(n_8928),
.B(n_139),
.Y(n_9352)
);

INVx1_ASAP7_75t_L g9353 ( 
.A(n_8871),
.Y(n_9353)
);

AND2x2_ASAP7_75t_L g9354 ( 
.A(n_9145),
.B(n_140),
.Y(n_9354)
);

AND2x2_ASAP7_75t_L g9355 ( 
.A(n_9000),
.B(n_140),
.Y(n_9355)
);

NAND2xp5_ASAP7_75t_SL g9356 ( 
.A(n_8758),
.B(n_141),
.Y(n_9356)
);

NAND2xp5_ASAP7_75t_L g9357 ( 
.A(n_8731),
.B(n_22),
.Y(n_9357)
);

AND2x2_ASAP7_75t_L g9358 ( 
.A(n_9065),
.B(n_9107),
.Y(n_9358)
);

INVx2_ASAP7_75t_SL g9359 ( 
.A(n_8846),
.Y(n_9359)
);

AND2x2_ASAP7_75t_L g9360 ( 
.A(n_8860),
.B(n_142),
.Y(n_9360)
);

AND2x2_ASAP7_75t_L g9361 ( 
.A(n_8816),
.B(n_142),
.Y(n_9361)
);

INVx2_ASAP7_75t_L g9362 ( 
.A(n_8865),
.Y(n_9362)
);

AND2x2_ASAP7_75t_L g9363 ( 
.A(n_8827),
.B(n_144),
.Y(n_9363)
);

NAND2xp5_ASAP7_75t_L g9364 ( 
.A(n_9043),
.B(n_23),
.Y(n_9364)
);

BUFx3_ASAP7_75t_L g9365 ( 
.A(n_8802),
.Y(n_9365)
);

INVx2_ASAP7_75t_L g9366 ( 
.A(n_8870),
.Y(n_9366)
);

NAND2xp5_ASAP7_75t_SL g9367 ( 
.A(n_8758),
.B(n_144),
.Y(n_9367)
);

NAND2xp5_ASAP7_75t_L g9368 ( 
.A(n_9043),
.B(n_23),
.Y(n_9368)
);

BUFx2_ASAP7_75t_L g9369 ( 
.A(n_9014),
.Y(n_9369)
);

INVx1_ASAP7_75t_L g9370 ( 
.A(n_8874),
.Y(n_9370)
);

AND2x2_ASAP7_75t_L g9371 ( 
.A(n_8850),
.B(n_145),
.Y(n_9371)
);

INVx1_ASAP7_75t_L g9372 ( 
.A(n_8875),
.Y(n_9372)
);

NAND2xp5_ASAP7_75t_L g9373 ( 
.A(n_9043),
.B(n_23),
.Y(n_9373)
);

NAND2xp5_ASAP7_75t_L g9374 ( 
.A(n_8883),
.B(n_24),
.Y(n_9374)
);

OR2x2_ASAP7_75t_L g9375 ( 
.A(n_8891),
.B(n_24),
.Y(n_9375)
);

HB1xp67_ASAP7_75t_L g9376 ( 
.A(n_8895),
.Y(n_9376)
);

INVx2_ASAP7_75t_L g9377 ( 
.A(n_8881),
.Y(n_9377)
);

AND2x2_ASAP7_75t_SL g9378 ( 
.A(n_9038),
.B(n_24),
.Y(n_9378)
);

INVx1_ASAP7_75t_L g9379 ( 
.A(n_8896),
.Y(n_9379)
);

INVx1_ASAP7_75t_L g9380 ( 
.A(n_8897),
.Y(n_9380)
);

NAND2xp5_ASAP7_75t_L g9381 ( 
.A(n_8909),
.B(n_25),
.Y(n_9381)
);

INVx1_ASAP7_75t_L g9382 ( 
.A(n_8911),
.Y(n_9382)
);

NAND2xp5_ASAP7_75t_L g9383 ( 
.A(n_8912),
.B(n_25),
.Y(n_9383)
);

NAND2xp5_ASAP7_75t_L g9384 ( 
.A(n_8927),
.B(n_26),
.Y(n_9384)
);

OAI21xp5_ASAP7_75t_L g9385 ( 
.A1(n_9066),
.A2(n_26),
.B(n_27),
.Y(n_9385)
);

OAI21xp5_ASAP7_75t_L g9386 ( 
.A1(n_8813),
.A2(n_26),
.B(n_27),
.Y(n_9386)
);

HB1xp67_ASAP7_75t_L g9387 ( 
.A(n_8931),
.Y(n_9387)
);

INVx1_ASAP7_75t_L g9388 ( 
.A(n_8934),
.Y(n_9388)
);

INVx2_ASAP7_75t_L g9389 ( 
.A(n_8902),
.Y(n_9389)
);

INVx3_ASAP7_75t_L g9390 ( 
.A(n_8914),
.Y(n_9390)
);

INVx2_ASAP7_75t_SL g9391 ( 
.A(n_8825),
.Y(n_9391)
);

INVx2_ASAP7_75t_L g9392 ( 
.A(n_8920),
.Y(n_9392)
);

INVx1_ASAP7_75t_L g9393 ( 
.A(n_8941),
.Y(n_9393)
);

BUFx3_ASAP7_75t_L g9394 ( 
.A(n_8832),
.Y(n_9394)
);

AND2x2_ASAP7_75t_SL g9395 ( 
.A(n_9201),
.B(n_27),
.Y(n_9395)
);

AND2x2_ASAP7_75t_L g9396 ( 
.A(n_9079),
.B(n_145),
.Y(n_9396)
);

AND2x2_ASAP7_75t_L g9397 ( 
.A(n_9119),
.B(n_8978),
.Y(n_9397)
);

OR2x2_ASAP7_75t_L g9398 ( 
.A(n_8947),
.B(n_28),
.Y(n_9398)
);

BUFx6f_ASAP7_75t_L g9399 ( 
.A(n_8833),
.Y(n_9399)
);

NAND2xp5_ASAP7_75t_L g9400 ( 
.A(n_8952),
.B(n_28),
.Y(n_9400)
);

OAI21xp5_ASAP7_75t_L g9401 ( 
.A1(n_8819),
.A2(n_29),
.B(n_30),
.Y(n_9401)
);

CKINVDCx5p33_ASAP7_75t_R g9402 ( 
.A(n_8778),
.Y(n_9402)
);

AND2x2_ASAP7_75t_L g9403 ( 
.A(n_9022),
.B(n_146),
.Y(n_9403)
);

AND2x2_ASAP7_75t_SL g9404 ( 
.A(n_8784),
.B(n_29),
.Y(n_9404)
);

AND2x2_ASAP7_75t_L g9405 ( 
.A(n_9067),
.B(n_147),
.Y(n_9405)
);

NAND2x1p5_ASAP7_75t_L g9406 ( 
.A(n_8837),
.B(n_147),
.Y(n_9406)
);

INVx2_ASAP7_75t_SL g9407 ( 
.A(n_9136),
.Y(n_9407)
);

AND2x2_ASAP7_75t_SL g9408 ( 
.A(n_8910),
.B(n_29),
.Y(n_9408)
);

INVx2_ASAP7_75t_L g9409 ( 
.A(n_8922),
.Y(n_9409)
);

INVx8_ASAP7_75t_L g9410 ( 
.A(n_8867),
.Y(n_9410)
);

BUFx6f_ASAP7_75t_L g9411 ( 
.A(n_9102),
.Y(n_9411)
);

INVx2_ASAP7_75t_L g9412 ( 
.A(n_8937),
.Y(n_9412)
);

AND2x2_ASAP7_75t_L g9413 ( 
.A(n_9144),
.B(n_148),
.Y(n_9413)
);

BUFx3_ASAP7_75t_L g9414 ( 
.A(n_8721),
.Y(n_9414)
);

NOR2xp67_ASAP7_75t_L g9415 ( 
.A(n_9183),
.B(n_9132),
.Y(n_9415)
);

HB1xp67_ASAP7_75t_L g9416 ( 
.A(n_8956),
.Y(n_9416)
);

OAI21xp5_ASAP7_75t_L g9417 ( 
.A1(n_8839),
.A2(n_30),
.B(n_31),
.Y(n_9417)
);

AND2x2_ASAP7_75t_L g9418 ( 
.A(n_9025),
.B(n_148),
.Y(n_9418)
);

NAND2xp5_ASAP7_75t_L g9419 ( 
.A(n_8960),
.B(n_30),
.Y(n_9419)
);

AND2x6_ASAP7_75t_L g9420 ( 
.A(n_8962),
.B(n_31),
.Y(n_9420)
);

NAND2xp5_ASAP7_75t_L g9421 ( 
.A(n_8964),
.B(n_32),
.Y(n_9421)
);

NAND2xp5_ASAP7_75t_SL g9422 ( 
.A(n_9172),
.B(n_149),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_8973),
.Y(n_9423)
);

INVx1_ASAP7_75t_L g9424 ( 
.A(n_8980),
.Y(n_9424)
);

BUFx6f_ASAP7_75t_L g9425 ( 
.A(n_9032),
.Y(n_9425)
);

BUFx3_ASAP7_75t_L g9426 ( 
.A(n_8856),
.Y(n_9426)
);

INVx1_ASAP7_75t_L g9427 ( 
.A(n_8990),
.Y(n_9427)
);

BUFx6f_ASAP7_75t_L g9428 ( 
.A(n_9221),
.Y(n_9428)
);

NAND2xp5_ASAP7_75t_L g9429 ( 
.A(n_8838),
.B(n_32),
.Y(n_9429)
);

INVxp67_ASAP7_75t_L g9430 ( 
.A(n_9154),
.Y(n_9430)
);

NOR2xp33_ASAP7_75t_L g9431 ( 
.A(n_8741),
.B(n_149),
.Y(n_9431)
);

INVx1_ASAP7_75t_L g9432 ( 
.A(n_9018),
.Y(n_9432)
);

INVx2_ASAP7_75t_L g9433 ( 
.A(n_8953),
.Y(n_9433)
);

HB1xp67_ASAP7_75t_L g9434 ( 
.A(n_9019),
.Y(n_9434)
);

INVx2_ASAP7_75t_L g9435 ( 
.A(n_8961),
.Y(n_9435)
);

INVx1_ASAP7_75t_L g9436 ( 
.A(n_9047),
.Y(n_9436)
);

INVxp67_ASAP7_75t_SL g9437 ( 
.A(n_8967),
.Y(n_9437)
);

INVx1_ASAP7_75t_L g9438 ( 
.A(n_9057),
.Y(n_9438)
);

BUFx3_ASAP7_75t_L g9439 ( 
.A(n_9125),
.Y(n_9439)
);

AND2x2_ASAP7_75t_L g9440 ( 
.A(n_8798),
.B(n_150),
.Y(n_9440)
);

AND2x4_ASAP7_75t_L g9441 ( 
.A(n_9120),
.B(n_150),
.Y(n_9441)
);

INVx2_ASAP7_75t_L g9442 ( 
.A(n_8988),
.Y(n_9442)
);

OR2x2_ASAP7_75t_L g9443 ( 
.A(n_9062),
.B(n_32),
.Y(n_9443)
);

NOR2xp33_ASAP7_75t_L g9444 ( 
.A(n_8726),
.B(n_151),
.Y(n_9444)
);

INVxp67_ASAP7_75t_SL g9445 ( 
.A(n_8722),
.Y(n_9445)
);

AND2x2_ASAP7_75t_SL g9446 ( 
.A(n_8948),
.B(n_33),
.Y(n_9446)
);

INVx2_ASAP7_75t_SL g9447 ( 
.A(n_9138),
.Y(n_9447)
);

INVx1_ASAP7_75t_L g9448 ( 
.A(n_9063),
.Y(n_9448)
);

AND2x2_ASAP7_75t_L g9449 ( 
.A(n_8733),
.B(n_151),
.Y(n_9449)
);

HB1xp67_ASAP7_75t_L g9450 ( 
.A(n_9133),
.Y(n_9450)
);

BUFx6f_ASAP7_75t_L g9451 ( 
.A(n_9204),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_9069),
.Y(n_9452)
);

NAND2xp5_ASAP7_75t_L g9453 ( 
.A(n_8747),
.B(n_8744),
.Y(n_9453)
);

NOR2xp33_ASAP7_75t_L g9454 ( 
.A(n_9028),
.B(n_152),
.Y(n_9454)
);

AND2x2_ASAP7_75t_L g9455 ( 
.A(n_8851),
.B(n_152),
.Y(n_9455)
);

NAND2xp5_ASAP7_75t_L g9456 ( 
.A(n_9134),
.B(n_33),
.Y(n_9456)
);

INVx1_ASAP7_75t_L g9457 ( 
.A(n_9078),
.Y(n_9457)
);

AND2x2_ASAP7_75t_L g9458 ( 
.A(n_8951),
.B(n_153),
.Y(n_9458)
);

INVx2_ASAP7_75t_L g9459 ( 
.A(n_8997),
.Y(n_9459)
);

OAI21xp5_ASAP7_75t_L g9460 ( 
.A1(n_8840),
.A2(n_8843),
.B(n_9024),
.Y(n_9460)
);

NOR2xp33_ASAP7_75t_L g9461 ( 
.A(n_8918),
.B(n_153),
.Y(n_9461)
);

NOR2xp33_ASAP7_75t_L g9462 ( 
.A(n_8779),
.B(n_8879),
.Y(n_9462)
);

HB1xp67_ASAP7_75t_L g9463 ( 
.A(n_9082),
.Y(n_9463)
);

AND2x2_ASAP7_75t_L g9464 ( 
.A(n_8951),
.B(n_154),
.Y(n_9464)
);

INVxp67_ASAP7_75t_SL g9465 ( 
.A(n_8751),
.Y(n_9465)
);

AND2x2_ASAP7_75t_L g9466 ( 
.A(n_8981),
.B(n_154),
.Y(n_9466)
);

HB1xp67_ASAP7_75t_L g9467 ( 
.A(n_9085),
.Y(n_9467)
);

NAND2xp5_ASAP7_75t_L g9468 ( 
.A(n_8749),
.B(n_8750),
.Y(n_9468)
);

NOR2xp33_ASAP7_75t_L g9469 ( 
.A(n_8907),
.B(n_155),
.Y(n_9469)
);

NAND2xp5_ASAP7_75t_L g9470 ( 
.A(n_8766),
.B(n_34),
.Y(n_9470)
);

INVx1_ASAP7_75t_SL g9471 ( 
.A(n_8977),
.Y(n_9471)
);

INVx2_ASAP7_75t_L g9472 ( 
.A(n_9013),
.Y(n_9472)
);

BUFx10_ASAP7_75t_L g9473 ( 
.A(n_8901),
.Y(n_9473)
);

NAND2xp5_ASAP7_75t_L g9474 ( 
.A(n_8773),
.B(n_34),
.Y(n_9474)
);

AND2x2_ASAP7_75t_L g9475 ( 
.A(n_9005),
.B(n_155),
.Y(n_9475)
);

AND2x2_ASAP7_75t_L g9476 ( 
.A(n_8975),
.B(n_156),
.Y(n_9476)
);

AND2x2_ASAP7_75t_L g9477 ( 
.A(n_9086),
.B(n_8796),
.Y(n_9477)
);

INVx1_ASAP7_75t_L g9478 ( 
.A(n_9091),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_9093),
.Y(n_9479)
);

OR2x2_ASAP7_75t_L g9480 ( 
.A(n_9100),
.B(n_9108),
.Y(n_9480)
);

INVx2_ASAP7_75t_SL g9481 ( 
.A(n_9218),
.Y(n_9481)
);

HB1xp67_ASAP7_75t_L g9482 ( 
.A(n_9112),
.Y(n_9482)
);

NOR2xp33_ASAP7_75t_L g9483 ( 
.A(n_8877),
.B(n_156),
.Y(n_9483)
);

AND2x2_ASAP7_75t_L g9484 ( 
.A(n_9053),
.B(n_157),
.Y(n_9484)
);

INVx2_ASAP7_75t_L g9485 ( 
.A(n_9015),
.Y(n_9485)
);

AND2x2_ASAP7_75t_L g9486 ( 
.A(n_8869),
.B(n_157),
.Y(n_9486)
);

INVx1_ASAP7_75t_L g9487 ( 
.A(n_9113),
.Y(n_9487)
);

HB1xp67_ASAP7_75t_L g9488 ( 
.A(n_9129),
.Y(n_9488)
);

OAI21x1_ASAP7_75t_L g9489 ( 
.A1(n_8725),
.A2(n_159),
.B(n_158),
.Y(n_9489)
);

INVx1_ASAP7_75t_L g9490 ( 
.A(n_9114),
.Y(n_9490)
);

INVx1_ASAP7_75t_L g9491 ( 
.A(n_9029),
.Y(n_9491)
);

INVxp67_ASAP7_75t_SL g9492 ( 
.A(n_8788),
.Y(n_9492)
);

INVx3_ASAP7_75t_L g9493 ( 
.A(n_8858),
.Y(n_9493)
);

INVx1_ASAP7_75t_L g9494 ( 
.A(n_9137),
.Y(n_9494)
);

OR2x2_ASAP7_75t_SL g9495 ( 
.A(n_9233),
.B(n_34),
.Y(n_9495)
);

NAND2x1p5_ASAP7_75t_L g9496 ( 
.A(n_9151),
.B(n_158),
.Y(n_9496)
);

BUFx2_ASAP7_75t_L g9497 ( 
.A(n_9171),
.Y(n_9497)
);

AND2x4_ASAP7_75t_L g9498 ( 
.A(n_9161),
.B(n_159),
.Y(n_9498)
);

NAND2xp5_ASAP7_75t_L g9499 ( 
.A(n_8945),
.B(n_35),
.Y(n_9499)
);

INVx1_ASAP7_75t_L g9500 ( 
.A(n_9141),
.Y(n_9500)
);

INVx2_ASAP7_75t_L g9501 ( 
.A(n_9017),
.Y(n_9501)
);

NAND2xp5_ASAP7_75t_L g9502 ( 
.A(n_9212),
.B(n_35),
.Y(n_9502)
);

NAND2xp5_ASAP7_75t_L g9503 ( 
.A(n_9219),
.B(n_35),
.Y(n_9503)
);

INVx1_ASAP7_75t_L g9504 ( 
.A(n_9178),
.Y(n_9504)
);

INVx1_ASAP7_75t_SL g9505 ( 
.A(n_8762),
.Y(n_9505)
);

INVx1_ASAP7_75t_L g9506 ( 
.A(n_9180),
.Y(n_9506)
);

AND2x2_ASAP7_75t_SL g9507 ( 
.A(n_9207),
.B(n_36),
.Y(n_9507)
);

AND2x2_ASAP7_75t_L g9508 ( 
.A(n_9208),
.B(n_160),
.Y(n_9508)
);

NAND2xp5_ASAP7_75t_L g9509 ( 
.A(n_8809),
.B(n_36),
.Y(n_9509)
);

OAI21xp5_ASAP7_75t_L g9510 ( 
.A1(n_8959),
.A2(n_36),
.B(n_37),
.Y(n_9510)
);

AND2x2_ASAP7_75t_L g9511 ( 
.A(n_8892),
.B(n_160),
.Y(n_9511)
);

HB1xp67_ASAP7_75t_L g9512 ( 
.A(n_9194),
.Y(n_9512)
);

AND2x2_ASAP7_75t_L g9513 ( 
.A(n_8916),
.B(n_161),
.Y(n_9513)
);

AND2x2_ASAP7_75t_L g9514 ( 
.A(n_8753),
.B(n_161),
.Y(n_9514)
);

INVx1_ASAP7_75t_L g9515 ( 
.A(n_9192),
.Y(n_9515)
);

INVx8_ASAP7_75t_L g9516 ( 
.A(n_9072),
.Y(n_9516)
);

AND2x2_ASAP7_75t_L g9517 ( 
.A(n_8760),
.B(n_162),
.Y(n_9517)
);

INVx1_ASAP7_75t_L g9518 ( 
.A(n_9199),
.Y(n_9518)
);

AND2x6_ASAP7_75t_L g9519 ( 
.A(n_9215),
.B(n_37),
.Y(n_9519)
);

AND2x2_ASAP7_75t_L g9520 ( 
.A(n_8942),
.B(n_162),
.Y(n_9520)
);

BUFx3_ASAP7_75t_L g9521 ( 
.A(n_8938),
.Y(n_9521)
);

NAND2xp5_ASAP7_75t_L g9522 ( 
.A(n_8789),
.B(n_37),
.Y(n_9522)
);

AND2x2_ASAP7_75t_L g9523 ( 
.A(n_9045),
.B(n_163),
.Y(n_9523)
);

INVx4_ASAP7_75t_L g9524 ( 
.A(n_8823),
.Y(n_9524)
);

AND2x2_ASAP7_75t_L g9525 ( 
.A(n_8872),
.B(n_163),
.Y(n_9525)
);

AND2x2_ASAP7_75t_L g9526 ( 
.A(n_8876),
.B(n_164),
.Y(n_9526)
);

BUFx6f_ASAP7_75t_L g9527 ( 
.A(n_8950),
.Y(n_9527)
);

AND2x2_ASAP7_75t_SL g9528 ( 
.A(n_8954),
.B(n_8834),
.Y(n_9528)
);

NAND2xp5_ASAP7_75t_L g9529 ( 
.A(n_8755),
.B(n_38),
.Y(n_9529)
);

INVx1_ASAP7_75t_L g9530 ( 
.A(n_9039),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_9049),
.Y(n_9531)
);

NAND2xp5_ASAP7_75t_L g9532 ( 
.A(n_8880),
.B(n_8737),
.Y(n_9532)
);

AND2x2_ASAP7_75t_L g9533 ( 
.A(n_8785),
.B(n_165),
.Y(n_9533)
);

OAI21xp5_ASAP7_75t_L g9534 ( 
.A1(n_8728),
.A2(n_38),
.B(n_39),
.Y(n_9534)
);

INVx1_ASAP7_75t_L g9535 ( 
.A(n_9051),
.Y(n_9535)
);

BUFx3_ASAP7_75t_L g9536 ( 
.A(n_9227),
.Y(n_9536)
);

INVx2_ASAP7_75t_L g9537 ( 
.A(n_9059),
.Y(n_9537)
);

AND2x2_ASAP7_75t_L g9538 ( 
.A(n_9147),
.B(n_165),
.Y(n_9538)
);

INVx1_ASAP7_75t_L g9539 ( 
.A(n_9064),
.Y(n_9539)
);

INVx1_ASAP7_75t_L g9540 ( 
.A(n_9068),
.Y(n_9540)
);

AND2x2_ASAP7_75t_L g9541 ( 
.A(n_8863),
.B(n_167),
.Y(n_9541)
);

BUFx4f_ASAP7_75t_L g9542 ( 
.A(n_9072),
.Y(n_9542)
);

INVx2_ASAP7_75t_L g9543 ( 
.A(n_9073),
.Y(n_9543)
);

INVx3_ASAP7_75t_L g9544 ( 
.A(n_9231),
.Y(n_9544)
);

INVx2_ASAP7_75t_SL g9545 ( 
.A(n_9164),
.Y(n_9545)
);

NAND2xp5_ASAP7_75t_L g9546 ( 
.A(n_9146),
.B(n_38),
.Y(n_9546)
);

INVx2_ASAP7_75t_L g9547 ( 
.A(n_9076),
.Y(n_9547)
);

NAND2xp5_ASAP7_75t_L g9548 ( 
.A(n_8783),
.B(n_40),
.Y(n_9548)
);

INVx3_ASAP7_75t_L g9549 ( 
.A(n_9104),
.Y(n_9549)
);

AND2x2_ASAP7_75t_L g9550 ( 
.A(n_9099),
.B(n_167),
.Y(n_9550)
);

INVx1_ASAP7_75t_L g9551 ( 
.A(n_9077),
.Y(n_9551)
);

NAND2xp5_ASAP7_75t_L g9552 ( 
.A(n_8853),
.B(n_40),
.Y(n_9552)
);

AND2x2_ASAP7_75t_L g9553 ( 
.A(n_8790),
.B(n_168),
.Y(n_9553)
);

BUFx5_ASAP7_75t_L g9554 ( 
.A(n_9060),
.Y(n_9554)
);

NAND2xp5_ASAP7_75t_SL g9555 ( 
.A(n_8764),
.B(n_168),
.Y(n_9555)
);

INVx1_ASAP7_75t_L g9556 ( 
.A(n_9096),
.Y(n_9556)
);

INVx1_ASAP7_75t_L g9557 ( 
.A(n_9105),
.Y(n_9557)
);

BUFx3_ASAP7_75t_L g9558 ( 
.A(n_9217),
.Y(n_9558)
);

INVx2_ASAP7_75t_L g9559 ( 
.A(n_9135),
.Y(n_9559)
);

OAI21xp5_ASAP7_75t_L g9560 ( 
.A1(n_8987),
.A2(n_41),
.B(n_42),
.Y(n_9560)
);

AND2x2_ASAP7_75t_L g9561 ( 
.A(n_8794),
.B(n_169),
.Y(n_9561)
);

HB1xp67_ASAP7_75t_L g9562 ( 
.A(n_9234),
.Y(n_9562)
);

OAI21xp5_ASAP7_75t_L g9563 ( 
.A1(n_8797),
.A2(n_41),
.B(n_42),
.Y(n_9563)
);

INVx1_ASAP7_75t_L g9564 ( 
.A(n_9148),
.Y(n_9564)
);

INVx1_ASAP7_75t_L g9565 ( 
.A(n_9152),
.Y(n_9565)
);

NAND2xp5_ASAP7_75t_L g9566 ( 
.A(n_8888),
.B(n_41),
.Y(n_9566)
);

INVx2_ASAP7_75t_L g9567 ( 
.A(n_9153),
.Y(n_9567)
);

AND2x2_ASAP7_75t_SL g9568 ( 
.A(n_9236),
.B(n_43),
.Y(n_9568)
);

AND2x2_ASAP7_75t_L g9569 ( 
.A(n_8864),
.B(n_170),
.Y(n_9569)
);

INVx3_ASAP7_75t_L g9570 ( 
.A(n_9235),
.Y(n_9570)
);

AND2x2_ASAP7_75t_L g9571 ( 
.A(n_8854),
.B(n_171),
.Y(n_9571)
);

NAND2xp5_ASAP7_75t_L g9572 ( 
.A(n_9156),
.B(n_43),
.Y(n_9572)
);

BUFx3_ASAP7_75t_L g9573 ( 
.A(n_9220),
.Y(n_9573)
);

INVx2_ASAP7_75t_L g9574 ( 
.A(n_9166),
.Y(n_9574)
);

INVx2_ASAP7_75t_L g9575 ( 
.A(n_9177),
.Y(n_9575)
);

AND2x2_ASAP7_75t_L g9576 ( 
.A(n_9149),
.B(n_171),
.Y(n_9576)
);

INVx1_ASAP7_75t_L g9577 ( 
.A(n_9182),
.Y(n_9577)
);

AND2x2_ASAP7_75t_L g9578 ( 
.A(n_8745),
.B(n_172),
.Y(n_9578)
);

OAI21xp5_ASAP7_75t_L g9579 ( 
.A1(n_8780),
.A2(n_43),
.B(n_44),
.Y(n_9579)
);

AND2x2_ASAP7_75t_L g9580 ( 
.A(n_9040),
.B(n_173),
.Y(n_9580)
);

AND2x2_ASAP7_75t_L g9581 ( 
.A(n_9225),
.B(n_173),
.Y(n_9581)
);

NAND2xp5_ASAP7_75t_L g9582 ( 
.A(n_9123),
.B(n_44),
.Y(n_9582)
);

INVx2_ASAP7_75t_L g9583 ( 
.A(n_9200),
.Y(n_9583)
);

NOR2xp33_ASAP7_75t_L g9584 ( 
.A(n_8886),
.B(n_174),
.Y(n_9584)
);

INVx2_ASAP7_75t_L g9585 ( 
.A(n_9206),
.Y(n_9585)
);

INVx1_ASAP7_75t_L g9586 ( 
.A(n_9209),
.Y(n_9586)
);

AND2x4_ASAP7_75t_L g9587 ( 
.A(n_9232),
.B(n_174),
.Y(n_9587)
);

INVx4_ASAP7_75t_L g9588 ( 
.A(n_9021),
.Y(n_9588)
);

HB1xp67_ASAP7_75t_L g9589 ( 
.A(n_9210),
.Y(n_9589)
);

AND2x2_ASAP7_75t_L g9590 ( 
.A(n_8822),
.B(n_175),
.Y(n_9590)
);

NOR2xp33_ASAP7_75t_L g9591 ( 
.A(n_8782),
.B(n_175),
.Y(n_9591)
);

AND2x2_ASAP7_75t_L g9592 ( 
.A(n_8792),
.B(n_176),
.Y(n_9592)
);

INVx1_ASAP7_75t_L g9593 ( 
.A(n_9213),
.Y(n_9593)
);

NAND2xp5_ASAP7_75t_L g9594 ( 
.A(n_8768),
.B(n_44),
.Y(n_9594)
);

INVx2_ASAP7_75t_L g9595 ( 
.A(n_9214),
.Y(n_9595)
);

NOR2xp33_ASAP7_75t_L g9596 ( 
.A(n_8808),
.B(n_176),
.Y(n_9596)
);

AND2x2_ASAP7_75t_L g9597 ( 
.A(n_9041),
.B(n_177),
.Y(n_9597)
);

NAND2xp5_ASAP7_75t_L g9598 ( 
.A(n_9002),
.B(n_45),
.Y(n_9598)
);

INVx1_ASAP7_75t_L g9599 ( 
.A(n_9196),
.Y(n_9599)
);

NAND2xp5_ASAP7_75t_L g9600 ( 
.A(n_9004),
.B(n_8887),
.Y(n_9600)
);

AND2x4_ASAP7_75t_L g9601 ( 
.A(n_8800),
.B(n_177),
.Y(n_9601)
);

INVx4_ASAP7_75t_L g9602 ( 
.A(n_8806),
.Y(n_9602)
);

INVx2_ASAP7_75t_L g9603 ( 
.A(n_9203),
.Y(n_9603)
);

OAI21x1_ASAP7_75t_L g9604 ( 
.A1(n_9001),
.A2(n_179),
.B(n_178),
.Y(n_9604)
);

AND2x4_ASAP7_75t_SL g9605 ( 
.A(n_9074),
.B(n_9095),
.Y(n_9605)
);

INVx1_ASAP7_75t_L g9606 ( 
.A(n_9202),
.Y(n_9606)
);

NOR2xp33_ASAP7_75t_SL g9607 ( 
.A(n_9116),
.B(n_45),
.Y(n_9607)
);

CKINVDCx5p33_ASAP7_75t_R g9608 ( 
.A(n_9169),
.Y(n_9608)
);

INVx1_ASAP7_75t_L g9609 ( 
.A(n_9205),
.Y(n_9609)
);

AND2x2_ASAP7_75t_L g9610 ( 
.A(n_8847),
.B(n_179),
.Y(n_9610)
);

BUFx3_ASAP7_75t_L g9611 ( 
.A(n_9110),
.Y(n_9611)
);

AND2x2_ASAP7_75t_L g9612 ( 
.A(n_9188),
.B(n_180),
.Y(n_9612)
);

INVx1_ASAP7_75t_L g9613 ( 
.A(n_9229),
.Y(n_9613)
);

INVx2_ASAP7_75t_L g9614 ( 
.A(n_9111),
.Y(n_9614)
);

OR2x2_ASAP7_75t_L g9615 ( 
.A(n_8893),
.B(n_46),
.Y(n_9615)
);

INVx4_ASAP7_75t_L g9616 ( 
.A(n_8932),
.Y(n_9616)
);

AND2x2_ASAP7_75t_L g9617 ( 
.A(n_8898),
.B(n_180),
.Y(n_9617)
);

INVx2_ASAP7_75t_L g9618 ( 
.A(n_9179),
.Y(n_9618)
);

INVx2_ASAP7_75t_L g9619 ( 
.A(n_9186),
.Y(n_9619)
);

INVx3_ASAP7_75t_L g9620 ( 
.A(n_9007),
.Y(n_9620)
);

BUFx6f_ASAP7_75t_L g9621 ( 
.A(n_8774),
.Y(n_9621)
);

AND2x2_ASAP7_75t_SL g9622 ( 
.A(n_9222),
.B(n_46),
.Y(n_9622)
);

NAND2xp5_ASAP7_75t_L g9623 ( 
.A(n_8903),
.B(n_46),
.Y(n_9623)
);

NAND2xp5_ASAP7_75t_L g9624 ( 
.A(n_8905),
.B(n_8906),
.Y(n_9624)
);

HB1xp67_ASAP7_75t_L g9625 ( 
.A(n_8759),
.Y(n_9625)
);

HB1xp67_ASAP7_75t_L g9626 ( 
.A(n_8770),
.Y(n_9626)
);

AND2x2_ASAP7_75t_L g9627 ( 
.A(n_8921),
.B(n_181),
.Y(n_9627)
);

INVx1_ASAP7_75t_L g9628 ( 
.A(n_9216),
.Y(n_9628)
);

NAND2xp5_ASAP7_75t_SL g9629 ( 
.A(n_8739),
.B(n_181),
.Y(n_9629)
);

AND2x2_ASAP7_75t_L g9630 ( 
.A(n_8925),
.B(n_182),
.Y(n_9630)
);

AND2x2_ASAP7_75t_L g9631 ( 
.A(n_8926),
.B(n_182),
.Y(n_9631)
);

INVx2_ASAP7_75t_SL g9632 ( 
.A(n_8946),
.Y(n_9632)
);

OR2x2_ASAP7_75t_L g9633 ( 
.A(n_8929),
.B(n_47),
.Y(n_9633)
);

INVx1_ASAP7_75t_L g9634 ( 
.A(n_9228),
.Y(n_9634)
);

NAND2xp5_ASAP7_75t_L g9635 ( 
.A(n_8933),
.B(n_47),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_9223),
.Y(n_9636)
);

NAND2xp5_ASAP7_75t_L g9637 ( 
.A(n_8935),
.B(n_47),
.Y(n_9637)
);

NAND2xp5_ASAP7_75t_L g9638 ( 
.A(n_8944),
.B(n_8971),
.Y(n_9638)
);

HB1xp67_ASAP7_75t_L g9639 ( 
.A(n_9191),
.Y(n_9639)
);

INVx2_ASAP7_75t_L g9640 ( 
.A(n_9128),
.Y(n_9640)
);

INVx1_ASAP7_75t_L g9641 ( 
.A(n_9195),
.Y(n_9641)
);

INVx1_ASAP7_75t_L g9642 ( 
.A(n_8982),
.Y(n_9642)
);

NOR2xp33_ASAP7_75t_L g9643 ( 
.A(n_8793),
.B(n_183),
.Y(n_9643)
);

INVx1_ASAP7_75t_L g9644 ( 
.A(n_8986),
.Y(n_9644)
);

AND2x2_ASAP7_75t_L g9645 ( 
.A(n_8972),
.B(n_183),
.Y(n_9645)
);

AND2x6_ASAP7_75t_L g9646 ( 
.A(n_9198),
.B(n_48),
.Y(n_9646)
);

INVx1_ASAP7_75t_L g9647 ( 
.A(n_8989),
.Y(n_9647)
);

NAND2xp5_ASAP7_75t_L g9648 ( 
.A(n_9016),
.B(n_48),
.Y(n_9648)
);

NAND2xp5_ASAP7_75t_L g9649 ( 
.A(n_9176),
.B(n_9142),
.Y(n_9649)
);

INVx2_ASAP7_75t_L g9650 ( 
.A(n_9083),
.Y(n_9650)
);

AND2x2_ASAP7_75t_L g9651 ( 
.A(n_9103),
.B(n_184),
.Y(n_9651)
);

INVx1_ASAP7_75t_L g9652 ( 
.A(n_9224),
.Y(n_9652)
);

INVx2_ASAP7_75t_L g9653 ( 
.A(n_9127),
.Y(n_9653)
);

NAND2xp5_ASAP7_75t_L g9654 ( 
.A(n_8958),
.B(n_48),
.Y(n_9654)
);

NAND2xp5_ASAP7_75t_L g9655 ( 
.A(n_9020),
.B(n_49),
.Y(n_9655)
);

INVx6_ASAP7_75t_L g9656 ( 
.A(n_8804),
.Y(n_9656)
);

INVx1_ASAP7_75t_L g9657 ( 
.A(n_8991),
.Y(n_9657)
);

BUFx6f_ASAP7_75t_L g9658 ( 
.A(n_9117),
.Y(n_9658)
);

INVx3_ASAP7_75t_L g9659 ( 
.A(n_9150),
.Y(n_9659)
);

INVx3_ASAP7_75t_L g9660 ( 
.A(n_9170),
.Y(n_9660)
);

INVx2_ASAP7_75t_L g9661 ( 
.A(n_9139),
.Y(n_9661)
);

AND2x2_ASAP7_75t_L g9662 ( 
.A(n_9162),
.B(n_9184),
.Y(n_9662)
);

AND2x4_ASAP7_75t_SL g9663 ( 
.A(n_9181),
.B(n_184),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_9189),
.Y(n_9664)
);

AND2x2_ASAP7_75t_L g9665 ( 
.A(n_9042),
.B(n_185),
.Y(n_9665)
);

INVx2_ASAP7_75t_L g9666 ( 
.A(n_9140),
.Y(n_9666)
);

HB1xp67_ASAP7_75t_L g9667 ( 
.A(n_9055),
.Y(n_9667)
);

NOR2xp33_ASAP7_75t_L g9668 ( 
.A(n_8801),
.B(n_185),
.Y(n_9668)
);

NAND2xp5_ASAP7_75t_SL g9669 ( 
.A(n_9061),
.B(n_186),
.Y(n_9669)
);

INVx1_ASAP7_75t_L g9670 ( 
.A(n_8841),
.Y(n_9670)
);

INVx1_ASAP7_75t_L g9671 ( 
.A(n_9173),
.Y(n_9671)
);

INVx3_ASAP7_75t_L g9672 ( 
.A(n_9101),
.Y(n_9672)
);

NOR2xp33_ASAP7_75t_L g9673 ( 
.A(n_9106),
.B(n_186),
.Y(n_9673)
);

INVx1_ASAP7_75t_SL g9674 ( 
.A(n_8814),
.Y(n_9674)
);

AND2x2_ASAP7_75t_L g9675 ( 
.A(n_9046),
.B(n_187),
.Y(n_9675)
);

AND2x4_ASAP7_75t_L g9676 ( 
.A(n_8815),
.B(n_187),
.Y(n_9676)
);

AND2x2_ASAP7_75t_L g9677 ( 
.A(n_9155),
.B(n_188),
.Y(n_9677)
);

AND2x2_ASAP7_75t_L g9678 ( 
.A(n_8811),
.B(n_8908),
.Y(n_9678)
);

HB1xp67_ASAP7_75t_L g9679 ( 
.A(n_8807),
.Y(n_9679)
);

HB1xp67_ASAP7_75t_L g9680 ( 
.A(n_8859),
.Y(n_9680)
);

OAI21xp5_ASAP7_75t_L g9681 ( 
.A1(n_9031),
.A2(n_50),
.B(n_51),
.Y(n_9681)
);

BUFx3_ASAP7_75t_L g9682 ( 
.A(n_9092),
.Y(n_9682)
);

INVx3_ASAP7_75t_L g9683 ( 
.A(n_9097),
.Y(n_9683)
);

BUFx8_ASAP7_75t_L g9684 ( 
.A(n_8817),
.Y(n_9684)
);

INVx2_ASAP7_75t_L g9685 ( 
.A(n_9157),
.Y(n_9685)
);

NOR2xp33_ASAP7_75t_L g9686 ( 
.A(n_8992),
.B(n_189),
.Y(n_9686)
);

HB1xp67_ASAP7_75t_L g9687 ( 
.A(n_9158),
.Y(n_9687)
);

NAND2xp5_ASAP7_75t_L g9688 ( 
.A(n_9033),
.B(n_50),
.Y(n_9688)
);

BUFx3_ASAP7_75t_L g9689 ( 
.A(n_9087),
.Y(n_9689)
);

INVx1_ASAP7_75t_L g9690 ( 
.A(n_9190),
.Y(n_9690)
);

INVx3_ASAP7_75t_L g9691 ( 
.A(n_8974),
.Y(n_9691)
);

NOR2xp33_ASAP7_75t_L g9692 ( 
.A(n_9009),
.B(n_189),
.Y(n_9692)
);

OAI21xp5_ASAP7_75t_L g9693 ( 
.A1(n_9010),
.A2(n_50),
.B(n_51),
.Y(n_9693)
);

INVx3_ASAP7_75t_L g9694 ( 
.A(n_8994),
.Y(n_9694)
);

INVx3_ASAP7_75t_L g9695 ( 
.A(n_8999),
.Y(n_9695)
);

HB1xp67_ASAP7_75t_L g9696 ( 
.A(n_9167),
.Y(n_9696)
);

INVx2_ASAP7_75t_L g9697 ( 
.A(n_9185),
.Y(n_9697)
);

BUFx3_ASAP7_75t_L g9698 ( 
.A(n_9006),
.Y(n_9698)
);

NAND2xp5_ASAP7_75t_L g9699 ( 
.A(n_9211),
.B(n_51),
.Y(n_9699)
);

AND2x2_ASAP7_75t_L g9700 ( 
.A(n_8878),
.B(n_190),
.Y(n_9700)
);

AND2x2_ASAP7_75t_L g9701 ( 
.A(n_9160),
.B(n_190),
.Y(n_9701)
);

INVx2_ASAP7_75t_L g9702 ( 
.A(n_9187),
.Y(n_9702)
);

AND2x2_ASAP7_75t_L g9703 ( 
.A(n_9115),
.B(n_191),
.Y(n_9703)
);

HB1xp67_ASAP7_75t_L g9704 ( 
.A(n_9124),
.Y(n_9704)
);

NAND2xp5_ASAP7_75t_L g9705 ( 
.A(n_8955),
.B(n_52),
.Y(n_9705)
);

AND2x2_ASAP7_75t_L g9706 ( 
.A(n_8884),
.B(n_191),
.Y(n_9706)
);

INVx4_ASAP7_75t_L g9707 ( 
.A(n_8818),
.Y(n_9707)
);

NOR2xp33_ASAP7_75t_L g9708 ( 
.A(n_8900),
.B(n_193),
.Y(n_9708)
);

AND2x2_ASAP7_75t_L g9709 ( 
.A(n_8913),
.B(n_193),
.Y(n_9709)
);

INVxp67_ASAP7_75t_SL g9710 ( 
.A(n_9058),
.Y(n_9710)
);

NAND2xp5_ASAP7_75t_L g9711 ( 
.A(n_8970),
.B(n_52),
.Y(n_9711)
);

HB1xp67_ASAP7_75t_L g9712 ( 
.A(n_8949),
.Y(n_9712)
);

INVx1_ASAP7_75t_L g9713 ( 
.A(n_9052),
.Y(n_9713)
);

INVx2_ASAP7_75t_L g9714 ( 
.A(n_8966),
.Y(n_9714)
);

AND2x2_ASAP7_75t_L g9715 ( 
.A(n_8979),
.B(n_194),
.Y(n_9715)
);

NOR2xp33_ASAP7_75t_L g9716 ( 
.A(n_8983),
.B(n_194),
.Y(n_9716)
);

INVx1_ASAP7_75t_L g9717 ( 
.A(n_9071),
.Y(n_9717)
);

INVxp33_ASAP7_75t_L g9718 ( 
.A(n_8821),
.Y(n_9718)
);

AND2x2_ASAP7_75t_L g9719 ( 
.A(n_8939),
.B(n_195),
.Y(n_9719)
);

AND2x2_ASAP7_75t_L g9720 ( 
.A(n_9168),
.B(n_196),
.Y(n_9720)
);

BUFx3_ASAP7_75t_L g9721 ( 
.A(n_9121),
.Y(n_9721)
);

AND2x2_ASAP7_75t_L g9722 ( 
.A(n_9174),
.B(n_197),
.Y(n_9722)
);

INVx1_ASAP7_75t_L g9723 ( 
.A(n_8976),
.Y(n_9723)
);

INVxp67_ASAP7_75t_SL g9724 ( 
.A(n_8984),
.Y(n_9724)
);

NAND2xp5_ASAP7_75t_L g9725 ( 
.A(n_9027),
.B(n_52),
.Y(n_9725)
);

NOR2xp33_ASAP7_75t_L g9726 ( 
.A(n_9003),
.B(n_197),
.Y(n_9726)
);

INVx2_ASAP7_75t_L g9727 ( 
.A(n_9012),
.Y(n_9727)
);

INVx4_ASAP7_75t_L g9728 ( 
.A(n_8866),
.Y(n_9728)
);

AND2x2_ASAP7_75t_L g9729 ( 
.A(n_9011),
.B(n_198),
.Y(n_9729)
);

BUFx3_ASAP7_75t_L g9730 ( 
.A(n_9159),
.Y(n_9730)
);

INVx2_ASAP7_75t_L g9731 ( 
.A(n_9026),
.Y(n_9731)
);

BUFx2_ASAP7_75t_L g9732 ( 
.A(n_9070),
.Y(n_9732)
);

BUFx3_ASAP7_75t_L g9733 ( 
.A(n_8915),
.Y(n_9733)
);

NAND2xp5_ASAP7_75t_L g9734 ( 
.A(n_8904),
.B(n_53),
.Y(n_9734)
);

NAND2xp5_ASAP7_75t_L g9735 ( 
.A(n_8924),
.B(n_53),
.Y(n_9735)
);

NAND2xp5_ASAP7_75t_L g9736 ( 
.A(n_9035),
.B(n_54),
.Y(n_9736)
);

AND2x2_ASAP7_75t_L g9737 ( 
.A(n_9036),
.B(n_198),
.Y(n_9737)
);

BUFx3_ASAP7_75t_L g9738 ( 
.A(n_8917),
.Y(n_9738)
);

INVxp67_ASAP7_75t_SL g9739 ( 
.A(n_9084),
.Y(n_9739)
);

HB1xp67_ASAP7_75t_L g9740 ( 
.A(n_9088),
.Y(n_9740)
);

AND2x4_ASAP7_75t_L g9741 ( 
.A(n_9089),
.B(n_199),
.Y(n_9741)
);

AND2x2_ASAP7_75t_L g9742 ( 
.A(n_9130),
.B(n_199),
.Y(n_9742)
);

INVx2_ASAP7_75t_SL g9743 ( 
.A(n_9094),
.Y(n_9743)
);

AND2x4_ASAP7_75t_L g9744 ( 
.A(n_8849),
.B(n_200),
.Y(n_9744)
);

AND2x2_ASAP7_75t_L g9745 ( 
.A(n_9044),
.B(n_200),
.Y(n_9745)
);

INVx2_ASAP7_75t_L g9746 ( 
.A(n_8882),
.Y(n_9746)
);

INVx1_ASAP7_75t_SL g9747 ( 
.A(n_9098),
.Y(n_9747)
);

AND2x2_ASAP7_75t_L g9748 ( 
.A(n_8732),
.B(n_201),
.Y(n_9748)
);

BUFx4f_ASAP7_75t_L g9749 ( 
.A(n_8730),
.Y(n_9749)
);

NAND2xp5_ASAP7_75t_L g9750 ( 
.A(n_8729),
.B(n_54),
.Y(n_9750)
);

NAND2xp5_ASAP7_75t_L g9751 ( 
.A(n_8729),
.B(n_54),
.Y(n_9751)
);

NAND2xp5_ASAP7_75t_SL g9752 ( 
.A(n_9034),
.B(n_201),
.Y(n_9752)
);

AND2x2_ASAP7_75t_L g9753 ( 
.A(n_8732),
.B(n_202),
.Y(n_9753)
);

NAND2xp5_ASAP7_75t_L g9754 ( 
.A(n_8729),
.B(n_55),
.Y(n_9754)
);

INVx2_ASAP7_75t_L g9755 ( 
.A(n_8723),
.Y(n_9755)
);

INVx1_ASAP7_75t_SL g9756 ( 
.A(n_9098),
.Y(n_9756)
);

AND2x2_ASAP7_75t_L g9757 ( 
.A(n_8732),
.B(n_203),
.Y(n_9757)
);

INVx1_ASAP7_75t_L g9758 ( 
.A(n_8889),
.Y(n_9758)
);

INVx1_ASAP7_75t_L g9759 ( 
.A(n_8889),
.Y(n_9759)
);

INVx2_ASAP7_75t_SL g9760 ( 
.A(n_8820),
.Y(n_9760)
);

INVx4_ASAP7_75t_L g9761 ( 
.A(n_8820),
.Y(n_9761)
);

INVx2_ASAP7_75t_L g9762 ( 
.A(n_8723),
.Y(n_9762)
);

INVx2_ASAP7_75t_L g9763 ( 
.A(n_8723),
.Y(n_9763)
);

NOR2xp33_ASAP7_75t_L g9764 ( 
.A(n_8727),
.B(n_203),
.Y(n_9764)
);

NAND2xp5_ASAP7_75t_SL g9765 ( 
.A(n_9034),
.B(n_204),
.Y(n_9765)
);

NAND2xp5_ASAP7_75t_L g9766 ( 
.A(n_8729),
.B(n_55),
.Y(n_9766)
);

INVx1_ASAP7_75t_L g9767 ( 
.A(n_8889),
.Y(n_9767)
);

NAND2xp5_ASAP7_75t_L g9768 ( 
.A(n_8729),
.B(n_55),
.Y(n_9768)
);

INVx1_ASAP7_75t_L g9769 ( 
.A(n_8889),
.Y(n_9769)
);

AND2x2_ASAP7_75t_L g9770 ( 
.A(n_8732),
.B(n_204),
.Y(n_9770)
);

NAND2xp5_ASAP7_75t_L g9771 ( 
.A(n_8729),
.B(n_56),
.Y(n_9771)
);

INVx3_ASAP7_75t_L g9772 ( 
.A(n_8820),
.Y(n_9772)
);

INVx1_ASAP7_75t_SL g9773 ( 
.A(n_9098),
.Y(n_9773)
);

INVx1_ASAP7_75t_L g9774 ( 
.A(n_8889),
.Y(n_9774)
);

OAI21xp5_ASAP7_75t_L g9775 ( 
.A1(n_9131),
.A2(n_56),
.B(n_57),
.Y(n_9775)
);

HB1xp67_ASAP7_75t_L g9776 ( 
.A(n_8830),
.Y(n_9776)
);

INVx1_ASAP7_75t_SL g9777 ( 
.A(n_9098),
.Y(n_9777)
);

NAND2xp5_ASAP7_75t_L g9778 ( 
.A(n_8729),
.B(n_56),
.Y(n_9778)
);

NAND2xp5_ASAP7_75t_SL g9779 ( 
.A(n_9034),
.B(n_205),
.Y(n_9779)
);

NOR2xp33_ASAP7_75t_L g9780 ( 
.A(n_8727),
.B(n_205),
.Y(n_9780)
);

AND2x2_ASAP7_75t_L g9781 ( 
.A(n_8732),
.B(n_206),
.Y(n_9781)
);

HB1xp67_ASAP7_75t_L g9782 ( 
.A(n_8830),
.Y(n_9782)
);

INVx1_ASAP7_75t_L g9783 ( 
.A(n_8889),
.Y(n_9783)
);

BUFx6f_ASAP7_75t_L g9784 ( 
.A(n_8820),
.Y(n_9784)
);

INVx1_ASAP7_75t_L g9785 ( 
.A(n_8889),
.Y(n_9785)
);

NAND2xp5_ASAP7_75t_L g9786 ( 
.A(n_8729),
.B(n_58),
.Y(n_9786)
);

INVx1_ASAP7_75t_L g9787 ( 
.A(n_8889),
.Y(n_9787)
);

INVx3_ASAP7_75t_L g9788 ( 
.A(n_8820),
.Y(n_9788)
);

INVxp67_ASAP7_75t_L g9789 ( 
.A(n_8787),
.Y(n_9789)
);

CKINVDCx5p33_ASAP7_75t_R g9790 ( 
.A(n_8836),
.Y(n_9790)
);

INVx1_ASAP7_75t_L g9791 ( 
.A(n_8889),
.Y(n_9791)
);

INVx1_ASAP7_75t_L g9792 ( 
.A(n_8889),
.Y(n_9792)
);

OAI21xp5_ASAP7_75t_L g9793 ( 
.A1(n_9131),
.A2(n_58),
.B(n_59),
.Y(n_9793)
);

AND2x2_ASAP7_75t_L g9794 ( 
.A(n_8732),
.B(n_207),
.Y(n_9794)
);

INVx3_ASAP7_75t_L g9795 ( 
.A(n_8820),
.Y(n_9795)
);

INVx1_ASAP7_75t_L g9796 ( 
.A(n_8889),
.Y(n_9796)
);

BUFx3_ASAP7_75t_L g9797 ( 
.A(n_9054),
.Y(n_9797)
);

NAND2xp5_ASAP7_75t_L g9798 ( 
.A(n_8729),
.B(n_59),
.Y(n_9798)
);

NOR2xp33_ASAP7_75t_L g9799 ( 
.A(n_8727),
.B(n_208),
.Y(n_9799)
);

NAND2xp5_ASAP7_75t_L g9800 ( 
.A(n_8729),
.B(n_59),
.Y(n_9800)
);

INVxp67_ASAP7_75t_SL g9801 ( 
.A(n_8830),
.Y(n_9801)
);

INVx2_ASAP7_75t_L g9802 ( 
.A(n_8723),
.Y(n_9802)
);

BUFx3_ASAP7_75t_L g9803 ( 
.A(n_9054),
.Y(n_9803)
);

NAND2xp5_ASAP7_75t_L g9804 ( 
.A(n_8729),
.B(n_60),
.Y(n_9804)
);

AND2x2_ASAP7_75t_L g9805 ( 
.A(n_8732),
.B(n_209),
.Y(n_9805)
);

INVx1_ASAP7_75t_L g9806 ( 
.A(n_8889),
.Y(n_9806)
);

INVx3_ASAP7_75t_L g9807 ( 
.A(n_8820),
.Y(n_9807)
);

BUFx3_ASAP7_75t_L g9808 ( 
.A(n_9054),
.Y(n_9808)
);

HB1xp67_ASAP7_75t_L g9809 ( 
.A(n_8830),
.Y(n_9809)
);

NAND2xp5_ASAP7_75t_L g9810 ( 
.A(n_8729),
.B(n_60),
.Y(n_9810)
);

AND2x2_ASAP7_75t_L g9811 ( 
.A(n_8732),
.B(n_210),
.Y(n_9811)
);

INVx2_ASAP7_75t_L g9812 ( 
.A(n_8723),
.Y(n_9812)
);

HB1xp67_ASAP7_75t_L g9813 ( 
.A(n_8830),
.Y(n_9813)
);

INVx2_ASAP7_75t_L g9814 ( 
.A(n_8723),
.Y(n_9814)
);

AND2x4_ASAP7_75t_L g9815 ( 
.A(n_8899),
.B(n_210),
.Y(n_9815)
);

AND2x2_ASAP7_75t_L g9816 ( 
.A(n_8732),
.B(n_211),
.Y(n_9816)
);

INVx1_ASAP7_75t_L g9817 ( 
.A(n_8889),
.Y(n_9817)
);

AND2x2_ASAP7_75t_L g9818 ( 
.A(n_8732),
.B(n_211),
.Y(n_9818)
);

AND2x2_ASAP7_75t_L g9819 ( 
.A(n_8732),
.B(n_212),
.Y(n_9819)
);

INVx3_ASAP7_75t_L g9820 ( 
.A(n_8820),
.Y(n_9820)
);

INVx1_ASAP7_75t_L g9821 ( 
.A(n_8889),
.Y(n_9821)
);

INVx1_ASAP7_75t_L g9822 ( 
.A(n_8889),
.Y(n_9822)
);

OR2x2_ASAP7_75t_L g9823 ( 
.A(n_8830),
.B(n_61),
.Y(n_9823)
);

INVx2_ASAP7_75t_L g9824 ( 
.A(n_8723),
.Y(n_9824)
);

AND2x2_ASAP7_75t_L g9825 ( 
.A(n_8732),
.B(n_212),
.Y(n_9825)
);

NOR2xp67_ASAP7_75t_L g9826 ( 
.A(n_9090),
.B(n_61),
.Y(n_9826)
);

NAND2xp5_ASAP7_75t_L g9827 ( 
.A(n_8729),
.B(n_61),
.Y(n_9827)
);

NOR2xp33_ASAP7_75t_L g9828 ( 
.A(n_8727),
.B(n_213),
.Y(n_9828)
);

INVx2_ASAP7_75t_L g9829 ( 
.A(n_8723),
.Y(n_9829)
);

NAND2xp5_ASAP7_75t_L g9830 ( 
.A(n_8729),
.B(n_62),
.Y(n_9830)
);

INVx2_ASAP7_75t_L g9831 ( 
.A(n_8723),
.Y(n_9831)
);

INVx3_ASAP7_75t_L g9832 ( 
.A(n_8820),
.Y(n_9832)
);

NAND2xp5_ASAP7_75t_L g9833 ( 
.A(n_8729),
.B(n_62),
.Y(n_9833)
);

AND2x4_ASAP7_75t_L g9834 ( 
.A(n_8899),
.B(n_213),
.Y(n_9834)
);

INVx2_ASAP7_75t_SL g9835 ( 
.A(n_8820),
.Y(n_9835)
);

AND2x2_ASAP7_75t_L g9836 ( 
.A(n_8732),
.B(n_214),
.Y(n_9836)
);

INVx3_ASAP7_75t_L g9837 ( 
.A(n_9761),
.Y(n_9837)
);

BUFx4f_ASAP7_75t_L g9838 ( 
.A(n_9784),
.Y(n_9838)
);

AOI21xp5_ASAP7_75t_L g9839 ( 
.A1(n_9258),
.A2(n_215),
.B(n_214),
.Y(n_9839)
);

NAND2xp5_ASAP7_75t_SL g9840 ( 
.A(n_9347),
.B(n_215),
.Y(n_9840)
);

AOI21xp5_ASAP7_75t_L g9841 ( 
.A1(n_9260),
.A2(n_217),
.B(n_216),
.Y(n_9841)
);

INVx2_ASAP7_75t_SL g9842 ( 
.A(n_9307),
.Y(n_9842)
);

AOI21xp5_ASAP7_75t_L g9843 ( 
.A1(n_9534),
.A2(n_9437),
.B(n_9465),
.Y(n_9843)
);

NOR3xp33_ASAP7_75t_L g9844 ( 
.A(n_9431),
.B(n_63),
.C(n_64),
.Y(n_9844)
);

A2O1A1Ixp33_ASAP7_75t_L g9845 ( 
.A1(n_9510),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_9845)
);

INVxp67_ASAP7_75t_L g9846 ( 
.A(n_9319),
.Y(n_9846)
);

NAND2xp5_ASAP7_75t_SL g9847 ( 
.A(n_9649),
.B(n_216),
.Y(n_9847)
);

NOR2xp33_ASAP7_75t_L g9848 ( 
.A(n_9605),
.B(n_217),
.Y(n_9848)
);

INVx3_ASAP7_75t_L g9849 ( 
.A(n_9784),
.Y(n_9849)
);

NAND2xp5_ASAP7_75t_L g9850 ( 
.A(n_9254),
.B(n_63),
.Y(n_9850)
);

NAND2xp5_ASAP7_75t_L g9851 ( 
.A(n_9257),
.B(n_65),
.Y(n_9851)
);

NAND2xp5_ASAP7_75t_L g9852 ( 
.A(n_9801),
.B(n_66),
.Y(n_9852)
);

INVx4_ASAP7_75t_L g9853 ( 
.A(n_9749),
.Y(n_9853)
);

A2O1A1Ixp33_ASAP7_75t_L g9854 ( 
.A1(n_9775),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_9854)
);

AOI21xp5_ASAP7_75t_L g9855 ( 
.A1(n_9263),
.A2(n_219),
.B(n_218),
.Y(n_9855)
);

INVx2_ASAP7_75t_L g9856 ( 
.A(n_9241),
.Y(n_9856)
);

AOI21xp5_ASAP7_75t_L g9857 ( 
.A1(n_9343),
.A2(n_220),
.B(n_219),
.Y(n_9857)
);

AOI21xp5_ASAP7_75t_L g9858 ( 
.A1(n_9356),
.A2(n_222),
.B(n_221),
.Y(n_9858)
);

AOI22xp5_ASAP7_75t_L g9859 ( 
.A1(n_9607),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_9859)
);

NAND2xp5_ASAP7_75t_L g9860 ( 
.A(n_9247),
.B(n_67),
.Y(n_9860)
);

NAND2xp5_ASAP7_75t_L g9861 ( 
.A(n_9273),
.B(n_68),
.Y(n_9861)
);

NAND2xp33_ASAP7_75t_L g9862 ( 
.A(n_9471),
.B(n_221),
.Y(n_9862)
);

O2A1O1Ixp33_ASAP7_75t_L g9863 ( 
.A1(n_9764),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_9863)
);

OAI21xp5_ASAP7_75t_L g9864 ( 
.A1(n_9780),
.A2(n_69),
.B(n_70),
.Y(n_9864)
);

NOR2x1_ASAP7_75t_L g9865 ( 
.A(n_9439),
.B(n_69),
.Y(n_9865)
);

A2O1A1Ixp33_ASAP7_75t_L g9866 ( 
.A1(n_9793),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_9866)
);

NAND2xp5_ASAP7_75t_SL g9867 ( 
.A(n_9473),
.B(n_222),
.Y(n_9867)
);

AOI21xp5_ASAP7_75t_L g9868 ( 
.A1(n_9367),
.A2(n_224),
.B(n_223),
.Y(n_9868)
);

AOI21x1_ASAP7_75t_L g9869 ( 
.A1(n_9652),
.A2(n_72),
.B(n_73),
.Y(n_9869)
);

AOI21xp5_ASAP7_75t_L g9870 ( 
.A1(n_9499),
.A2(n_224),
.B(n_223),
.Y(n_9870)
);

NAND2xp5_ASAP7_75t_L g9871 ( 
.A(n_9758),
.B(n_73),
.Y(n_9871)
);

INVxp67_ASAP7_75t_L g9872 ( 
.A(n_9679),
.Y(n_9872)
);

BUFx10_ASAP7_75t_L g9873 ( 
.A(n_9790),
.Y(n_9873)
);

OAI21xp5_ASAP7_75t_L g9874 ( 
.A1(n_9799),
.A2(n_74),
.B(n_75),
.Y(n_9874)
);

OAI21xp5_ASAP7_75t_L g9875 ( 
.A1(n_9828),
.A2(n_74),
.B(n_75),
.Y(n_9875)
);

AOI21xp5_ASAP7_75t_L g9876 ( 
.A1(n_9460),
.A2(n_226),
.B(n_225),
.Y(n_9876)
);

AOI21xp5_ASAP7_75t_L g9877 ( 
.A1(n_9555),
.A2(n_228),
.B(n_226),
.Y(n_9877)
);

AOI21xp5_ASAP7_75t_L g9878 ( 
.A1(n_9710),
.A2(n_229),
.B(n_228),
.Y(n_9878)
);

O2A1O1Ixp33_ASAP7_75t_L g9879 ( 
.A1(n_9584),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_9879)
);

AOI21xp5_ASAP7_75t_L g9880 ( 
.A1(n_9600),
.A2(n_231),
.B(n_230),
.Y(n_9880)
);

AOI21xp5_ASAP7_75t_L g9881 ( 
.A1(n_9327),
.A2(n_231),
.B(n_230),
.Y(n_9881)
);

HB1xp67_ASAP7_75t_L g9882 ( 
.A(n_9242),
.Y(n_9882)
);

OAI21xp5_ASAP7_75t_L g9883 ( 
.A1(n_9385),
.A2(n_9275),
.B(n_9483),
.Y(n_9883)
);

NAND2xp5_ASAP7_75t_L g9884 ( 
.A(n_9759),
.B(n_76),
.Y(n_9884)
);

AOI21xp5_ASAP7_75t_L g9885 ( 
.A1(n_9629),
.A2(n_233),
.B(n_232),
.Y(n_9885)
);

NAND2xp5_ASAP7_75t_L g9886 ( 
.A(n_9767),
.B(n_76),
.Y(n_9886)
);

INVxp67_ASAP7_75t_L g9887 ( 
.A(n_9698),
.Y(n_9887)
);

INVx2_ASAP7_75t_L g9888 ( 
.A(n_9255),
.Y(n_9888)
);

AND2x4_ASAP7_75t_L g9889 ( 
.A(n_9261),
.B(n_233),
.Y(n_9889)
);

OAI21xp33_ASAP7_75t_L g9890 ( 
.A1(n_9708),
.A2(n_77),
.B(n_78),
.Y(n_9890)
);

NAND2xp5_ASAP7_75t_SL g9891 ( 
.A(n_9425),
.B(n_234),
.Y(n_9891)
);

AOI22xp33_ASAP7_75t_L g9892 ( 
.A1(n_9404),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_9892)
);

OAI321xp33_ASAP7_75t_L g9893 ( 
.A1(n_9563),
.A2(n_80),
.A3(n_82),
.B1(n_78),
.B2(n_79),
.C(n_81),
.Y(n_9893)
);

INVx2_ASAP7_75t_L g9894 ( 
.A(n_9262),
.Y(n_9894)
);

INVx1_ASAP7_75t_L g9895 ( 
.A(n_9286),
.Y(n_9895)
);

O2A1O1Ixp5_ASAP7_75t_L g9896 ( 
.A1(n_9422),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_9896)
);

AOI21xp5_ASAP7_75t_L g9897 ( 
.A1(n_9329),
.A2(n_9717),
.B(n_9713),
.Y(n_9897)
);

NAND2xp5_ASAP7_75t_L g9898 ( 
.A(n_9769),
.B(n_80),
.Y(n_9898)
);

AOI21xp5_ASAP7_75t_L g9899 ( 
.A1(n_9594),
.A2(n_235),
.B(n_234),
.Y(n_9899)
);

NAND2xp5_ASAP7_75t_SL g9900 ( 
.A(n_9425),
.B(n_235),
.Y(n_9900)
);

INVx2_ASAP7_75t_SL g9901 ( 
.A(n_9307),
.Y(n_9901)
);

INVx2_ASAP7_75t_L g9902 ( 
.A(n_9265),
.Y(n_9902)
);

AOI21xp5_ASAP7_75t_L g9903 ( 
.A1(n_9492),
.A2(n_237),
.B(n_236),
.Y(n_9903)
);

NAND2xp5_ASAP7_75t_L g9904 ( 
.A(n_9774),
.B(n_81),
.Y(n_9904)
);

NOR2xp33_ASAP7_75t_L g9905 ( 
.A(n_9252),
.B(n_236),
.Y(n_9905)
);

AOI21xp5_ASAP7_75t_L g9906 ( 
.A1(n_9445),
.A2(n_239),
.B(n_238),
.Y(n_9906)
);

NAND2xp5_ASAP7_75t_L g9907 ( 
.A(n_9783),
.B(n_82),
.Y(n_9907)
);

AOI21x1_ASAP7_75t_L g9908 ( 
.A1(n_9626),
.A2(n_82),
.B(n_83),
.Y(n_9908)
);

AOI21xp5_ASAP7_75t_L g9909 ( 
.A1(n_9746),
.A2(n_240),
.B(n_238),
.Y(n_9909)
);

INVx3_ASAP7_75t_L g9910 ( 
.A(n_9331),
.Y(n_9910)
);

NAND2xp5_ASAP7_75t_SL g9911 ( 
.A(n_9453),
.B(n_241),
.Y(n_9911)
);

NAND2xp33_ASAP7_75t_L g9912 ( 
.A(n_9662),
.B(n_241),
.Y(n_9912)
);

AND2x2_ASAP7_75t_L g9913 ( 
.A(n_9272),
.B(n_242),
.Y(n_9913)
);

AOI21xp5_ASAP7_75t_L g9914 ( 
.A1(n_9560),
.A2(n_244),
.B(n_243),
.Y(n_9914)
);

INVx2_ASAP7_75t_L g9915 ( 
.A(n_9291),
.Y(n_9915)
);

NAND2xp5_ASAP7_75t_SL g9916 ( 
.A(n_9468),
.B(n_243),
.Y(n_9916)
);

A2O1A1Ixp33_ASAP7_75t_L g9917 ( 
.A1(n_9716),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_9917)
);

AO21x1_ASAP7_75t_L g9918 ( 
.A1(n_9285),
.A2(n_83),
.B(n_85),
.Y(n_9918)
);

NAND2xp5_ASAP7_75t_L g9919 ( 
.A(n_9785),
.B(n_85),
.Y(n_9919)
);

NAND2xp5_ASAP7_75t_L g9920 ( 
.A(n_9787),
.B(n_86),
.Y(n_9920)
);

INVx1_ASAP7_75t_L g9921 ( 
.A(n_9290),
.Y(n_9921)
);

O2A1O1Ixp33_ASAP7_75t_L g9922 ( 
.A1(n_9316),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_9922)
);

AOI22xp33_ASAP7_75t_L g9923 ( 
.A1(n_9296),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_9923)
);

HB1xp67_ASAP7_75t_L g9924 ( 
.A(n_9776),
.Y(n_9924)
);

NOR2xp33_ASAP7_75t_L g9925 ( 
.A(n_9747),
.B(n_244),
.Y(n_9925)
);

AOI21xp5_ASAP7_75t_L g9926 ( 
.A1(n_9386),
.A2(n_246),
.B(n_245),
.Y(n_9926)
);

NAND2xp5_ASAP7_75t_SL g9927 ( 
.A(n_9264),
.B(n_245),
.Y(n_9927)
);

NAND2xp5_ASAP7_75t_L g9928 ( 
.A(n_9791),
.B(n_87),
.Y(n_9928)
);

OAI21xp33_ASAP7_75t_L g9929 ( 
.A1(n_9469),
.A2(n_88),
.B(n_90),
.Y(n_9929)
);

NOR2xp33_ASAP7_75t_L g9930 ( 
.A(n_9756),
.B(n_9773),
.Y(n_9930)
);

A2O1A1Ixp33_ASAP7_75t_L g9931 ( 
.A1(n_9686),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_9931)
);

AOI21x1_ASAP7_75t_L g9932 ( 
.A1(n_9582),
.A2(n_90),
.B(n_91),
.Y(n_9932)
);

NAND2xp5_ASAP7_75t_L g9933 ( 
.A(n_9792),
.B(n_9796),
.Y(n_9933)
);

NOR2xp67_ASAP7_75t_L g9934 ( 
.A(n_9430),
.B(n_91),
.Y(n_9934)
);

NAND2xp5_ASAP7_75t_L g9935 ( 
.A(n_9806),
.B(n_92),
.Y(n_9935)
);

NAND2xp5_ASAP7_75t_L g9936 ( 
.A(n_9817),
.B(n_93),
.Y(n_9936)
);

AOI22xp5_ASAP7_75t_L g9937 ( 
.A1(n_9395),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_9937)
);

AOI21xp5_ASAP7_75t_L g9938 ( 
.A1(n_9401),
.A2(n_247),
.B(n_246),
.Y(n_9938)
);

OAI22xp5_ASAP7_75t_L g9939 ( 
.A1(n_9732),
.A2(n_248),
.B1(n_249),
.B2(n_247),
.Y(n_9939)
);

NOR2xp33_ASAP7_75t_L g9940 ( 
.A(n_9777),
.B(n_248),
.Y(n_9940)
);

NAND2xp5_ASAP7_75t_L g9941 ( 
.A(n_9821),
.B(n_94),
.Y(n_9941)
);

NAND2xp5_ASAP7_75t_L g9942 ( 
.A(n_9822),
.B(n_94),
.Y(n_9942)
);

NAND2xp5_ASAP7_75t_SL g9943 ( 
.A(n_9505),
.B(n_250),
.Y(n_9943)
);

NOR2xp33_ASAP7_75t_L g9944 ( 
.A(n_9524),
.B(n_250),
.Y(n_9944)
);

NAND2xp5_ASAP7_75t_L g9945 ( 
.A(n_9782),
.B(n_95),
.Y(n_9945)
);

AOI21xp5_ASAP7_75t_L g9946 ( 
.A1(n_9417),
.A2(n_252),
.B(n_251),
.Y(n_9946)
);

INVx1_ASAP7_75t_L g9947 ( 
.A(n_9295),
.Y(n_9947)
);

NAND2xp5_ASAP7_75t_L g9948 ( 
.A(n_9809),
.B(n_95),
.Y(n_9948)
);

AOI21xp5_ASAP7_75t_L g9949 ( 
.A1(n_9624),
.A2(n_9638),
.B(n_9664),
.Y(n_9949)
);

OAI21xp5_ASAP7_75t_L g9950 ( 
.A1(n_9681),
.A2(n_9692),
.B(n_9693),
.Y(n_9950)
);

AOI21xp5_ASAP7_75t_L g9951 ( 
.A1(n_9813),
.A2(n_254),
.B(n_251),
.Y(n_9951)
);

O2A1O1Ixp33_ASAP7_75t_SL g9952 ( 
.A1(n_9734),
.A2(n_256),
.B(n_257),
.C(n_255),
.Y(n_9952)
);

INVx1_ASAP7_75t_L g9953 ( 
.A(n_9376),
.Y(n_9953)
);

HB1xp67_ASAP7_75t_L g9954 ( 
.A(n_9248),
.Y(n_9954)
);

NAND2xp5_ASAP7_75t_L g9955 ( 
.A(n_9244),
.B(n_96),
.Y(n_9955)
);

INVx4_ASAP7_75t_L g9956 ( 
.A(n_9348),
.Y(n_9956)
);

NAND2xp5_ASAP7_75t_L g9957 ( 
.A(n_9450),
.B(n_96),
.Y(n_9957)
);

NAND2xp5_ASAP7_75t_L g9958 ( 
.A(n_9249),
.B(n_9387),
.Y(n_9958)
);

O2A1O1Ixp33_ASAP7_75t_L g9959 ( 
.A1(n_9268),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_9959)
);

INVx2_ASAP7_75t_L g9960 ( 
.A(n_9292),
.Y(n_9960)
);

OAI21xp5_ASAP7_75t_L g9961 ( 
.A1(n_9743),
.A2(n_97),
.B(n_99),
.Y(n_9961)
);

NAND2xp5_ASAP7_75t_L g9962 ( 
.A(n_9416),
.B(n_99),
.Y(n_9962)
);

INVx2_ASAP7_75t_L g9963 ( 
.A(n_9299),
.Y(n_9963)
);

AOI21xp5_ASAP7_75t_L g9964 ( 
.A1(n_9650),
.A2(n_256),
.B(n_255),
.Y(n_9964)
);

AOI21xp5_ASAP7_75t_L g9965 ( 
.A1(n_9237),
.A2(n_258),
.B(n_257),
.Y(n_9965)
);

A2O1A1Ixp33_ASAP7_75t_L g9966 ( 
.A1(n_9579),
.A2(n_9591),
.B(n_9668),
.C(n_9643),
.Y(n_9966)
);

AOI21xp5_ASAP7_75t_L g9967 ( 
.A1(n_9634),
.A2(n_260),
.B(n_259),
.Y(n_9967)
);

AOI21xp5_ASAP7_75t_L g9968 ( 
.A1(n_9489),
.A2(n_262),
.B(n_261),
.Y(n_9968)
);

NOR2xp33_ASAP7_75t_L g9969 ( 
.A(n_9240),
.B(n_263),
.Y(n_9969)
);

NAND2xp5_ASAP7_75t_L g9970 ( 
.A(n_9434),
.B(n_99),
.Y(n_9970)
);

INVx1_ASAP7_75t_L g9971 ( 
.A(n_9463),
.Y(n_9971)
);

BUFx3_ASAP7_75t_L g9972 ( 
.A(n_9287),
.Y(n_9972)
);

OR2x2_ASAP7_75t_L g9973 ( 
.A(n_9467),
.B(n_263),
.Y(n_9973)
);

NOR2xp67_ASAP7_75t_L g9974 ( 
.A(n_9694),
.B(n_100),
.Y(n_9974)
);

AOI22xp33_ASAP7_75t_L g9975 ( 
.A1(n_9622),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_9975)
);

AOI21x1_ASAP7_75t_L g9976 ( 
.A1(n_9589),
.A2(n_100),
.B(n_101),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_9482),
.Y(n_9977)
);

INVx3_ASAP7_75t_L g9978 ( 
.A(n_9331),
.Y(n_9978)
);

NAND3xp33_ASAP7_75t_L g9979 ( 
.A(n_9596),
.B(n_101),
.C(n_102),
.Y(n_9979)
);

BUFx6f_ASAP7_75t_L g9980 ( 
.A(n_9287),
.Y(n_9980)
);

NAND2xp5_ASAP7_75t_L g9981 ( 
.A(n_9490),
.B(n_102),
.Y(n_9981)
);

HB1xp67_ASAP7_75t_L g9982 ( 
.A(n_9488),
.Y(n_9982)
);

INVx2_ASAP7_75t_SL g9983 ( 
.A(n_9334),
.Y(n_9983)
);

NOR2xp33_ASAP7_75t_L g9984 ( 
.A(n_9789),
.B(n_264),
.Y(n_9984)
);

NAND2xp5_ASAP7_75t_L g9985 ( 
.A(n_9276),
.B(n_103),
.Y(n_9985)
);

AOI21xp5_ASAP7_75t_L g9986 ( 
.A1(n_9628),
.A2(n_266),
.B(n_265),
.Y(n_9986)
);

NAND2xp5_ASAP7_75t_L g9987 ( 
.A(n_9278),
.B(n_103),
.Y(n_9987)
);

AOI21xp5_ASAP7_75t_L g9988 ( 
.A1(n_9750),
.A2(n_9754),
.B(n_9751),
.Y(n_9988)
);

O2A1O1Ixp33_ASAP7_75t_L g9989 ( 
.A1(n_9752),
.A2(n_9779),
.B(n_9765),
.C(n_9705),
.Y(n_9989)
);

HB1xp67_ASAP7_75t_L g9990 ( 
.A(n_9625),
.Y(n_9990)
);

INVx2_ASAP7_75t_L g9991 ( 
.A(n_9305),
.Y(n_9991)
);

NAND2xp5_ASAP7_75t_L g9992 ( 
.A(n_9280),
.B(n_103),
.Y(n_9992)
);

AOI21xp5_ASAP7_75t_L g9993 ( 
.A1(n_9766),
.A2(n_267),
.B(n_265),
.Y(n_9993)
);

NOR2xp33_ASAP7_75t_L g9994 ( 
.A(n_9695),
.B(n_267),
.Y(n_9994)
);

CKINVDCx8_ASAP7_75t_R g9995 ( 
.A(n_9410),
.Y(n_9995)
);

OAI22xp5_ASAP7_75t_L g9996 ( 
.A1(n_9730),
.A2(n_269),
.B1(n_270),
.B2(n_268),
.Y(n_9996)
);

NAND2xp5_ASAP7_75t_L g9997 ( 
.A(n_9282),
.B(n_104),
.Y(n_9997)
);

AND2x4_ASAP7_75t_L g9998 ( 
.A(n_9411),
.B(n_268),
.Y(n_9998)
);

NAND2xp5_ASAP7_75t_L g9999 ( 
.A(n_9297),
.B(n_104),
.Y(n_9999)
);

AO32x1_ASAP7_75t_L g10000 ( 
.A1(n_9289),
.A2(n_107),
.A3(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_10000)
);

INVx1_ASAP7_75t_L g10001 ( 
.A(n_9512),
.Y(n_10001)
);

INVx1_ASAP7_75t_L g10002 ( 
.A(n_9301),
.Y(n_10002)
);

AND2x2_ASAP7_75t_L g10003 ( 
.A(n_9748),
.B(n_269),
.Y(n_10003)
);

HB1xp67_ASAP7_75t_L g10004 ( 
.A(n_9562),
.Y(n_10004)
);

INVx1_ASAP7_75t_L g10005 ( 
.A(n_9302),
.Y(n_10005)
);

OAI21xp5_ASAP7_75t_L g10006 ( 
.A1(n_9598),
.A2(n_105),
.B(n_107),
.Y(n_10006)
);

O2A1O1Ixp33_ASAP7_75t_L g10007 ( 
.A1(n_9735),
.A2(n_108),
.B(n_105),
.C(n_107),
.Y(n_10007)
);

NAND3xp33_ASAP7_75t_L g10008 ( 
.A(n_9461),
.B(n_109),
.C(n_110),
.Y(n_10008)
);

O2A1O1Ixp33_ASAP7_75t_L g10009 ( 
.A1(n_9298),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_10009)
);

HB1xp67_ASAP7_75t_L g10010 ( 
.A(n_9304),
.Y(n_10010)
);

NAND2xp5_ASAP7_75t_L g10011 ( 
.A(n_9335),
.B(n_109),
.Y(n_10011)
);

NAND2xp5_ASAP7_75t_L g10012 ( 
.A(n_9337),
.B(n_110),
.Y(n_10012)
);

NAND2xp5_ASAP7_75t_L g10013 ( 
.A(n_9353),
.B(n_111),
.Y(n_10013)
);

A2O1A1Ixp33_ASAP7_75t_L g10014 ( 
.A1(n_9462),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_10014)
);

NAND3xp33_ASAP7_75t_L g10015 ( 
.A(n_9651),
.B(n_112),
.C(n_113),
.Y(n_10015)
);

AOI21xp5_ASAP7_75t_L g10016 ( 
.A1(n_9768),
.A2(n_271),
.B(n_270),
.Y(n_10016)
);

OAI21xp33_ASAP7_75t_L g10017 ( 
.A1(n_9725),
.A2(n_113),
.B(n_114),
.Y(n_10017)
);

OAI21xp5_ASAP7_75t_L g10018 ( 
.A1(n_9293),
.A2(n_114),
.B(n_115),
.Y(n_10018)
);

AOI21xp5_ASAP7_75t_L g10019 ( 
.A1(n_9771),
.A2(n_272),
.B(n_271),
.Y(n_10019)
);

NAND2xp5_ASAP7_75t_L g10020 ( 
.A(n_9370),
.B(n_114),
.Y(n_10020)
);

NOR3xp33_ASAP7_75t_L g10021 ( 
.A(n_9711),
.B(n_115),
.C(n_116),
.Y(n_10021)
);

OAI21xp5_ASAP7_75t_L g10022 ( 
.A1(n_9313),
.A2(n_115),
.B(n_116),
.Y(n_10022)
);

OAI21x1_ASAP7_75t_L g10023 ( 
.A1(n_9604),
.A2(n_116),
.B(n_117),
.Y(n_10023)
);

A2O1A1Ixp33_ASAP7_75t_L g10024 ( 
.A1(n_9721),
.A2(n_9744),
.B(n_9678),
.C(n_9446),
.Y(n_10024)
);

AOI21xp5_ASAP7_75t_L g10025 ( 
.A1(n_9778),
.A2(n_274),
.B(n_273),
.Y(n_10025)
);

INVx1_ASAP7_75t_L g10026 ( 
.A(n_9372),
.Y(n_10026)
);

NAND2xp5_ASAP7_75t_SL g10027 ( 
.A(n_9621),
.B(n_273),
.Y(n_10027)
);

O2A1O1Ixp33_ASAP7_75t_L g10028 ( 
.A1(n_9311),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_10028)
);

AOI21xp5_ASAP7_75t_L g10029 ( 
.A1(n_9786),
.A2(n_275),
.B(n_274),
.Y(n_10029)
);

NOR3xp33_ASAP7_75t_L g10030 ( 
.A(n_9332),
.B(n_117),
.C(n_118),
.Y(n_10030)
);

NAND2xp5_ASAP7_75t_L g10031 ( 
.A(n_9379),
.B(n_118),
.Y(n_10031)
);

AOI21xp5_ASAP7_75t_L g10032 ( 
.A1(n_9798),
.A2(n_276),
.B(n_275),
.Y(n_10032)
);

NAND2xp5_ASAP7_75t_L g10033 ( 
.A(n_9380),
.B(n_119),
.Y(n_10033)
);

AOI21xp33_ASAP7_75t_L g10034 ( 
.A1(n_9690),
.A2(n_120),
.B(n_121),
.Y(n_10034)
);

NOR3xp33_ASAP7_75t_L g10035 ( 
.A(n_9673),
.B(n_120),
.C(n_121),
.Y(n_10035)
);

NAND3xp33_ASAP7_75t_L g10036 ( 
.A(n_9726),
.B(n_120),
.C(n_121),
.Y(n_10036)
);

O2A1O1Ixp33_ASAP7_75t_L g10037 ( 
.A1(n_9364),
.A2(n_122),
.B(n_277),
.C(n_276),
.Y(n_10037)
);

INVx3_ASAP7_75t_L g10038 ( 
.A(n_9334),
.Y(n_10038)
);

INVx2_ASAP7_75t_L g10039 ( 
.A(n_9308),
.Y(n_10039)
);

OAI21x1_ASAP7_75t_L g10040 ( 
.A1(n_9423),
.A2(n_122),
.B(n_278),
.Y(n_10040)
);

NOR2xp33_ASAP7_75t_L g10041 ( 
.A(n_9350),
.B(n_278),
.Y(n_10041)
);

NOR2x1_ASAP7_75t_L g10042 ( 
.A(n_9521),
.B(n_122),
.Y(n_10042)
);

AOI21xp5_ASAP7_75t_L g10043 ( 
.A1(n_9800),
.A2(n_279),
.B(n_280),
.Y(n_10043)
);

INVx1_ASAP7_75t_L g10044 ( 
.A(n_9382),
.Y(n_10044)
);

INVx1_ASAP7_75t_L g10045 ( 
.A(n_9388),
.Y(n_10045)
);

A2O1A1Ixp33_ASAP7_75t_L g10046 ( 
.A1(n_9568),
.A2(n_282),
.B(n_279),
.C(n_281),
.Y(n_10046)
);

AOI21xp5_ASAP7_75t_L g10047 ( 
.A1(n_9804),
.A2(n_281),
.B(n_282),
.Y(n_10047)
);

NAND2xp5_ASAP7_75t_L g10048 ( 
.A(n_9393),
.B(n_283),
.Y(n_10048)
);

A2O1A1Ixp33_ASAP7_75t_L g10049 ( 
.A1(n_9578),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_10049)
);

OAI21xp5_ASAP7_75t_L g10050 ( 
.A1(n_9654),
.A2(n_285),
.B(n_286),
.Y(n_10050)
);

BUFx12f_ASAP7_75t_L g10051 ( 
.A(n_9341),
.Y(n_10051)
);

AOI21xp5_ASAP7_75t_L g10052 ( 
.A1(n_9810),
.A2(n_286),
.B(n_287),
.Y(n_10052)
);

AOI21xp5_ASAP7_75t_L g10053 ( 
.A1(n_9827),
.A2(n_287),
.B(n_288),
.Y(n_10053)
);

AOI21x1_ASAP7_75t_L g10054 ( 
.A1(n_9613),
.A2(n_288),
.B(n_289),
.Y(n_10054)
);

AND2x2_ASAP7_75t_SL g10055 ( 
.A(n_9279),
.B(n_290),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_L g10056 ( 
.A(n_9432),
.B(n_290),
.Y(n_10056)
);

BUFx3_ASAP7_75t_L g10057 ( 
.A(n_9318),
.Y(n_10057)
);

OAI321xp33_ASAP7_75t_L g10058 ( 
.A1(n_9699),
.A2(n_9315),
.A3(n_9541),
.B1(n_9373),
.B2(n_9368),
.C(n_9706),
.Y(n_10058)
);

AOI21xp5_ASAP7_75t_L g10059 ( 
.A1(n_9830),
.A2(n_9833),
.B(n_9532),
.Y(n_10059)
);

NOR2xp33_ASAP7_75t_L g10060 ( 
.A(n_9728),
.B(n_291),
.Y(n_10060)
);

AOI21xp5_ASAP7_75t_L g10061 ( 
.A1(n_9586),
.A2(n_291),
.B(n_292),
.Y(n_10061)
);

NAND2xp5_ASAP7_75t_L g10062 ( 
.A(n_9424),
.B(n_292),
.Y(n_10062)
);

NOR2xp33_ASAP7_75t_L g10063 ( 
.A(n_9454),
.B(n_293),
.Y(n_10063)
);

AOI21xp5_ASAP7_75t_L g10064 ( 
.A1(n_9593),
.A2(n_294),
.B(n_295),
.Y(n_10064)
);

NAND2xp5_ASAP7_75t_L g10065 ( 
.A(n_9427),
.B(n_294),
.Y(n_10065)
);

AOI21xp5_ASAP7_75t_L g10066 ( 
.A1(n_9357),
.A2(n_295),
.B(n_296),
.Y(n_10066)
);

NAND2xp5_ASAP7_75t_L g10067 ( 
.A(n_9436),
.B(n_297),
.Y(n_10067)
);

NAND2xp5_ASAP7_75t_SL g10068 ( 
.A(n_9621),
.B(n_297),
.Y(n_10068)
);

AOI21xp5_ASAP7_75t_L g10069 ( 
.A1(n_9259),
.A2(n_298),
.B(n_299),
.Y(n_10069)
);

OAI22xp5_ASAP7_75t_L g10070 ( 
.A1(n_9408),
.A2(n_9507),
.B1(n_9466),
.B2(n_9475),
.Y(n_10070)
);

INVx2_ASAP7_75t_L g10071 ( 
.A(n_9310),
.Y(n_10071)
);

NAND2xp5_ASAP7_75t_L g10072 ( 
.A(n_9438),
.B(n_298),
.Y(n_10072)
);

OAI22xp5_ASAP7_75t_L g10073 ( 
.A1(n_9677),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_10073)
);

AOI21xp5_ASAP7_75t_L g10074 ( 
.A1(n_9657),
.A2(n_300),
.B(n_301),
.Y(n_10074)
);

NAND2xp33_ASAP7_75t_L g10075 ( 
.A(n_9608),
.B(n_302),
.Y(n_10075)
);

NAND2xp5_ASAP7_75t_L g10076 ( 
.A(n_9448),
.B(n_302),
.Y(n_10076)
);

INVx2_ASAP7_75t_SL g10077 ( 
.A(n_9399),
.Y(n_10077)
);

AOI21xp5_ASAP7_75t_L g10078 ( 
.A1(n_9670),
.A2(n_9636),
.B(n_9474),
.Y(n_10078)
);

OAI21xp5_ASAP7_75t_L g10079 ( 
.A1(n_9742),
.A2(n_303),
.B(n_305),
.Y(n_10079)
);

NOR2xp33_ASAP7_75t_L g10080 ( 
.A(n_9616),
.B(n_303),
.Y(n_10080)
);

INVx1_ASAP7_75t_L g10081 ( 
.A(n_9452),
.Y(n_10081)
);

AO32x1_ASAP7_75t_L g10082 ( 
.A1(n_9545),
.A2(n_307),
.A3(n_305),
.B1(n_306),
.B2(n_308),
.Y(n_10082)
);

INVx3_ASAP7_75t_L g10083 ( 
.A(n_9309),
.Y(n_10083)
);

OAI21xp5_ASAP7_75t_L g10084 ( 
.A1(n_9745),
.A2(n_9703),
.B(n_9520),
.Y(n_10084)
);

NOR3xp33_ASAP7_75t_L g10085 ( 
.A(n_9736),
.B(n_306),
.C(n_307),
.Y(n_10085)
);

NAND2xp5_ASAP7_75t_L g10086 ( 
.A(n_9457),
.B(n_308),
.Y(n_10086)
);

CKINVDCx10_ASAP7_75t_R g10087 ( 
.A(n_9309),
.Y(n_10087)
);

NAND2xp5_ASAP7_75t_L g10088 ( 
.A(n_9478),
.B(n_309),
.Y(n_10088)
);

NOR2xp33_ASAP7_75t_L g10089 ( 
.A(n_9691),
.B(n_310),
.Y(n_10089)
);

NAND2xp5_ASAP7_75t_L g10090 ( 
.A(n_9479),
.B(n_311),
.Y(n_10090)
);

NAND2xp5_ASAP7_75t_L g10091 ( 
.A(n_9487),
.B(n_312),
.Y(n_10091)
);

OR2x6_ASAP7_75t_SL g10092 ( 
.A(n_9402),
.B(n_312),
.Y(n_10092)
);

OAI22xp5_ASAP7_75t_L g10093 ( 
.A1(n_9538),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_10093)
);

AOI21xp5_ASAP7_75t_L g10094 ( 
.A1(n_9470),
.A2(n_314),
.B(n_315),
.Y(n_10094)
);

AND2x2_ASAP7_75t_L g10095 ( 
.A(n_9753),
.B(n_316),
.Y(n_10095)
);

AND2x2_ASAP7_75t_L g10096 ( 
.A(n_9836),
.B(n_9757),
.Y(n_10096)
);

NOR2xp33_ASAP7_75t_SL g10097 ( 
.A(n_9528),
.B(n_316),
.Y(n_10097)
);

OAI21x1_ASAP7_75t_L g10098 ( 
.A1(n_9491),
.A2(n_317),
.B(n_318),
.Y(n_10098)
);

AND2x6_ASAP7_75t_SL g10099 ( 
.A(n_9444),
.B(n_317),
.Y(n_10099)
);

HB1xp67_ASAP7_75t_L g10100 ( 
.A(n_9595),
.Y(n_10100)
);

AOI21xp5_ASAP7_75t_L g10101 ( 
.A1(n_9599),
.A2(n_318),
.B(n_319),
.Y(n_10101)
);

AO22x1_ASAP7_75t_L g10102 ( 
.A1(n_9330),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_10102)
);

OAI22xp5_ASAP7_75t_L g10103 ( 
.A1(n_9709),
.A2(n_9715),
.B1(n_9288),
.B2(n_9508),
.Y(n_10103)
);

AOI21xp5_ASAP7_75t_L g10104 ( 
.A1(n_9374),
.A2(n_321),
.B(n_322),
.Y(n_10104)
);

OAI321xp33_ASAP7_75t_L g10105 ( 
.A1(n_9729),
.A2(n_324),
.A3(n_328),
.B1(n_322),
.B2(n_323),
.C(n_327),
.Y(n_10105)
);

INVx2_ASAP7_75t_L g10106 ( 
.A(n_9325),
.Y(n_10106)
);

NAND2xp5_ASAP7_75t_L g10107 ( 
.A(n_9642),
.B(n_323),
.Y(n_10107)
);

NAND2xp5_ASAP7_75t_L g10108 ( 
.A(n_9644),
.B(n_324),
.Y(n_10108)
);

INVx2_ASAP7_75t_L g10109 ( 
.A(n_9333),
.Y(n_10109)
);

INVx1_ASAP7_75t_L g10110 ( 
.A(n_9480),
.Y(n_10110)
);

OAI21xp5_ASAP7_75t_L g10111 ( 
.A1(n_9720),
.A2(n_328),
.B(n_329),
.Y(n_10111)
);

NAND2xp5_ASAP7_75t_L g10112 ( 
.A(n_9647),
.B(n_329),
.Y(n_10112)
);

O2A1O1Ixp33_ASAP7_75t_L g10113 ( 
.A1(n_9655),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_10113)
);

BUFx6f_ASAP7_75t_L g10114 ( 
.A(n_9348),
.Y(n_10114)
);

NAND2xp5_ASAP7_75t_L g10115 ( 
.A(n_9680),
.B(n_330),
.Y(n_10115)
);

AOI21x1_ASAP7_75t_L g10116 ( 
.A1(n_9667),
.A2(n_331),
.B(n_332),
.Y(n_10116)
);

NAND2xp5_ASAP7_75t_L g10117 ( 
.A(n_9314),
.B(n_333),
.Y(n_10117)
);

AOI21xp5_ASAP7_75t_L g10118 ( 
.A1(n_9381),
.A2(n_333),
.B(n_334),
.Y(n_10118)
);

NAND2xp5_ASAP7_75t_SL g10119 ( 
.A(n_9554),
.B(n_335),
.Y(n_10119)
);

NOR2xp33_ASAP7_75t_L g10120 ( 
.A(n_9707),
.B(n_335),
.Y(n_10120)
);

AOI21xp5_ASAP7_75t_L g10121 ( 
.A1(n_9383),
.A2(n_336),
.B(n_337),
.Y(n_10121)
);

NAND2xp5_ASAP7_75t_L g10122 ( 
.A(n_9477),
.B(n_337),
.Y(n_10122)
);

NAND2xp5_ASAP7_75t_SL g10123 ( 
.A(n_9554),
.B(n_338),
.Y(n_10123)
);

O2A1O1Ixp33_ASAP7_75t_L g10124 ( 
.A1(n_9688),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_10124)
);

AOI21xp5_ASAP7_75t_L g10125 ( 
.A1(n_9384),
.A2(n_339),
.B(n_341),
.Y(n_10125)
);

NOR2xp33_ASAP7_75t_L g10126 ( 
.A(n_9588),
.B(n_9267),
.Y(n_10126)
);

OAI21xp33_ASAP7_75t_L g10127 ( 
.A1(n_9719),
.A2(n_341),
.B(n_342),
.Y(n_10127)
);

OAI21xp5_ASAP7_75t_L g10128 ( 
.A1(n_9722),
.A2(n_342),
.B(n_343),
.Y(n_10128)
);

INVx2_ASAP7_75t_L g10129 ( 
.A(n_9336),
.Y(n_10129)
);

OAI21xp5_ASAP7_75t_L g10130 ( 
.A1(n_9700),
.A2(n_343),
.B(n_344),
.Y(n_10130)
);

AOI21xp5_ASAP7_75t_L g10131 ( 
.A1(n_9400),
.A2(n_344),
.B(n_345),
.Y(n_10131)
);

AOI22xp5_ASAP7_75t_L g10132 ( 
.A1(n_9646),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_10132)
);

INVx2_ASAP7_75t_SL g10133 ( 
.A(n_9399),
.Y(n_10133)
);

AND2x2_ASAP7_75t_L g10134 ( 
.A(n_9770),
.B(n_346),
.Y(n_10134)
);

NOR2x1_ASAP7_75t_L g10135 ( 
.A(n_9823),
.B(n_348),
.Y(n_10135)
);

NAND2x1p5_ASAP7_75t_L g10136 ( 
.A(n_9542),
.B(n_9245),
.Y(n_10136)
);

AOI21xp5_ASAP7_75t_L g10137 ( 
.A1(n_9419),
.A2(n_350),
.B(n_351),
.Y(n_10137)
);

O2A1O1Ixp33_ASAP7_75t_SL g10138 ( 
.A1(n_9271),
.A2(n_9407),
.B(n_9447),
.C(n_9623),
.Y(n_10138)
);

INVx2_ASAP7_75t_SL g10139 ( 
.A(n_9340),
.Y(n_10139)
);

NOR2xp33_ASAP7_75t_L g10140 ( 
.A(n_9281),
.B(n_350),
.Y(n_10140)
);

AND2x2_ASAP7_75t_SL g10141 ( 
.A(n_9378),
.B(n_351),
.Y(n_10141)
);

AOI21xp5_ASAP7_75t_L g10142 ( 
.A1(n_9421),
.A2(n_9529),
.B(n_9641),
.Y(n_10142)
);

INVx1_ASAP7_75t_SL g10143 ( 
.A(n_9284),
.Y(n_10143)
);

AND3x2_ASAP7_75t_L g10144 ( 
.A(n_9253),
.B(n_352),
.C(n_353),
.Y(n_10144)
);

INVx1_ASAP7_75t_L g10145 ( 
.A(n_9494),
.Y(n_10145)
);

AOI21xp5_ASAP7_75t_L g10146 ( 
.A1(n_9724),
.A2(n_352),
.B(n_354),
.Y(n_10146)
);

AOI21xp5_ASAP7_75t_L g10147 ( 
.A1(n_9739),
.A2(n_355),
.B(n_356),
.Y(n_10147)
);

AOI21xp5_ASAP7_75t_L g10148 ( 
.A1(n_9606),
.A2(n_355),
.B(n_356),
.Y(n_10148)
);

NOR2xp33_ASAP7_75t_L g10149 ( 
.A(n_9283),
.B(n_357),
.Y(n_10149)
);

AOI21xp5_ASAP7_75t_L g10150 ( 
.A1(n_9609),
.A2(n_358),
.B(n_359),
.Y(n_10150)
);

AOI21xp5_ASAP7_75t_L g10151 ( 
.A1(n_9239),
.A2(n_359),
.B(n_360),
.Y(n_10151)
);

AOI21xp5_ASAP7_75t_L g10152 ( 
.A1(n_9669),
.A2(n_360),
.B(n_361),
.Y(n_10152)
);

AOI21xp5_ASAP7_75t_L g10153 ( 
.A1(n_9635),
.A2(n_9648),
.B(n_9637),
.Y(n_10153)
);

AOI21xp5_ASAP7_75t_L g10154 ( 
.A1(n_9522),
.A2(n_361),
.B(n_362),
.Y(n_10154)
);

AOI21xp5_ASAP7_75t_L g10155 ( 
.A1(n_9548),
.A2(n_362),
.B(n_363),
.Y(n_10155)
);

AND2x4_ASAP7_75t_L g10156 ( 
.A(n_9411),
.B(n_363),
.Y(n_10156)
);

INVx2_ASAP7_75t_L g10157 ( 
.A(n_9338),
.Y(n_10157)
);

A2O1A1Ixp33_ASAP7_75t_L g10158 ( 
.A1(n_9701),
.A2(n_9523),
.B(n_9321),
.C(n_9663),
.Y(n_10158)
);

NAND2xp5_ASAP7_75t_L g10159 ( 
.A(n_9640),
.B(n_364),
.Y(n_10159)
);

BUFx12f_ASAP7_75t_L g10160 ( 
.A(n_9684),
.Y(n_10160)
);

OAI22xp5_ASAP7_75t_L g10161 ( 
.A1(n_9546),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_10161)
);

AND2x2_ASAP7_75t_L g10162 ( 
.A(n_9781),
.B(n_9794),
.Y(n_10162)
);

NAND2xp5_ASAP7_75t_L g10163 ( 
.A(n_9443),
.B(n_365),
.Y(n_10163)
);

OAI22x1_ASAP7_75t_L g10164 ( 
.A1(n_9602),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_10164)
);

INVx1_ASAP7_75t_L g10165 ( 
.A(n_9500),
.Y(n_10165)
);

AOI21xp5_ASAP7_75t_L g10166 ( 
.A1(n_9572),
.A2(n_368),
.B(n_369),
.Y(n_10166)
);

AOI21xp5_ASAP7_75t_L g10167 ( 
.A1(n_9456),
.A2(n_369),
.B(n_370),
.Y(n_10167)
);

AOI21x1_ASAP7_75t_L g10168 ( 
.A1(n_9671),
.A2(n_370),
.B(n_371),
.Y(n_10168)
);

NAND2xp5_ASAP7_75t_L g10169 ( 
.A(n_9375),
.B(n_371),
.Y(n_10169)
);

AOI21xp5_ASAP7_75t_L g10170 ( 
.A1(n_9723),
.A2(n_372),
.B(n_373),
.Y(n_10170)
);

AO21x1_ASAP7_75t_L g10171 ( 
.A1(n_9612),
.A2(n_372),
.B(n_373),
.Y(n_10171)
);

NOR2xp33_ASAP7_75t_L g10172 ( 
.A(n_9303),
.B(n_374),
.Y(n_10172)
);

INVx3_ASAP7_75t_L g10173 ( 
.A(n_9797),
.Y(n_10173)
);

A2O1A1Ixp33_ASAP7_75t_L g10174 ( 
.A1(n_9597),
.A2(n_9610),
.B(n_9476),
.C(n_9429),
.Y(n_10174)
);

OAI21xp33_ASAP7_75t_L g10175 ( 
.A1(n_9533),
.A2(n_374),
.B(n_375),
.Y(n_10175)
);

O2A1O1Ixp33_ASAP7_75t_L g10176 ( 
.A1(n_9552),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_10176)
);

AOI22xp33_ASAP7_75t_L g10177 ( 
.A1(n_9519),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_10177)
);

AOI21xp5_ASAP7_75t_L g10178 ( 
.A1(n_9653),
.A2(n_378),
.B(n_379),
.Y(n_10178)
);

INVx1_ASAP7_75t_SL g10179 ( 
.A(n_9358),
.Y(n_10179)
);

AOI21xp5_ASAP7_75t_L g10180 ( 
.A1(n_9661),
.A2(n_379),
.B(n_380),
.Y(n_10180)
);

NAND2xp5_ASAP7_75t_L g10181 ( 
.A(n_9398),
.B(n_380),
.Y(n_10181)
);

AOI21x1_ASAP7_75t_L g10182 ( 
.A1(n_9639),
.A2(n_382),
.B(n_383),
.Y(n_10182)
);

AOI21xp5_ASAP7_75t_L g10183 ( 
.A1(n_9666),
.A2(n_382),
.B(n_383),
.Y(n_10183)
);

NAND2xp5_ASAP7_75t_L g10184 ( 
.A(n_9330),
.B(n_384),
.Y(n_10184)
);

NOR2xp33_ASAP7_75t_L g10185 ( 
.A(n_9718),
.B(n_384),
.Y(n_10185)
);

NAND2xp5_ASAP7_75t_L g10186 ( 
.A(n_9330),
.B(n_385),
.Y(n_10186)
);

AND2x2_ASAP7_75t_L g10187 ( 
.A(n_9805),
.B(n_385),
.Y(n_10187)
);

HB1xp67_ASAP7_75t_L g10188 ( 
.A(n_9570),
.Y(n_10188)
);

NAND2xp5_ASAP7_75t_L g10189 ( 
.A(n_9349),
.B(n_386),
.Y(n_10189)
);

AOI21xp5_ASAP7_75t_L g10190 ( 
.A1(n_9685),
.A2(n_386),
.B(n_387),
.Y(n_10190)
);

AOI21x1_ASAP7_75t_L g10191 ( 
.A1(n_9415),
.A2(n_387),
.B(n_388),
.Y(n_10191)
);

AOI22xp5_ASAP7_75t_L g10192 ( 
.A1(n_9646),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_10192)
);

NAND2xp5_ASAP7_75t_L g10193 ( 
.A(n_9349),
.B(n_389),
.Y(n_10193)
);

AND2x2_ASAP7_75t_L g10194 ( 
.A(n_9811),
.B(n_390),
.Y(n_10194)
);

INVx2_ASAP7_75t_L g10195 ( 
.A(n_9339),
.Y(n_10195)
);

INVxp67_ASAP7_75t_L g10196 ( 
.A(n_9497),
.Y(n_10196)
);

AOI21xp5_ASAP7_75t_L g10197 ( 
.A1(n_9697),
.A2(n_391),
.B(n_392),
.Y(n_10197)
);

O2A1O1Ixp33_ASAP7_75t_L g10198 ( 
.A1(n_9361),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_10198)
);

NAND2xp5_ASAP7_75t_L g10199 ( 
.A(n_9349),
.B(n_395),
.Y(n_10199)
);

INVx2_ASAP7_75t_L g10200 ( 
.A(n_9345),
.Y(n_10200)
);

INVx3_ASAP7_75t_L g10201 ( 
.A(n_9803),
.Y(n_10201)
);

AND2x2_ASAP7_75t_L g10202 ( 
.A(n_9816),
.B(n_396),
.Y(n_10202)
);

INVx2_ASAP7_75t_L g10203 ( 
.A(n_9362),
.Y(n_10203)
);

INVx2_ASAP7_75t_SL g10204 ( 
.A(n_9451),
.Y(n_10204)
);

BUFx4f_ASAP7_75t_L g10205 ( 
.A(n_9410),
.Y(n_10205)
);

NAND2xp5_ASAP7_75t_L g10206 ( 
.A(n_9420),
.B(n_396),
.Y(n_10206)
);

AND2x4_ASAP7_75t_L g10207 ( 
.A(n_9558),
.B(n_397),
.Y(n_10207)
);

OR2x6_ASAP7_75t_L g10208 ( 
.A(n_9516),
.B(n_398),
.Y(n_10208)
);

INVx1_ASAP7_75t_L g10209 ( 
.A(n_9504),
.Y(n_10209)
);

NAND3xp33_ASAP7_75t_L g10210 ( 
.A(n_9351),
.B(n_399),
.C(n_400),
.Y(n_10210)
);

AND2x2_ASAP7_75t_L g10211 ( 
.A(n_9818),
.B(n_399),
.Y(n_10211)
);

INVx4_ASAP7_75t_L g10212 ( 
.A(n_9243),
.Y(n_10212)
);

NAND2xp5_ASAP7_75t_SL g10213 ( 
.A(n_9554),
.B(n_400),
.Y(n_10213)
);

NAND2xp5_ASAP7_75t_L g10214 ( 
.A(n_9420),
.B(n_9449),
.Y(n_10214)
);

NAND2xp5_ASAP7_75t_SL g10215 ( 
.A(n_9527),
.B(n_401),
.Y(n_10215)
);

AOI21xp5_ASAP7_75t_L g10216 ( 
.A1(n_9702),
.A2(n_401),
.B(n_402),
.Y(n_10216)
);

OAI22xp5_ASAP7_75t_L g10217 ( 
.A1(n_9615),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_10217)
);

AOI21xp5_ASAP7_75t_L g10218 ( 
.A1(n_9714),
.A2(n_403),
.B(n_404),
.Y(n_10218)
);

AOI21xp5_ASAP7_75t_L g10219 ( 
.A1(n_9727),
.A2(n_9731),
.B(n_9441),
.Y(n_10219)
);

O2A1O1Ixp33_ASAP7_75t_L g10220 ( 
.A1(n_9363),
.A2(n_9371),
.B(n_9526),
.C(n_9525),
.Y(n_10220)
);

INVx2_ASAP7_75t_L g10221 ( 
.A(n_9366),
.Y(n_10221)
);

NAND2xp5_ASAP7_75t_L g10222 ( 
.A(n_9420),
.B(n_405),
.Y(n_10222)
);

AOI21xp5_ASAP7_75t_L g10223 ( 
.A1(n_9614),
.A2(n_405),
.B(n_406),
.Y(n_10223)
);

NAND2xp5_ASAP7_75t_L g10224 ( 
.A(n_9344),
.B(n_407),
.Y(n_10224)
);

INVx1_ASAP7_75t_L g10225 ( 
.A(n_9506),
.Y(n_10225)
);

NAND2xp5_ASAP7_75t_SL g10226 ( 
.A(n_9527),
.B(n_407),
.Y(n_10226)
);

NAND2xp5_ASAP7_75t_L g10227 ( 
.A(n_9659),
.B(n_408),
.Y(n_10227)
);

AOI21xp5_ASAP7_75t_L g10228 ( 
.A1(n_9618),
.A2(n_9619),
.B(n_9683),
.Y(n_10228)
);

BUFx6f_ASAP7_75t_L g10229 ( 
.A(n_9808),
.Y(n_10229)
);

BUFx3_ASAP7_75t_L g10230 ( 
.A(n_9414),
.Y(n_10230)
);

AOI21xp5_ASAP7_75t_L g10231 ( 
.A1(n_9515),
.A2(n_9518),
.B(n_9481),
.Y(n_10231)
);

NAND2xp5_ASAP7_75t_L g10232 ( 
.A(n_9660),
.B(n_408),
.Y(n_10232)
);

OR2x6_ASAP7_75t_L g10233 ( 
.A(n_9516),
.B(n_409),
.Y(n_10233)
);

AOI21xp5_ASAP7_75t_L g10234 ( 
.A1(n_9342),
.A2(n_409),
.B(n_410),
.Y(n_10234)
);

INVx1_ASAP7_75t_L g10235 ( 
.A(n_9530),
.Y(n_10235)
);

NAND2xp5_ASAP7_75t_L g10236 ( 
.A(n_9277),
.B(n_411),
.Y(n_10236)
);

BUFx4f_ASAP7_75t_L g10237 ( 
.A(n_9549),
.Y(n_10237)
);

AOI21xp5_ASAP7_75t_L g10238 ( 
.A1(n_9712),
.A2(n_411),
.B(n_412),
.Y(n_10238)
);

NAND2xp5_ASAP7_75t_L g10239 ( 
.A(n_9519),
.B(n_412),
.Y(n_10239)
);

NAND2xp5_ASAP7_75t_L g10240 ( 
.A(n_9519),
.B(n_413),
.Y(n_10240)
);

NOR2xp33_ASAP7_75t_L g10241 ( 
.A(n_9656),
.B(n_9733),
.Y(n_10241)
);

BUFx2_ASAP7_75t_SL g10242 ( 
.A(n_9346),
.Y(n_10242)
);

CKINVDCx5p33_ASAP7_75t_R g10243 ( 
.A(n_9426),
.Y(n_10243)
);

INVx2_ASAP7_75t_L g10244 ( 
.A(n_9377),
.Y(n_10244)
);

NAND2xp5_ASAP7_75t_L g10245 ( 
.A(n_9312),
.B(n_413),
.Y(n_10245)
);

AOI21xp5_ASAP7_75t_L g10246 ( 
.A1(n_9740),
.A2(n_414),
.B(n_415),
.Y(n_10246)
);

NAND2xp5_ASAP7_75t_L g10247 ( 
.A(n_9306),
.B(n_414),
.Y(n_10247)
);

NAND2xp5_ASAP7_75t_L g10248 ( 
.A(n_9369),
.B(n_415),
.Y(n_10248)
);

INVxp67_ASAP7_75t_L g10249 ( 
.A(n_9536),
.Y(n_10249)
);

A2O1A1Ixp33_ASAP7_75t_L g10250 ( 
.A1(n_9617),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_10250)
);

NAND2xp5_ASAP7_75t_L g10251 ( 
.A(n_9819),
.B(n_416),
.Y(n_10251)
);

HB1xp67_ASAP7_75t_L g10252 ( 
.A(n_9573),
.Y(n_10252)
);

O2A1O1Ixp5_ASAP7_75t_L g10253 ( 
.A1(n_9741),
.A2(n_419),
.B(n_417),
.C(n_418),
.Y(n_10253)
);

AOI21xp5_ASAP7_75t_L g10254 ( 
.A1(n_9238),
.A2(n_420),
.B(n_421),
.Y(n_10254)
);

OAI22xp5_ASAP7_75t_L g10255 ( 
.A1(n_9633),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_10255)
);

INVx2_ASAP7_75t_L g10256 ( 
.A(n_9389),
.Y(n_10256)
);

AOI21xp5_ASAP7_75t_L g10257 ( 
.A1(n_9687),
.A2(n_423),
.B(n_424),
.Y(n_10257)
);

OAI22xp5_ASAP7_75t_L g10258 ( 
.A1(n_9682),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_10258)
);

NOR3xp33_ASAP7_75t_L g10259 ( 
.A(n_9550),
.B(n_425),
.C(n_426),
.Y(n_10259)
);

NOR2xp33_ASAP7_75t_R g10260 ( 
.A(n_9772),
.B(n_427),
.Y(n_10260)
);

NAND2xp5_ASAP7_75t_SL g10261 ( 
.A(n_9672),
.B(n_427),
.Y(n_10261)
);

HB1xp67_ASAP7_75t_L g10262 ( 
.A(n_9696),
.Y(n_10262)
);

NOR3xp33_ASAP7_75t_L g10263 ( 
.A(n_9632),
.B(n_428),
.C(n_429),
.Y(n_10263)
);

NAND2xp5_ASAP7_75t_L g10264 ( 
.A(n_9825),
.B(n_429),
.Y(n_10264)
);

NAND3xp33_ASAP7_75t_L g10265 ( 
.A(n_9580),
.B(n_430),
.C(n_431),
.Y(n_10265)
);

AOI21xp5_ASAP7_75t_L g10266 ( 
.A1(n_9502),
.A2(n_430),
.B(n_432),
.Y(n_10266)
);

NAND2xp5_ASAP7_75t_L g10267 ( 
.A(n_9294),
.B(n_433),
.Y(n_10267)
);

AOI21xp5_ASAP7_75t_L g10268 ( 
.A1(n_9503),
.A2(n_433),
.B(n_434),
.Y(n_10268)
);

OAI21xp5_ASAP7_75t_L g10269 ( 
.A1(n_9646),
.A2(n_434),
.B(n_435),
.Y(n_10269)
);

BUFx12f_ASAP7_75t_L g10270 ( 
.A(n_9269),
.Y(n_10270)
);

NAND2xp5_ASAP7_75t_L g10271 ( 
.A(n_9620),
.B(n_435),
.Y(n_10271)
);

AOI21xp5_ASAP7_75t_L g10272 ( 
.A1(n_9627),
.A2(n_436),
.B(n_437),
.Y(n_10272)
);

AOI21xp5_ASAP7_75t_L g10273 ( 
.A1(n_9630),
.A2(n_436),
.B(n_437),
.Y(n_10273)
);

BUFx3_ASAP7_75t_L g10274 ( 
.A(n_9365),
.Y(n_10274)
);

INVxp67_ASAP7_75t_L g10275 ( 
.A(n_9611),
.Y(n_10275)
);

NOR2xp67_ASAP7_75t_L g10276 ( 
.A(n_9493),
.B(n_438),
.Y(n_10276)
);

NAND2xp5_ASAP7_75t_L g10277 ( 
.A(n_9514),
.B(n_438),
.Y(n_10277)
);

OAI22xp5_ASAP7_75t_L g10278 ( 
.A1(n_9495),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_10278)
);

NAND2xp5_ASAP7_75t_L g10279 ( 
.A(n_9517),
.B(n_439),
.Y(n_10279)
);

OAI21xp5_ASAP7_75t_L g10280 ( 
.A1(n_9440),
.A2(n_441),
.B(n_442),
.Y(n_10280)
);

BUFx6f_ASAP7_75t_L g10281 ( 
.A(n_9394),
.Y(n_10281)
);

BUFx4f_ASAP7_75t_L g10282 ( 
.A(n_9788),
.Y(n_10282)
);

INVx1_ASAP7_75t_L g10283 ( 
.A(n_9531),
.Y(n_10283)
);

AOI21xp5_ASAP7_75t_L g10284 ( 
.A1(n_9631),
.A2(n_9645),
.B(n_9359),
.Y(n_10284)
);

NAND2xp33_ASAP7_75t_SL g10285 ( 
.A(n_9390),
.B(n_442),
.Y(n_10285)
);

A2O1A1Ixp33_ASAP7_75t_L g10286 ( 
.A1(n_9326),
.A2(n_446),
.B(n_444),
.C(n_445),
.Y(n_10286)
);

INVx1_ASAP7_75t_L g10287 ( 
.A(n_9535),
.Y(n_10287)
);

AOI21xp5_ASAP7_75t_L g10288 ( 
.A1(n_9539),
.A2(n_444),
.B(n_445),
.Y(n_10288)
);

OAI21xp5_ASAP7_75t_L g10289 ( 
.A1(n_9569),
.A2(n_446),
.B(n_447),
.Y(n_10289)
);

OAI22xp5_ASAP7_75t_L g10290 ( 
.A1(n_9704),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_10290)
);

OAI21xp5_ASAP7_75t_L g10291 ( 
.A1(n_9592),
.A2(n_448),
.B(n_449),
.Y(n_10291)
);

AOI21xp33_ASAP7_75t_L g10292 ( 
.A1(n_9603),
.A2(n_450),
.B(n_451),
.Y(n_10292)
);

A2O1A1Ixp33_ASAP7_75t_L g10293 ( 
.A1(n_9251),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_10293)
);

AOI21xp5_ASAP7_75t_L g10294 ( 
.A1(n_9540),
.A2(n_452),
.B(n_453),
.Y(n_10294)
);

INVx2_ASAP7_75t_SL g10295 ( 
.A(n_9451),
.Y(n_10295)
);

INVx2_ASAP7_75t_L g10296 ( 
.A(n_9392),
.Y(n_10296)
);

AND2x2_ASAP7_75t_L g10297 ( 
.A(n_9274),
.B(n_9581),
.Y(n_10297)
);

INVx1_ASAP7_75t_SL g10298 ( 
.A(n_9397),
.Y(n_10298)
);

NAND2xp5_ASAP7_75t_L g10299 ( 
.A(n_9511),
.B(n_453),
.Y(n_10299)
);

NAND2xp5_ASAP7_75t_L g10300 ( 
.A(n_9513),
.B(n_454),
.Y(n_10300)
);

NAND2xp5_ASAP7_75t_SL g10301 ( 
.A(n_9428),
.B(n_454),
.Y(n_10301)
);

NAND2xp5_ASAP7_75t_SL g10302 ( 
.A(n_9428),
.B(n_455),
.Y(n_10302)
);

AOI21xp5_ASAP7_75t_L g10303 ( 
.A1(n_9551),
.A2(n_455),
.B(n_456),
.Y(n_10303)
);

OAI21xp5_ASAP7_75t_L g10304 ( 
.A1(n_9553),
.A2(n_456),
.B(n_457),
.Y(n_10304)
);

NAND2xp5_ASAP7_75t_L g10305 ( 
.A(n_9266),
.B(n_458),
.Y(n_10305)
);

NAND2xp5_ASAP7_75t_L g10306 ( 
.A(n_9266),
.B(n_458),
.Y(n_10306)
);

OAI21xp5_ASAP7_75t_L g10307 ( 
.A1(n_9561),
.A2(n_459),
.B(n_460),
.Y(n_10307)
);

AOI21xp5_ASAP7_75t_L g10308 ( 
.A1(n_9556),
.A2(n_460),
.B(n_461),
.Y(n_10308)
);

AOI21xp5_ASAP7_75t_L g10309 ( 
.A1(n_9557),
.A2(n_462),
.B(n_463),
.Y(n_10309)
);

A2O1A1Ixp33_ASAP7_75t_L g10310 ( 
.A1(n_9826),
.A2(n_464),
.B(n_462),
.C(n_463),
.Y(n_10310)
);

NAND2xp5_ASAP7_75t_SL g10311 ( 
.A(n_9544),
.B(n_464),
.Y(n_10311)
);

INVx2_ASAP7_75t_L g10312 ( 
.A(n_9409),
.Y(n_10312)
);

NAND2xp5_ASAP7_75t_SL g10313 ( 
.A(n_9689),
.B(n_465),
.Y(n_10313)
);

INVx1_ASAP7_75t_L g10314 ( 
.A(n_9564),
.Y(n_10314)
);

INVx2_ASAP7_75t_L g10315 ( 
.A(n_9412),
.Y(n_10315)
);

BUFx3_ASAP7_75t_L g10316 ( 
.A(n_9246),
.Y(n_10316)
);

AOI22xp5_ASAP7_75t_L g10317 ( 
.A1(n_9266),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_10317)
);

INVx1_ASAP7_75t_L g10318 ( 
.A(n_9565),
.Y(n_10318)
);

OAI21xp5_ASAP7_75t_L g10319 ( 
.A1(n_9571),
.A2(n_467),
.B(n_468),
.Y(n_10319)
);

AOI21x1_ASAP7_75t_L g10320 ( 
.A1(n_9509),
.A2(n_469),
.B(n_470),
.Y(n_10320)
);

AOI21x1_ASAP7_75t_L g10321 ( 
.A1(n_9352),
.A2(n_469),
.B(n_470),
.Y(n_10321)
);

NAND2xp5_ASAP7_75t_SL g10322 ( 
.A(n_9658),
.B(n_471),
.Y(n_10322)
);

BUFx6f_ASAP7_75t_L g10323 ( 
.A(n_9256),
.Y(n_10323)
);

AOI22xp5_ASAP7_75t_L g10324 ( 
.A1(n_9601),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_10324)
);

AND2x2_ASAP7_75t_L g10325 ( 
.A(n_9250),
.B(n_472),
.Y(n_10325)
);

AOI21xp5_ASAP7_75t_L g10326 ( 
.A1(n_9577),
.A2(n_473),
.B(n_474),
.Y(n_10326)
);

AOI21xp5_ASAP7_75t_L g10327 ( 
.A1(n_9433),
.A2(n_474),
.B(n_475),
.Y(n_10327)
);

NAND2xp5_ASAP7_75t_L g10328 ( 
.A(n_9435),
.B(n_475),
.Y(n_10328)
);

AOI21xp5_ASAP7_75t_L g10329 ( 
.A1(n_9442),
.A2(n_476),
.B(n_477),
.Y(n_10329)
);

OAI22xp5_ASAP7_75t_L g10330 ( 
.A1(n_9738),
.A2(n_9674),
.B1(n_9486),
.B2(n_9455),
.Y(n_10330)
);

HB1xp67_ASAP7_75t_L g10331 ( 
.A(n_9459),
.Y(n_10331)
);

OAI321xp33_ASAP7_75t_L g10332 ( 
.A1(n_9458),
.A2(n_479),
.A3(n_481),
.B1(n_477),
.B2(n_478),
.C(n_480),
.Y(n_10332)
);

NAND2xp5_ASAP7_75t_SL g10333 ( 
.A(n_9658),
.B(n_9391),
.Y(n_10333)
);

INVx3_ASAP7_75t_L g10334 ( 
.A(n_9795),
.Y(n_10334)
);

AOI21xp5_ASAP7_75t_L g10335 ( 
.A1(n_9472),
.A2(n_478),
.B(n_482),
.Y(n_10335)
);

NAND2x1p5_ASAP7_75t_L g10336 ( 
.A(n_9807),
.B(n_482),
.Y(n_10336)
);

BUFx12f_ASAP7_75t_L g10337 ( 
.A(n_9760),
.Y(n_10337)
);

BUFx6f_ASAP7_75t_L g10338 ( 
.A(n_9820),
.Y(n_10338)
);

INVx1_ASAP7_75t_L g10339 ( 
.A(n_9485),
.Y(n_10339)
);

AOI22xp5_ASAP7_75t_L g10340 ( 
.A1(n_9676),
.A2(n_487),
.B1(n_484),
.B2(n_485),
.Y(n_10340)
);

BUFx6f_ASAP7_75t_L g10341 ( 
.A(n_9835),
.Y(n_10341)
);

NAND2xp5_ASAP7_75t_L g10342 ( 
.A(n_9501),
.B(n_484),
.Y(n_10342)
);

INVx2_ASAP7_75t_L g10343 ( 
.A(n_9537),
.Y(n_10343)
);

INVx2_ASAP7_75t_L g10344 ( 
.A(n_9543),
.Y(n_10344)
);

INVx3_ASAP7_75t_L g10345 ( 
.A(n_9832),
.Y(n_10345)
);

NAND2xp5_ASAP7_75t_L g10346 ( 
.A(n_9547),
.B(n_485),
.Y(n_10346)
);

OAI21xp5_ASAP7_75t_L g10347 ( 
.A1(n_9576),
.A2(n_487),
.B(n_488),
.Y(n_10347)
);

AOI21xp5_ASAP7_75t_L g10348 ( 
.A1(n_9559),
.A2(n_488),
.B(n_489),
.Y(n_10348)
);

A2O1A1Ixp33_ASAP7_75t_L g10349 ( 
.A1(n_9665),
.A2(n_491),
.B(n_489),
.C(n_490),
.Y(n_10349)
);

BUFx4f_ASAP7_75t_L g10350 ( 
.A(n_9815),
.Y(n_10350)
);

BUFx3_ASAP7_75t_L g10351 ( 
.A(n_9320),
.Y(n_10351)
);

NAND2xp5_ASAP7_75t_L g10352 ( 
.A(n_9567),
.B(n_9574),
.Y(n_10352)
);

AOI22xp5_ASAP7_75t_L g10353 ( 
.A1(n_9464),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_10353)
);

O2A1O1Ixp33_ASAP7_75t_SL g10354 ( 
.A1(n_9566),
.A2(n_494),
.B(n_492),
.C(n_493),
.Y(n_10354)
);

O2A1O1Ixp33_ASAP7_75t_SL g10355 ( 
.A1(n_9496),
.A2(n_496),
.B(n_493),
.C(n_495),
.Y(n_10355)
);

A2O1A1Ixp33_ASAP7_75t_L g10356 ( 
.A1(n_9675),
.A2(n_497),
.B(n_495),
.C(n_496),
.Y(n_10356)
);

NAND2xp5_ASAP7_75t_L g10357 ( 
.A(n_9575),
.B(n_497),
.Y(n_10357)
);

AOI22xp5_ASAP7_75t_SL g10358 ( 
.A1(n_9484),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_10358)
);

INVx2_ASAP7_75t_L g10359 ( 
.A(n_9583),
.Y(n_10359)
);

AOI21xp5_ASAP7_75t_L g10360 ( 
.A1(n_9585),
.A2(n_500),
.B(n_501),
.Y(n_10360)
);

BUFx6f_ASAP7_75t_L g10361 ( 
.A(n_9834),
.Y(n_10361)
);

NOR2xp33_ASAP7_75t_L g10362 ( 
.A(n_9300),
.B(n_502),
.Y(n_10362)
);

NAND2xp5_ASAP7_75t_L g10363 ( 
.A(n_9755),
.B(n_503),
.Y(n_10363)
);

NOR2xp33_ASAP7_75t_SL g10364 ( 
.A(n_9413),
.B(n_503),
.Y(n_10364)
);

AOI21xp5_ASAP7_75t_L g10365 ( 
.A1(n_9762),
.A2(n_504),
.B(n_505),
.Y(n_10365)
);

NAND2xp5_ASAP7_75t_L g10366 ( 
.A(n_9763),
.B(n_504),
.Y(n_10366)
);

A2O1A1Ixp33_ASAP7_75t_L g10367 ( 
.A1(n_9587),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_10367)
);

NAND2xp5_ASAP7_75t_L g10368 ( 
.A(n_9802),
.B(n_506),
.Y(n_10368)
);

NAND2xp5_ASAP7_75t_L g10369 ( 
.A(n_9812),
.B(n_507),
.Y(n_10369)
);

AOI21xp5_ASAP7_75t_L g10370 ( 
.A1(n_9814),
.A2(n_508),
.B(n_509),
.Y(n_10370)
);

AOI21xp5_ASAP7_75t_L g10371 ( 
.A1(n_9824),
.A2(n_508),
.B(n_509),
.Y(n_10371)
);

INVx2_ASAP7_75t_L g10372 ( 
.A(n_9829),
.Y(n_10372)
);

NAND2xp5_ASAP7_75t_L g10373 ( 
.A(n_9831),
.B(n_510),
.Y(n_10373)
);

AOI21xp5_ASAP7_75t_L g10374 ( 
.A1(n_9590),
.A2(n_511),
.B(n_512),
.Y(n_10374)
);

AOI21xp5_ASAP7_75t_L g10375 ( 
.A1(n_9737),
.A2(n_512),
.B(n_513),
.Y(n_10375)
);

A2O1A1Ixp33_ASAP7_75t_L g10376 ( 
.A1(n_9323),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_10376)
);

AOI21xp5_ASAP7_75t_L g10377 ( 
.A1(n_9322),
.A2(n_514),
.B(n_516),
.Y(n_10377)
);

NAND2xp5_ASAP7_75t_L g10378 ( 
.A(n_9328),
.B(n_516),
.Y(n_10378)
);

AOI21x1_ASAP7_75t_L g10379 ( 
.A1(n_9355),
.A2(n_9324),
.B(n_9418),
.Y(n_10379)
);

AOI21xp5_ASAP7_75t_L g10380 ( 
.A1(n_9317),
.A2(n_517),
.B(n_518),
.Y(n_10380)
);

NAND2xp5_ASAP7_75t_L g10381 ( 
.A(n_9354),
.B(n_517),
.Y(n_10381)
);

AOI21xp5_ASAP7_75t_L g10382 ( 
.A1(n_9406),
.A2(n_518),
.B(n_519),
.Y(n_10382)
);

INVx2_ASAP7_75t_L g10383 ( 
.A(n_9360),
.Y(n_10383)
);

AND2x2_ASAP7_75t_L g10384 ( 
.A(n_9403),
.B(n_519),
.Y(n_10384)
);

AO21x1_ASAP7_75t_L g10385 ( 
.A1(n_9498),
.A2(n_9270),
.B(n_9405),
.Y(n_10385)
);

OAI22xp5_ASAP7_75t_L g10386 ( 
.A1(n_9396),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_10386)
);

AOI21xp5_ASAP7_75t_L g10387 ( 
.A1(n_9258),
.A2(n_521),
.B(n_523),
.Y(n_10387)
);

AND2x2_ASAP7_75t_L g10388 ( 
.A(n_9272),
.B(n_523),
.Y(n_10388)
);

NAND2xp5_ASAP7_75t_L g10389 ( 
.A(n_9254),
.B(n_524),
.Y(n_10389)
);

AOI22xp5_ASAP7_75t_L g10390 ( 
.A1(n_9258),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_10390)
);

AO32x1_ASAP7_75t_L g10391 ( 
.A1(n_9285),
.A2(n_528),
.A3(n_526),
.B1(n_527),
.B2(n_529),
.Y(n_10391)
);

NAND2xp5_ASAP7_75t_L g10392 ( 
.A(n_9254),
.B(n_528),
.Y(n_10392)
);

AOI21x1_ASAP7_75t_L g10393 ( 
.A1(n_9347),
.A2(n_530),
.B(n_531),
.Y(n_10393)
);

INVx1_ASAP7_75t_L g10394 ( 
.A(n_9286),
.Y(n_10394)
);

A2O1A1Ixp33_ASAP7_75t_L g10395 ( 
.A1(n_9258),
.A2(n_532),
.B(n_530),
.C(n_531),
.Y(n_10395)
);

AOI21x1_ASAP7_75t_L g10396 ( 
.A1(n_9347),
.A2(n_532),
.B(n_533),
.Y(n_10396)
);

INVx2_ASAP7_75t_SL g10397 ( 
.A(n_9307),
.Y(n_10397)
);

HB1xp67_ASAP7_75t_L g10398 ( 
.A(n_9242),
.Y(n_10398)
);

INVx2_ASAP7_75t_L g10399 ( 
.A(n_9241),
.Y(n_10399)
);

AO32x2_ASAP7_75t_L g10400 ( 
.A1(n_9545),
.A2(n_535),
.A3(n_533),
.B1(n_534),
.B2(n_536),
.Y(n_10400)
);

AOI21x1_ASAP7_75t_L g10401 ( 
.A1(n_9347),
.A2(n_535),
.B(n_536),
.Y(n_10401)
);

NAND2xp5_ASAP7_75t_SL g10402 ( 
.A(n_9258),
.B(n_538),
.Y(n_10402)
);

OAI22xp5_ASAP7_75t_L g10403 ( 
.A1(n_9732),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.Y(n_10403)
);

OAI22xp5_ASAP7_75t_L g10404 ( 
.A1(n_9732),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_10404)
);

AND2x4_ASAP7_75t_L g10405 ( 
.A(n_9261),
.B(n_542),
.Y(n_10405)
);

NAND2xp5_ASAP7_75t_L g10406 ( 
.A(n_9254),
.B(n_543),
.Y(n_10406)
);

INVx1_ASAP7_75t_L g10407 ( 
.A(n_9286),
.Y(n_10407)
);

AOI22xp33_ASAP7_75t_SL g10408 ( 
.A1(n_9404),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_10408)
);

AOI21xp5_ASAP7_75t_L g10409 ( 
.A1(n_9258),
.A2(n_544),
.B(n_545),
.Y(n_10409)
);

O2A1O1Ixp5_ASAP7_75t_L g10410 ( 
.A1(n_9258),
.A2(n_548),
.B(n_546),
.C(n_547),
.Y(n_10410)
);

NOR2x1p5_ASAP7_75t_SL g10411 ( 
.A(n_9652),
.B(n_546),
.Y(n_10411)
);

O2A1O1Ixp33_ASAP7_75t_L g10412 ( 
.A1(n_9258),
.A2(n_550),
.B(n_547),
.C(n_549),
.Y(n_10412)
);

BUFx3_ASAP7_75t_L g10413 ( 
.A(n_9287),
.Y(n_10413)
);

NAND2xp5_ASAP7_75t_L g10414 ( 
.A(n_9254),
.B(n_549),
.Y(n_10414)
);

A2O1A1Ixp33_ASAP7_75t_L g10415 ( 
.A1(n_9258),
.A2(n_554),
.B(n_551),
.C(n_552),
.Y(n_10415)
);

INVx2_ASAP7_75t_L g10416 ( 
.A(n_9241),
.Y(n_10416)
);

AOI21xp5_ASAP7_75t_L g10417 ( 
.A1(n_9258),
.A2(n_552),
.B(n_555),
.Y(n_10417)
);

HB1xp67_ASAP7_75t_L g10418 ( 
.A(n_9242),
.Y(n_10418)
);

OAI22x1_ASAP7_75t_L g10419 ( 
.A1(n_9285),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_10419)
);

OR2x6_ASAP7_75t_L g10420 ( 
.A(n_9309),
.B(n_558),
.Y(n_10420)
);

AOI22xp33_ASAP7_75t_L g10421 ( 
.A1(n_9404),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.Y(n_10421)
);

NAND2x1p5_ASAP7_75t_L g10422 ( 
.A(n_9749),
.B(n_561),
.Y(n_10422)
);

NOR2xp33_ASAP7_75t_L g10423 ( 
.A(n_9258),
.B(n_562),
.Y(n_10423)
);

AOI22xp5_ASAP7_75t_L g10424 ( 
.A1(n_9258),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_10424)
);

OAI22xp5_ASAP7_75t_L g10425 ( 
.A1(n_9732),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_10425)
);

NAND2xp5_ASAP7_75t_SL g10426 ( 
.A(n_9258),
.B(n_566),
.Y(n_10426)
);

BUFx4f_ASAP7_75t_L g10427 ( 
.A(n_9784),
.Y(n_10427)
);

NAND2xp5_ASAP7_75t_L g10428 ( 
.A(n_9254),
.B(n_566),
.Y(n_10428)
);

A2O1A1Ixp33_ASAP7_75t_L g10429 ( 
.A1(n_9258),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_10429)
);

AOI21xp5_ASAP7_75t_L g10430 ( 
.A1(n_9258),
.A2(n_567),
.B(n_568),
.Y(n_10430)
);

A2O1A1Ixp33_ASAP7_75t_L g10431 ( 
.A1(n_9258),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_10431)
);

BUFx2_ASAP7_75t_L g10432 ( 
.A(n_9801),
.Y(n_10432)
);

INVx3_ASAP7_75t_L g10433 ( 
.A(n_9761),
.Y(n_10433)
);

AND2x2_ASAP7_75t_L g10434 ( 
.A(n_9272),
.B(n_570),
.Y(n_10434)
);

NOR3xp33_ASAP7_75t_L g10435 ( 
.A(n_9258),
.B(n_571),
.C(n_572),
.Y(n_10435)
);

INVx2_ASAP7_75t_L g10436 ( 
.A(n_9241),
.Y(n_10436)
);

BUFx4f_ASAP7_75t_SL g10437 ( 
.A(n_9341),
.Y(n_10437)
);

OAI22xp5_ASAP7_75t_L g10438 ( 
.A1(n_9732),
.A2(n_576),
.B1(n_573),
.B2(n_574),
.Y(n_10438)
);

NAND2xp5_ASAP7_75t_L g10439 ( 
.A(n_9254),
.B(n_573),
.Y(n_10439)
);

BUFx4f_ASAP7_75t_L g10440 ( 
.A(n_9784),
.Y(n_10440)
);

INVx2_ASAP7_75t_L g10441 ( 
.A(n_9241),
.Y(n_10441)
);

NAND2xp5_ASAP7_75t_SL g10442 ( 
.A(n_9258),
.B(n_576),
.Y(n_10442)
);

AOI21xp5_ASAP7_75t_L g10443 ( 
.A1(n_9258),
.A2(n_577),
.B(n_578),
.Y(n_10443)
);

OA21x2_ASAP7_75t_L g10444 ( 
.A1(n_9465),
.A2(n_577),
.B(n_578),
.Y(n_10444)
);

AOI21xp5_ASAP7_75t_L g10445 ( 
.A1(n_9258),
.A2(n_579),
.B(n_580),
.Y(n_10445)
);

INVx1_ASAP7_75t_L g10446 ( 
.A(n_9286),
.Y(n_10446)
);

NAND2xp5_ASAP7_75t_L g10447 ( 
.A(n_9254),
.B(n_579),
.Y(n_10447)
);

AO31x2_ASAP7_75t_L g10448 ( 
.A1(n_9652),
.A2(n_583),
.A3(n_581),
.B(n_582),
.Y(n_10448)
);

OAI22xp5_ASAP7_75t_L g10449 ( 
.A1(n_9732),
.A2(n_584),
.B1(n_581),
.B2(n_583),
.Y(n_10449)
);

NAND2xp5_ASAP7_75t_L g10450 ( 
.A(n_9254),
.B(n_584),
.Y(n_10450)
);

NAND2xp5_ASAP7_75t_L g10451 ( 
.A(n_9254),
.B(n_585),
.Y(n_10451)
);

NOR2xp67_ASAP7_75t_L g10452 ( 
.A(n_9430),
.B(n_585),
.Y(n_10452)
);

AOI21xp5_ASAP7_75t_L g10453 ( 
.A1(n_9258),
.A2(n_586),
.B(n_587),
.Y(n_10453)
);

INVx2_ASAP7_75t_L g10454 ( 
.A(n_9241),
.Y(n_10454)
);

BUFx6f_ASAP7_75t_L g10455 ( 
.A(n_9784),
.Y(n_10455)
);

AOI21xp5_ASAP7_75t_L g10456 ( 
.A1(n_9258),
.A2(n_587),
.B(n_588),
.Y(n_10456)
);

INVx3_ASAP7_75t_L g10457 ( 
.A(n_9761),
.Y(n_10457)
);

BUFx4f_ASAP7_75t_SL g10458 ( 
.A(n_9341),
.Y(n_10458)
);

AOI21x1_ASAP7_75t_L g10459 ( 
.A1(n_9347),
.A2(n_588),
.B(n_589),
.Y(n_10459)
);

AOI22xp5_ASAP7_75t_L g10460 ( 
.A1(n_9258),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_10460)
);

AOI21xp5_ASAP7_75t_L g10461 ( 
.A1(n_9258),
.A2(n_590),
.B(n_591),
.Y(n_10461)
);

NAND2xp5_ASAP7_75t_SL g10462 ( 
.A(n_9258),
.B(n_592),
.Y(n_10462)
);

NAND2xp5_ASAP7_75t_L g10463 ( 
.A(n_9254),
.B(n_593),
.Y(n_10463)
);

NAND2xp5_ASAP7_75t_L g10464 ( 
.A(n_9254),
.B(n_593),
.Y(n_10464)
);

OAI22xp5_ASAP7_75t_L g10465 ( 
.A1(n_9732),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.Y(n_10465)
);

NAND2xp5_ASAP7_75t_SL g10466 ( 
.A(n_9258),
.B(n_594),
.Y(n_10466)
);

INVxp67_ASAP7_75t_L g10467 ( 
.A(n_9319),
.Y(n_10467)
);

O2A1O1Ixp33_ASAP7_75t_SL g10468 ( 
.A1(n_9258),
.A2(n_597),
.B(n_595),
.C(n_596),
.Y(n_10468)
);

NAND2xp5_ASAP7_75t_L g10469 ( 
.A(n_9254),
.B(n_597),
.Y(n_10469)
);

AOI21xp5_ASAP7_75t_L g10470 ( 
.A1(n_9258),
.A2(n_598),
.B(n_599),
.Y(n_10470)
);

INVxp67_ASAP7_75t_L g10471 ( 
.A(n_9319),
.Y(n_10471)
);

AOI21xp5_ASAP7_75t_L g10472 ( 
.A1(n_9258),
.A2(n_598),
.B(n_599),
.Y(n_10472)
);

NAND2xp5_ASAP7_75t_L g10473 ( 
.A(n_9254),
.B(n_600),
.Y(n_10473)
);

INVx1_ASAP7_75t_L g10474 ( 
.A(n_9286),
.Y(n_10474)
);

AOI21xp5_ASAP7_75t_L g10475 ( 
.A1(n_9258),
.A2(n_600),
.B(n_601),
.Y(n_10475)
);

NOR2xp33_ASAP7_75t_L g10476 ( 
.A(n_9258),
.B(n_601),
.Y(n_10476)
);

INVxp67_ASAP7_75t_L g10477 ( 
.A(n_9319),
.Y(n_10477)
);

AND2x2_ASAP7_75t_L g10478 ( 
.A(n_9272),
.B(n_602),
.Y(n_10478)
);

O2A1O1Ixp33_ASAP7_75t_L g10479 ( 
.A1(n_9258),
.A2(n_604),
.B(n_602),
.C(n_603),
.Y(n_10479)
);

AOI21xp5_ASAP7_75t_L g10480 ( 
.A1(n_9258),
.A2(n_603),
.B(n_605),
.Y(n_10480)
);

AOI21xp5_ASAP7_75t_L g10481 ( 
.A1(n_9258),
.A2(n_605),
.B(n_606),
.Y(n_10481)
);

AOI33xp33_ASAP7_75t_L g10482 ( 
.A1(n_9508),
.A2(n_608),
.A3(n_610),
.B1(n_606),
.B2(n_607),
.B3(n_609),
.Y(n_10482)
);

AOI21xp5_ASAP7_75t_L g10483 ( 
.A1(n_9258),
.A2(n_607),
.B(n_609),
.Y(n_10483)
);

BUFx6f_ASAP7_75t_L g10484 ( 
.A(n_9784),
.Y(n_10484)
);

AOI21xp5_ASAP7_75t_L g10485 ( 
.A1(n_9258),
.A2(n_610),
.B(n_611),
.Y(n_10485)
);

NAND2xp5_ASAP7_75t_L g10486 ( 
.A(n_9254),
.B(n_611),
.Y(n_10486)
);

HB1xp67_ASAP7_75t_L g10487 ( 
.A(n_9242),
.Y(n_10487)
);

AOI21xp5_ASAP7_75t_L g10488 ( 
.A1(n_9258),
.A2(n_612),
.B(n_613),
.Y(n_10488)
);

NAND2xp5_ASAP7_75t_L g10489 ( 
.A(n_9254),
.B(n_612),
.Y(n_10489)
);

NAND2xp5_ASAP7_75t_L g10490 ( 
.A(n_9254),
.B(n_613),
.Y(n_10490)
);

INVx2_ASAP7_75t_L g10491 ( 
.A(n_9241),
.Y(n_10491)
);

NAND2xp5_ASAP7_75t_SL g10492 ( 
.A(n_9258),
.B(n_614),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_9286),
.Y(n_10493)
);

AOI21xp5_ASAP7_75t_L g10494 ( 
.A1(n_9258),
.A2(n_614),
.B(n_615),
.Y(n_10494)
);

INVx1_ASAP7_75t_L g10495 ( 
.A(n_9286),
.Y(n_10495)
);

AOI21xp5_ASAP7_75t_L g10496 ( 
.A1(n_9258),
.A2(n_615),
.B(n_616),
.Y(n_10496)
);

AOI21xp5_ASAP7_75t_L g10497 ( 
.A1(n_9258),
.A2(n_616),
.B(n_617),
.Y(n_10497)
);

INVx1_ASAP7_75t_L g10498 ( 
.A(n_9286),
.Y(n_10498)
);

O2A1O1Ixp33_ASAP7_75t_L g10499 ( 
.A1(n_9258),
.A2(n_619),
.B(n_617),
.C(n_618),
.Y(n_10499)
);

NOR3xp33_ASAP7_75t_L g10500 ( 
.A(n_9258),
.B(n_619),
.C(n_620),
.Y(n_10500)
);

NAND2xp5_ASAP7_75t_L g10501 ( 
.A(n_9254),
.B(n_620),
.Y(n_10501)
);

OAI21xp5_ASAP7_75t_L g10502 ( 
.A1(n_9258),
.A2(n_621),
.B(n_622),
.Y(n_10502)
);

OAI22xp5_ASAP7_75t_L g10503 ( 
.A1(n_9732),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_10503)
);

INVx2_ASAP7_75t_L g10504 ( 
.A(n_9241),
.Y(n_10504)
);

AOI21xp5_ASAP7_75t_L g10505 ( 
.A1(n_9258),
.A2(n_624),
.B(n_625),
.Y(n_10505)
);

BUFx2_ASAP7_75t_L g10506 ( 
.A(n_9801),
.Y(n_10506)
);

INVx2_ASAP7_75t_L g10507 ( 
.A(n_9241),
.Y(n_10507)
);

NAND2x1p5_ASAP7_75t_L g10508 ( 
.A(n_9749),
.B(n_625),
.Y(n_10508)
);

OAI22xp5_ASAP7_75t_L g10509 ( 
.A1(n_9732),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_10509)
);

AOI21xp5_ASAP7_75t_L g10510 ( 
.A1(n_9258),
.A2(n_626),
.B(n_628),
.Y(n_10510)
);

NOR2xp33_ASAP7_75t_L g10511 ( 
.A(n_9258),
.B(n_629),
.Y(n_10511)
);

A2O1A1Ixp33_ASAP7_75t_L g10512 ( 
.A1(n_9258),
.A2(n_631),
.B(n_629),
.C(n_630),
.Y(n_10512)
);

AND2x2_ASAP7_75t_L g10513 ( 
.A(n_9272),
.B(n_630),
.Y(n_10513)
);

INVx2_ASAP7_75t_L g10514 ( 
.A(n_9241),
.Y(n_10514)
);

A2O1A1Ixp33_ASAP7_75t_L g10515 ( 
.A1(n_9258),
.A2(n_635),
.B(n_631),
.C(n_633),
.Y(n_10515)
);

BUFx6f_ASAP7_75t_L g10516 ( 
.A(n_9784),
.Y(n_10516)
);

INVx2_ASAP7_75t_L g10517 ( 
.A(n_9241),
.Y(n_10517)
);

NAND2xp5_ASAP7_75t_SL g10518 ( 
.A(n_9258),
.B(n_633),
.Y(n_10518)
);

HB1xp67_ASAP7_75t_L g10519 ( 
.A(n_9242),
.Y(n_10519)
);

AOI21xp5_ASAP7_75t_L g10520 ( 
.A1(n_9258),
.A2(n_635),
.B(n_636),
.Y(n_10520)
);

AOI21xp5_ASAP7_75t_L g10521 ( 
.A1(n_9258),
.A2(n_637),
.B(n_638),
.Y(n_10521)
);

INVx1_ASAP7_75t_L g10522 ( 
.A(n_9286),
.Y(n_10522)
);

INVx1_ASAP7_75t_L g10523 ( 
.A(n_9286),
.Y(n_10523)
);

INVx1_ASAP7_75t_L g10524 ( 
.A(n_9286),
.Y(n_10524)
);

AOI21x1_ASAP7_75t_L g10525 ( 
.A1(n_9347),
.A2(n_637),
.B(n_639),
.Y(n_10525)
);

NAND2xp5_ASAP7_75t_SL g10526 ( 
.A(n_9258),
.B(n_639),
.Y(n_10526)
);

NAND2xp5_ASAP7_75t_L g10527 ( 
.A(n_9254),
.B(n_640),
.Y(n_10527)
);

INVx2_ASAP7_75t_L g10528 ( 
.A(n_9241),
.Y(n_10528)
);

NAND2x1_ASAP7_75t_L g10529 ( 
.A(n_9652),
.B(n_641),
.Y(n_10529)
);

OA22x2_ASAP7_75t_L g10530 ( 
.A1(n_9258),
.A2(n_643),
.B1(n_641),
.B2(n_642),
.Y(n_10530)
);

AOI21xp5_ASAP7_75t_L g10531 ( 
.A1(n_9258),
.A2(n_642),
.B(n_643),
.Y(n_10531)
);

AOI21x1_ASAP7_75t_L g10532 ( 
.A1(n_9347),
.A2(n_644),
.B(n_645),
.Y(n_10532)
);

O2A1O1Ixp33_ASAP7_75t_L g10533 ( 
.A1(n_9258),
.A2(n_646),
.B(n_644),
.C(n_645),
.Y(n_10533)
);

BUFx6f_ASAP7_75t_L g10534 ( 
.A(n_9784),
.Y(n_10534)
);

BUFx2_ASAP7_75t_L g10535 ( 
.A(n_9801),
.Y(n_10535)
);

A2O1A1Ixp33_ASAP7_75t_L g10536 ( 
.A1(n_9258),
.A2(n_648),
.B(n_646),
.C(n_647),
.Y(n_10536)
);

OAI22xp5_ASAP7_75t_L g10537 ( 
.A1(n_9732),
.A2(n_650),
.B1(n_648),
.B2(n_649),
.Y(n_10537)
);

INVx1_ASAP7_75t_L g10538 ( 
.A(n_9286),
.Y(n_10538)
);

NOR2xp67_ASAP7_75t_L g10539 ( 
.A(n_9430),
.B(n_650),
.Y(n_10539)
);

AOI21xp5_ASAP7_75t_L g10540 ( 
.A1(n_9258),
.A2(n_651),
.B(n_652),
.Y(n_10540)
);

NAND2xp5_ASAP7_75t_L g10541 ( 
.A(n_9254),
.B(n_652),
.Y(n_10541)
);

INVx1_ASAP7_75t_L g10542 ( 
.A(n_9286),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_9286),
.Y(n_10543)
);

AOI21xp5_ASAP7_75t_L g10544 ( 
.A1(n_9258),
.A2(n_653),
.B(n_654),
.Y(n_10544)
);

AOI21xp5_ASAP7_75t_L g10545 ( 
.A1(n_9258),
.A2(n_653),
.B(n_654),
.Y(n_10545)
);

INVx1_ASAP7_75t_L g10546 ( 
.A(n_9286),
.Y(n_10546)
);

NAND2xp5_ASAP7_75t_SL g10547 ( 
.A(n_9258),
.B(n_655),
.Y(n_10547)
);

OAI321xp33_ASAP7_75t_L g10548 ( 
.A1(n_9258),
.A2(n_657),
.A3(n_659),
.B1(n_655),
.B2(n_656),
.C(n_658),
.Y(n_10548)
);

HB1xp67_ASAP7_75t_L g10549 ( 
.A(n_9242),
.Y(n_10549)
);

AOI21xp5_ASAP7_75t_L g10550 ( 
.A1(n_9258),
.A2(n_657),
.B(n_658),
.Y(n_10550)
);

A2O1A1Ixp33_ASAP7_75t_L g10551 ( 
.A1(n_9258),
.A2(n_662),
.B(n_660),
.C(n_661),
.Y(n_10551)
);

NOR2xp33_ASAP7_75t_L g10552 ( 
.A(n_9258),
.B(n_660),
.Y(n_10552)
);

NAND2xp5_ASAP7_75t_L g10553 ( 
.A(n_9254),
.B(n_661),
.Y(n_10553)
);

AOI21xp5_ASAP7_75t_L g10554 ( 
.A1(n_9258),
.A2(n_663),
.B(n_664),
.Y(n_10554)
);

NOR2xp33_ASAP7_75t_L g10555 ( 
.A(n_9258),
.B(n_664),
.Y(n_10555)
);

AO22x1_ASAP7_75t_L g10556 ( 
.A1(n_9258),
.A2(n_667),
.B1(n_665),
.B2(n_666),
.Y(n_10556)
);

INVx4_ASAP7_75t_L g10557 ( 
.A(n_9749),
.Y(n_10557)
);

INVx1_ASAP7_75t_L g10558 ( 
.A(n_9286),
.Y(n_10558)
);

A2O1A1Ixp33_ASAP7_75t_L g10559 ( 
.A1(n_9258),
.A2(n_669),
.B(n_667),
.C(n_668),
.Y(n_10559)
);

AOI21xp5_ASAP7_75t_L g10560 ( 
.A1(n_9258),
.A2(n_668),
.B(n_669),
.Y(n_10560)
);

AOI21xp5_ASAP7_75t_L g10561 ( 
.A1(n_9258),
.A2(n_670),
.B(n_671),
.Y(n_10561)
);

INVx3_ASAP7_75t_L g10562 ( 
.A(n_9761),
.Y(n_10562)
);

BUFx3_ASAP7_75t_L g10563 ( 
.A(n_9287),
.Y(n_10563)
);

AOI22xp5_ASAP7_75t_L g10564 ( 
.A1(n_9258),
.A2(n_673),
.B1(n_671),
.B2(n_672),
.Y(n_10564)
);

OAI22xp5_ASAP7_75t_L g10565 ( 
.A1(n_10423),
.A2(n_674),
.B1(n_672),
.B2(n_673),
.Y(n_10565)
);

O2A1O1Ixp33_ASAP7_75t_L g10566 ( 
.A1(n_9966),
.A2(n_9883),
.B(n_10511),
.C(n_10476),
.Y(n_10566)
);

AND2x4_ASAP7_75t_L g10567 ( 
.A(n_10252),
.B(n_674),
.Y(n_10567)
);

AOI22xp33_ASAP7_75t_L g10568 ( 
.A1(n_9950),
.A2(n_677),
.B1(n_675),
.B2(n_676),
.Y(n_10568)
);

INVx1_ASAP7_75t_L g10569 ( 
.A(n_10010),
.Y(n_10569)
);

AOI21x1_ASAP7_75t_L g10570 ( 
.A1(n_10078),
.A2(n_675),
.B(n_676),
.Y(n_10570)
);

INVx2_ASAP7_75t_L g10571 ( 
.A(n_10235),
.Y(n_10571)
);

INVx1_ASAP7_75t_SL g10572 ( 
.A(n_10230),
.Y(n_10572)
);

AND2x4_ASAP7_75t_L g10573 ( 
.A(n_10432),
.B(n_677),
.Y(n_10573)
);

BUFx6f_ASAP7_75t_L g10574 ( 
.A(n_10114),
.Y(n_10574)
);

AOI21xp5_ASAP7_75t_L g10575 ( 
.A1(n_9912),
.A2(n_678),
.B(n_679),
.Y(n_10575)
);

OAI22x1_ASAP7_75t_L g10576 ( 
.A1(n_9887),
.A2(n_680),
.B1(n_678),
.B2(n_679),
.Y(n_10576)
);

NAND2xp5_ASAP7_75t_L g10577 ( 
.A(n_10506),
.B(n_680),
.Y(n_10577)
);

NAND2xp5_ASAP7_75t_L g10578 ( 
.A(n_10535),
.B(n_9882),
.Y(n_10578)
);

A2O1A1Ixp33_ASAP7_75t_L g10579 ( 
.A1(n_9879),
.A2(n_683),
.B(n_681),
.C(n_682),
.Y(n_10579)
);

OAI22xp5_ASAP7_75t_L g10580 ( 
.A1(n_10552),
.A2(n_683),
.B1(n_681),
.B2(n_682),
.Y(n_10580)
);

INVx2_ASAP7_75t_L g10581 ( 
.A(n_10283),
.Y(n_10581)
);

AOI21xp5_ASAP7_75t_L g10582 ( 
.A1(n_9843),
.A2(n_684),
.B(n_686),
.Y(n_10582)
);

AOI22xp33_ASAP7_75t_L g10583 ( 
.A1(n_9844),
.A2(n_688),
.B1(n_684),
.B2(n_687),
.Y(n_10583)
);

A2O1A1Ixp33_ASAP7_75t_SL g10584 ( 
.A1(n_10555),
.A2(n_690),
.B(n_688),
.C(n_689),
.Y(n_10584)
);

OR2x6_ASAP7_75t_L g10585 ( 
.A(n_10219),
.B(n_689),
.Y(n_10585)
);

AOI21xp5_ASAP7_75t_L g10586 ( 
.A1(n_9897),
.A2(n_9840),
.B(n_9949),
.Y(n_10586)
);

INVx1_ASAP7_75t_L g10587 ( 
.A(n_9982),
.Y(n_10587)
);

BUFx3_ASAP7_75t_L g10588 ( 
.A(n_10057),
.Y(n_10588)
);

INVx2_ASAP7_75t_SL g10589 ( 
.A(n_10281),
.Y(n_10589)
);

NOR2xp33_ASAP7_75t_L g10590 ( 
.A(n_10281),
.B(n_690),
.Y(n_10590)
);

INVx2_ASAP7_75t_SL g10591 ( 
.A(n_10274),
.Y(n_10591)
);

INVx2_ASAP7_75t_SL g10592 ( 
.A(n_9980),
.Y(n_10592)
);

NAND2xp33_ASAP7_75t_SL g10593 ( 
.A(n_10260),
.B(n_10482),
.Y(n_10593)
);

NAND2xp5_ASAP7_75t_L g10594 ( 
.A(n_9924),
.B(n_691),
.Y(n_10594)
);

BUFx6f_ASAP7_75t_L g10595 ( 
.A(n_10114),
.Y(n_10595)
);

NAND2xp5_ASAP7_75t_SL g10596 ( 
.A(n_10024),
.B(n_691),
.Y(n_10596)
);

AOI21xp5_ASAP7_75t_L g10597 ( 
.A1(n_10502),
.A2(n_692),
.B(n_693),
.Y(n_10597)
);

AOI22xp5_ASAP7_75t_L g10598 ( 
.A1(n_9890),
.A2(n_694),
.B1(n_692),
.B2(n_693),
.Y(n_10598)
);

OAI22xp5_ASAP7_75t_SL g10599 ( 
.A1(n_10141),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_10599)
);

NAND2xp5_ASAP7_75t_SL g10600 ( 
.A(n_10059),
.B(n_695),
.Y(n_10600)
);

AND2x6_ASAP7_75t_L g10601 ( 
.A(n_10083),
.B(n_696),
.Y(n_10601)
);

O2A1O1Ixp33_ASAP7_75t_L g10602 ( 
.A1(n_9917),
.A2(n_10435),
.B(n_10500),
.C(n_9931),
.Y(n_10602)
);

BUFx3_ASAP7_75t_L g10603 ( 
.A(n_9972),
.Y(n_10603)
);

AOI21xp5_ASAP7_75t_L g10604 ( 
.A1(n_9914),
.A2(n_697),
.B(n_698),
.Y(n_10604)
);

NAND2xp5_ASAP7_75t_L g10605 ( 
.A(n_10398),
.B(n_698),
.Y(n_10605)
);

NAND3xp33_ASAP7_75t_L g10606 ( 
.A(n_9979),
.B(n_699),
.C(n_700),
.Y(n_10606)
);

NAND2xp5_ASAP7_75t_L g10607 ( 
.A(n_10418),
.B(n_699),
.Y(n_10607)
);

AOI21x1_ASAP7_75t_L g10608 ( 
.A1(n_9908),
.A2(n_9869),
.B(n_9932),
.Y(n_10608)
);

BUFx3_ASAP7_75t_L g10609 ( 
.A(n_10413),
.Y(n_10609)
);

CKINVDCx5p33_ASAP7_75t_R g10610 ( 
.A(n_10051),
.Y(n_10610)
);

AOI21xp5_ASAP7_75t_L g10611 ( 
.A1(n_10548),
.A2(n_700),
.B(n_701),
.Y(n_10611)
);

BUFx12f_ASAP7_75t_L g10612 ( 
.A(n_10160),
.Y(n_10612)
);

NOR2xp33_ASAP7_75t_R g10613 ( 
.A(n_10437),
.B(n_702),
.Y(n_10613)
);

NOR2xp67_ASAP7_75t_L g10614 ( 
.A(n_10487),
.B(n_702),
.Y(n_10614)
);

HB1xp67_ASAP7_75t_L g10615 ( 
.A(n_9990),
.Y(n_10615)
);

INVx4_ASAP7_75t_L g10616 ( 
.A(n_10205),
.Y(n_10616)
);

OR2x2_ASAP7_75t_L g10617 ( 
.A(n_10519),
.B(n_703),
.Y(n_10617)
);

BUFx3_ASAP7_75t_L g10618 ( 
.A(n_10563),
.Y(n_10618)
);

A2O1A1Ixp33_ASAP7_75t_SL g10619 ( 
.A1(n_10409),
.A2(n_706),
.B(n_704),
.C(n_705),
.Y(n_10619)
);

CKINVDCx5p33_ASAP7_75t_R g10620 ( 
.A(n_10087),
.Y(n_10620)
);

NAND2xp5_ASAP7_75t_L g10621 ( 
.A(n_10549),
.B(n_704),
.Y(n_10621)
);

NAND2xp5_ASAP7_75t_L g10622 ( 
.A(n_9954),
.B(n_705),
.Y(n_10622)
);

OAI21xp5_ASAP7_75t_L g10623 ( 
.A1(n_9839),
.A2(n_706),
.B(n_707),
.Y(n_10623)
);

NAND2xp5_ASAP7_75t_SL g10624 ( 
.A(n_10284),
.B(n_707),
.Y(n_10624)
);

NOR2xp33_ASAP7_75t_L g10625 ( 
.A(n_10173),
.B(n_708),
.Y(n_10625)
);

O2A1O1Ixp33_ASAP7_75t_L g10626 ( 
.A1(n_10046),
.A2(n_711),
.B(n_709),
.C(n_710),
.Y(n_10626)
);

HB1xp67_ASAP7_75t_L g10627 ( 
.A(n_10262),
.Y(n_10627)
);

INVx5_ASAP7_75t_L g10628 ( 
.A(n_10420),
.Y(n_10628)
);

BUFx6f_ASAP7_75t_L g10629 ( 
.A(n_9980),
.Y(n_10629)
);

BUFx3_ASAP7_75t_L g10630 ( 
.A(n_10229),
.Y(n_10630)
);

A2O1A1Ixp33_ASAP7_75t_L g10631 ( 
.A1(n_9922),
.A2(n_711),
.B(n_709),
.C(n_710),
.Y(n_10631)
);

NOR2xp33_ASAP7_75t_L g10632 ( 
.A(n_10201),
.B(n_712),
.Y(n_10632)
);

NOR2xp33_ASAP7_75t_R g10633 ( 
.A(n_10458),
.B(n_9995),
.Y(n_10633)
);

NAND2xp5_ASAP7_75t_L g10634 ( 
.A(n_10004),
.B(n_712),
.Y(n_10634)
);

INVx2_ASAP7_75t_L g10635 ( 
.A(n_10287),
.Y(n_10635)
);

INVx2_ASAP7_75t_L g10636 ( 
.A(n_10314),
.Y(n_10636)
);

NAND2xp5_ASAP7_75t_L g10637 ( 
.A(n_9872),
.B(n_713),
.Y(n_10637)
);

AOI21xp5_ASAP7_75t_L g10638 ( 
.A1(n_9893),
.A2(n_10479),
.B(n_10412),
.Y(n_10638)
);

A2O1A1Ixp33_ASAP7_75t_SL g10639 ( 
.A1(n_10430),
.A2(n_715),
.B(n_713),
.C(n_714),
.Y(n_10639)
);

NOR2xp33_ASAP7_75t_L g10640 ( 
.A(n_10041),
.B(n_714),
.Y(n_10640)
);

AND2x4_ASAP7_75t_L g10641 ( 
.A(n_10196),
.B(n_716),
.Y(n_10641)
);

INVx2_ASAP7_75t_L g10642 ( 
.A(n_10318),
.Y(n_10642)
);

NAND2xp5_ASAP7_75t_SL g10643 ( 
.A(n_9988),
.B(n_716),
.Y(n_10643)
);

OAI21xp5_ASAP7_75t_L g10644 ( 
.A1(n_10387),
.A2(n_10443),
.B(n_10417),
.Y(n_10644)
);

A2O1A1Ixp33_ASAP7_75t_L g10645 ( 
.A1(n_9863),
.A2(n_719),
.B(n_717),
.C(n_718),
.Y(n_10645)
);

AOI21xp5_ASAP7_75t_L g10646 ( 
.A1(n_10499),
.A2(n_718),
.B(n_719),
.Y(n_10646)
);

AO21x1_ASAP7_75t_L g10647 ( 
.A1(n_10084),
.A2(n_720),
.B(n_722),
.Y(n_10647)
);

AOI21xp5_ASAP7_75t_L g10648 ( 
.A1(n_10533),
.A2(n_720),
.B(n_722),
.Y(n_10648)
);

INVx1_ASAP7_75t_L g10649 ( 
.A(n_10558),
.Y(n_10649)
);

AND2x6_ASAP7_75t_L g10650 ( 
.A(n_10179),
.B(n_723),
.Y(n_10650)
);

INVx2_ASAP7_75t_SL g10651 ( 
.A(n_10351),
.Y(n_10651)
);

INVx5_ASAP7_75t_L g10652 ( 
.A(n_10420),
.Y(n_10652)
);

NOR2xp33_ASAP7_75t_L g10653 ( 
.A(n_10063),
.B(n_723),
.Y(n_10653)
);

INVxp67_ASAP7_75t_L g10654 ( 
.A(n_9958),
.Y(n_10654)
);

INVx1_ASAP7_75t_L g10655 ( 
.A(n_9895),
.Y(n_10655)
);

AOI21xp5_ASAP7_75t_L g10656 ( 
.A1(n_10402),
.A2(n_724),
.B(n_725),
.Y(n_10656)
);

AOI21xp5_ASAP7_75t_L g10657 ( 
.A1(n_10426),
.A2(n_724),
.B(n_725),
.Y(n_10657)
);

AND2x4_ASAP7_75t_L g10658 ( 
.A(n_10249),
.B(n_726),
.Y(n_10658)
);

OAI22xp5_ASAP7_75t_L g10659 ( 
.A1(n_10132),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_10659)
);

INVx3_ASAP7_75t_L g10660 ( 
.A(n_9910),
.Y(n_10660)
);

NAND2xp5_ASAP7_75t_SL g10661 ( 
.A(n_10214),
.B(n_728),
.Y(n_10661)
);

NOR2xp33_ASAP7_75t_R g10662 ( 
.A(n_10243),
.B(n_729),
.Y(n_10662)
);

NOR2xp33_ASAP7_75t_L g10663 ( 
.A(n_10212),
.B(n_729),
.Y(n_10663)
);

AOI21xp5_ASAP7_75t_L g10664 ( 
.A1(n_10442),
.A2(n_730),
.B(n_731),
.Y(n_10664)
);

OAI22xp5_ASAP7_75t_L g10665 ( 
.A1(n_10192),
.A2(n_733),
.B1(n_730),
.B2(n_732),
.Y(n_10665)
);

INVx2_ASAP7_75t_L g10666 ( 
.A(n_10331),
.Y(n_10666)
);

BUFx3_ASAP7_75t_L g10667 ( 
.A(n_10229),
.Y(n_10667)
);

NAND2xp5_ASAP7_75t_L g10668 ( 
.A(n_9921),
.B(n_732),
.Y(n_10668)
);

CKINVDCx20_ASAP7_75t_R g10669 ( 
.A(n_9838),
.Y(n_10669)
);

AOI21xp5_ASAP7_75t_L g10670 ( 
.A1(n_10462),
.A2(n_734),
.B(n_735),
.Y(n_10670)
);

NAND2x1p5_ASAP7_75t_L g10671 ( 
.A(n_10350),
.B(n_9853),
.Y(n_10671)
);

O2A1O1Ixp33_ASAP7_75t_L g10672 ( 
.A1(n_10466),
.A2(n_737),
.B(n_734),
.C(n_736),
.Y(n_10672)
);

AOI21xp5_ASAP7_75t_L g10673 ( 
.A1(n_10492),
.A2(n_737),
.B(n_738),
.Y(n_10673)
);

NAND2xp5_ASAP7_75t_L g10674 ( 
.A(n_9947),
.B(n_738),
.Y(n_10674)
);

NAND3xp33_ASAP7_75t_SL g10675 ( 
.A(n_10035),
.B(n_740),
.C(n_742),
.Y(n_10675)
);

O2A1O1Ixp5_ASAP7_75t_L g10676 ( 
.A1(n_10556),
.A2(n_743),
.B(n_740),
.C(n_742),
.Y(n_10676)
);

O2A1O1Ixp33_ASAP7_75t_L g10677 ( 
.A1(n_10518),
.A2(n_746),
.B(n_744),
.C(n_745),
.Y(n_10677)
);

INVx3_ASAP7_75t_L g10678 ( 
.A(n_9978),
.Y(n_10678)
);

NOR2xp33_ASAP7_75t_L g10679 ( 
.A(n_10323),
.B(n_744),
.Y(n_10679)
);

NAND3xp33_ASAP7_75t_SL g10680 ( 
.A(n_9864),
.B(n_746),
.C(n_747),
.Y(n_10680)
);

INVx3_ASAP7_75t_L g10681 ( 
.A(n_10038),
.Y(n_10681)
);

O2A1O1Ixp33_ASAP7_75t_SL g10682 ( 
.A1(n_10526),
.A2(n_750),
.B(n_747),
.C(n_749),
.Y(n_10682)
);

NAND2xp5_ASAP7_75t_L g10683 ( 
.A(n_9953),
.B(n_749),
.Y(n_10683)
);

NOR3xp33_ASAP7_75t_SL g10684 ( 
.A(n_10547),
.B(n_750),
.C(n_751),
.Y(n_10684)
);

INVx2_ASAP7_75t_L g10685 ( 
.A(n_10145),
.Y(n_10685)
);

OAI22xp5_ASAP7_75t_SL g10686 ( 
.A1(n_10055),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.Y(n_10686)
);

INVx1_ASAP7_75t_L g10687 ( 
.A(n_9971),
.Y(n_10687)
);

OAI22xp5_ASAP7_75t_L g10688 ( 
.A1(n_10317),
.A2(n_755),
.B1(n_752),
.B2(n_754),
.Y(n_10688)
);

INVx4_ASAP7_75t_L g10689 ( 
.A(n_10427),
.Y(n_10689)
);

AND2x2_ASAP7_75t_L g10690 ( 
.A(n_10096),
.B(n_755),
.Y(n_10690)
);

BUFx6f_ASAP7_75t_L g10691 ( 
.A(n_10440),
.Y(n_10691)
);

NAND2xp5_ASAP7_75t_L g10692 ( 
.A(n_9977),
.B(n_10394),
.Y(n_10692)
);

INVx5_ASAP7_75t_L g10693 ( 
.A(n_10557),
.Y(n_10693)
);

AOI22xp5_ASAP7_75t_L g10694 ( 
.A1(n_9929),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.Y(n_10694)
);

AOI21x1_ASAP7_75t_SL g10695 ( 
.A1(n_9962),
.A2(n_9970),
.B(n_9948),
.Y(n_10695)
);

AND2x2_ASAP7_75t_L g10696 ( 
.A(n_10162),
.B(n_756),
.Y(n_10696)
);

NAND2xp5_ASAP7_75t_L g10697 ( 
.A(n_10407),
.B(n_759),
.Y(n_10697)
);

NAND2xp5_ASAP7_75t_SL g10698 ( 
.A(n_10385),
.B(n_759),
.Y(n_10698)
);

OR2x6_ASAP7_75t_L g10699 ( 
.A(n_10242),
.B(n_760),
.Y(n_10699)
);

INVx3_ASAP7_75t_L g10700 ( 
.A(n_10338),
.Y(n_10700)
);

INVx2_ASAP7_75t_L g10701 ( 
.A(n_10165),
.Y(n_10701)
);

INVx5_ASAP7_75t_L g10702 ( 
.A(n_10208),
.Y(n_10702)
);

AOI21xp5_ASAP7_75t_L g10703 ( 
.A1(n_9881),
.A2(n_10138),
.B(n_9876),
.Y(n_10703)
);

INVx2_ASAP7_75t_SL g10704 ( 
.A(n_10139),
.Y(n_10704)
);

INVx4_ASAP7_75t_L g10705 ( 
.A(n_10455),
.Y(n_10705)
);

A2O1A1Ixp33_ASAP7_75t_L g10706 ( 
.A1(n_9874),
.A2(n_762),
.B(n_760),
.C(n_761),
.Y(n_10706)
);

NOR2xp33_ASAP7_75t_L g10707 ( 
.A(n_10323),
.B(n_761),
.Y(n_10707)
);

AND2x2_ASAP7_75t_L g10708 ( 
.A(n_9846),
.B(n_10467),
.Y(n_10708)
);

BUFx4f_ASAP7_75t_L g10709 ( 
.A(n_10136),
.Y(n_10709)
);

NAND2xp33_ASAP7_75t_SL g10710 ( 
.A(n_9973),
.B(n_762),
.Y(n_10710)
);

NOR2xp67_ASAP7_75t_SL g10711 ( 
.A(n_10015),
.B(n_10265),
.Y(n_10711)
);

O2A1O1Ixp33_ASAP7_75t_L g10712 ( 
.A1(n_9875),
.A2(n_765),
.B(n_763),
.C(n_764),
.Y(n_10712)
);

NOR2xp33_ASAP7_75t_L g10713 ( 
.A(n_10341),
.B(n_765),
.Y(n_10713)
);

NAND2xp33_ASAP7_75t_SL g10714 ( 
.A(n_10184),
.B(n_766),
.Y(n_10714)
);

NAND2xp5_ASAP7_75t_L g10715 ( 
.A(n_10446),
.B(n_766),
.Y(n_10715)
);

NAND2xp5_ASAP7_75t_L g10716 ( 
.A(n_10474),
.B(n_768),
.Y(n_10716)
);

BUFx2_ASAP7_75t_L g10717 ( 
.A(n_10188),
.Y(n_10717)
);

O2A1O1Ixp33_ASAP7_75t_SL g10718 ( 
.A1(n_10395),
.A2(n_770),
.B(n_768),
.C(n_769),
.Y(n_10718)
);

NAND2xp5_ASAP7_75t_SL g10719 ( 
.A(n_10058),
.B(n_769),
.Y(n_10719)
);

AOI21xp5_ASAP7_75t_L g10720 ( 
.A1(n_9926),
.A2(n_770),
.B(n_771),
.Y(n_10720)
);

CKINVDCx11_ASAP7_75t_R g10721 ( 
.A(n_10092),
.Y(n_10721)
);

OAI22xp5_ASAP7_75t_L g10722 ( 
.A1(n_10177),
.A2(n_773),
.B1(n_771),
.B2(n_772),
.Y(n_10722)
);

AOI21xp5_ASAP7_75t_L g10723 ( 
.A1(n_9938),
.A2(n_773),
.B(n_774),
.Y(n_10723)
);

BUFx6f_ASAP7_75t_L g10724 ( 
.A(n_10455),
.Y(n_10724)
);

BUFx12f_ASAP7_75t_L g10725 ( 
.A(n_9873),
.Y(n_10725)
);

INVx1_ASAP7_75t_L g10726 ( 
.A(n_10493),
.Y(n_10726)
);

OAI21xp33_ASAP7_75t_SL g10727 ( 
.A1(n_10530),
.A2(n_775),
.B(n_776),
.Y(n_10727)
);

NAND2xp5_ASAP7_75t_L g10728 ( 
.A(n_10495),
.B(n_775),
.Y(n_10728)
);

NAND2xp5_ASAP7_75t_SL g10729 ( 
.A(n_10275),
.B(n_777),
.Y(n_10729)
);

NAND2xp5_ASAP7_75t_SL g10730 ( 
.A(n_10142),
.B(n_777),
.Y(n_10730)
);

NAND3xp33_ASAP7_75t_L g10731 ( 
.A(n_10085),
.B(n_778),
.C(n_779),
.Y(n_10731)
);

NAND2xp5_ASAP7_75t_L g10732 ( 
.A(n_10498),
.B(n_780),
.Y(n_10732)
);

A2O1A1Ixp33_ASAP7_75t_L g10733 ( 
.A1(n_10007),
.A2(n_782),
.B(n_780),
.C(n_781),
.Y(n_10733)
);

O2A1O1Ixp33_ASAP7_75t_L g10734 ( 
.A1(n_10014),
.A2(n_783),
.B(n_781),
.C(n_782),
.Y(n_10734)
);

BUFx2_ASAP7_75t_L g10735 ( 
.A(n_10522),
.Y(n_10735)
);

OR2x2_ASAP7_75t_L g10736 ( 
.A(n_10001),
.B(n_783),
.Y(n_10736)
);

O2A1O1Ixp33_ASAP7_75t_L g10737 ( 
.A1(n_9862),
.A2(n_786),
.B(n_784),
.C(n_785),
.Y(n_10737)
);

NAND2xp5_ASAP7_75t_L g10738 ( 
.A(n_10523),
.B(n_784),
.Y(n_10738)
);

AND2x4_ASAP7_75t_L g10739 ( 
.A(n_10110),
.B(n_785),
.Y(n_10739)
);

NOR2xp33_ASAP7_75t_L g10740 ( 
.A(n_10341),
.B(n_786),
.Y(n_10740)
);

NAND3xp33_ASAP7_75t_L g10741 ( 
.A(n_10445),
.B(n_787),
.C(n_788),
.Y(n_10741)
);

NAND2xp5_ASAP7_75t_SL g10742 ( 
.A(n_10097),
.B(n_787),
.Y(n_10742)
);

AOI21xp5_ASAP7_75t_L g10743 ( 
.A1(n_9946),
.A2(n_788),
.B(n_789),
.Y(n_10743)
);

AOI21xp5_ASAP7_75t_L g10744 ( 
.A1(n_10468),
.A2(n_790),
.B(n_791),
.Y(n_10744)
);

INVx2_ASAP7_75t_SL g10745 ( 
.A(n_10316),
.Y(n_10745)
);

NAND2xp5_ASAP7_75t_L g10746 ( 
.A(n_10524),
.B(n_10538),
.Y(n_10746)
);

NAND2xp5_ASAP7_75t_L g10747 ( 
.A(n_10542),
.B(n_10543),
.Y(n_10747)
);

INVxp67_ASAP7_75t_L g10748 ( 
.A(n_10100),
.Y(n_10748)
);

AOI21xp5_ASAP7_75t_L g10749 ( 
.A1(n_10391),
.A2(n_790),
.B(n_791),
.Y(n_10749)
);

AOI21xp5_ASAP7_75t_L g10750 ( 
.A1(n_10391),
.A2(n_792),
.B(n_793),
.Y(n_10750)
);

AO32x2_ASAP7_75t_L g10751 ( 
.A1(n_10330),
.A2(n_10103),
.A3(n_10070),
.B1(n_10278),
.B2(n_9939),
.Y(n_10751)
);

INVx4_ASAP7_75t_L g10752 ( 
.A(n_10484),
.Y(n_10752)
);

NOR2xp33_ASAP7_75t_R g10753 ( 
.A(n_10237),
.B(n_792),
.Y(n_10753)
);

NOR2xp33_ASAP7_75t_L g10754 ( 
.A(n_9849),
.B(n_793),
.Y(n_10754)
);

BUFx12f_ASAP7_75t_L g10755 ( 
.A(n_9956),
.Y(n_10755)
);

NAND2xp5_ASAP7_75t_SL g10756 ( 
.A(n_10379),
.B(n_794),
.Y(n_10756)
);

AOI21xp5_ASAP7_75t_L g10757 ( 
.A1(n_10105),
.A2(n_794),
.B(n_795),
.Y(n_10757)
);

NAND2xp5_ASAP7_75t_L g10758 ( 
.A(n_10546),
.B(n_796),
.Y(n_10758)
);

BUFx6f_ASAP7_75t_L g10759 ( 
.A(n_10484),
.Y(n_10759)
);

BUFx6f_ASAP7_75t_L g10760 ( 
.A(n_10516),
.Y(n_10760)
);

CKINVDCx5p33_ASAP7_75t_R g10761 ( 
.A(n_10270),
.Y(n_10761)
);

INVx3_ASAP7_75t_L g10762 ( 
.A(n_10338),
.Y(n_10762)
);

AOI21xp5_ASAP7_75t_L g10763 ( 
.A1(n_10453),
.A2(n_796),
.B(n_797),
.Y(n_10763)
);

AOI21xp5_ASAP7_75t_L g10764 ( 
.A1(n_10456),
.A2(n_797),
.B(n_798),
.Y(n_10764)
);

NAND2xp5_ASAP7_75t_L g10765 ( 
.A(n_10471),
.B(n_799),
.Y(n_10765)
);

INVx1_ASAP7_75t_L g10766 ( 
.A(n_10002),
.Y(n_10766)
);

O2A1O1Ixp33_ASAP7_75t_L g10767 ( 
.A1(n_10415),
.A2(n_801),
.B(n_799),
.C(n_800),
.Y(n_10767)
);

OAI22xp5_ASAP7_75t_L g10768 ( 
.A1(n_10390),
.A2(n_802),
.B1(n_800),
.B2(n_801),
.Y(n_10768)
);

NAND2xp5_ASAP7_75t_SL g10769 ( 
.A(n_10338),
.B(n_802),
.Y(n_10769)
);

NAND2xp5_ASAP7_75t_L g10770 ( 
.A(n_10477),
.B(n_803),
.Y(n_10770)
);

NAND2xp5_ASAP7_75t_L g10771 ( 
.A(n_10005),
.B(n_803),
.Y(n_10771)
);

AOI21xp5_ASAP7_75t_L g10772 ( 
.A1(n_10461),
.A2(n_804),
.B(n_806),
.Y(n_10772)
);

INVx1_ASAP7_75t_L g10773 ( 
.A(n_10026),
.Y(n_10773)
);

OAI22xp5_ASAP7_75t_L g10774 ( 
.A1(n_10424),
.A2(n_808),
.B1(n_804),
.B2(n_807),
.Y(n_10774)
);

INVx1_ASAP7_75t_L g10775 ( 
.A(n_10044),
.Y(n_10775)
);

INVx3_ASAP7_75t_L g10776 ( 
.A(n_10516),
.Y(n_10776)
);

A2O1A1Ixp33_ASAP7_75t_L g10777 ( 
.A1(n_10009),
.A2(n_809),
.B(n_807),
.C(n_808),
.Y(n_10777)
);

AOI22xp33_ASAP7_75t_L g10778 ( 
.A1(n_9918),
.A2(n_812),
.B1(n_810),
.B2(n_811),
.Y(n_10778)
);

INVx2_ASAP7_75t_L g10779 ( 
.A(n_10209),
.Y(n_10779)
);

NAND2xp5_ASAP7_75t_L g10780 ( 
.A(n_10045),
.B(n_10081),
.Y(n_10780)
);

HB1xp67_ASAP7_75t_L g10781 ( 
.A(n_10225),
.Y(n_10781)
);

AND2x2_ASAP7_75t_L g10782 ( 
.A(n_10297),
.B(n_811),
.Y(n_10782)
);

NAND2xp5_ASAP7_75t_SL g10783 ( 
.A(n_10153),
.B(n_10220),
.Y(n_10783)
);

NOR2xp33_ASAP7_75t_L g10784 ( 
.A(n_9930),
.B(n_813),
.Y(n_10784)
);

BUFx6f_ASAP7_75t_L g10785 ( 
.A(n_10534),
.Y(n_10785)
);

AOI21xp5_ASAP7_75t_L g10786 ( 
.A1(n_10470),
.A2(n_813),
.B(n_814),
.Y(n_10786)
);

INVx5_ASAP7_75t_L g10787 ( 
.A(n_10208),
.Y(n_10787)
);

NAND2xp5_ASAP7_75t_L g10788 ( 
.A(n_9933),
.B(n_814),
.Y(n_10788)
);

AOI21xp5_ASAP7_75t_L g10789 ( 
.A1(n_10472),
.A2(n_815),
.B(n_816),
.Y(n_10789)
);

AOI22xp5_ASAP7_75t_L g10790 ( 
.A1(n_10127),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.Y(n_10790)
);

NAND2xp5_ASAP7_75t_L g10791 ( 
.A(n_9852),
.B(n_817),
.Y(n_10791)
);

BUFx2_ASAP7_75t_L g10792 ( 
.A(n_10337),
.Y(n_10792)
);

INVx3_ASAP7_75t_L g10793 ( 
.A(n_10534),
.Y(n_10793)
);

BUFx4f_ASAP7_75t_L g10794 ( 
.A(n_10361),
.Y(n_10794)
);

O2A1O1Ixp5_ASAP7_75t_L g10795 ( 
.A1(n_10102),
.A2(n_822),
.B(n_818),
.C(n_821),
.Y(n_10795)
);

AOI21xp5_ASAP7_75t_L g10796 ( 
.A1(n_10475),
.A2(n_821),
.B(n_822),
.Y(n_10796)
);

BUFx2_ASAP7_75t_L g10797 ( 
.A(n_10077),
.Y(n_10797)
);

INVx4_ASAP7_75t_L g10798 ( 
.A(n_10361),
.Y(n_10798)
);

INVx1_ASAP7_75t_L g10799 ( 
.A(n_10339),
.Y(n_10799)
);

INVx2_ASAP7_75t_L g10800 ( 
.A(n_9856),
.Y(n_10800)
);

INVx2_ASAP7_75t_L g10801 ( 
.A(n_9888),
.Y(n_10801)
);

O2A1O1Ixp33_ASAP7_75t_L g10802 ( 
.A1(n_10429),
.A2(n_825),
.B(n_823),
.C(n_824),
.Y(n_10802)
);

NAND2x1p5_ASAP7_75t_L g10803 ( 
.A(n_10143),
.B(n_10333),
.Y(n_10803)
);

BUFx6f_ASAP7_75t_L g10804 ( 
.A(n_10282),
.Y(n_10804)
);

BUFx4f_ASAP7_75t_L g10805 ( 
.A(n_10233),
.Y(n_10805)
);

A2O1A1Ixp33_ASAP7_75t_L g10806 ( 
.A1(n_10028),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_10806)
);

A2O1A1Ixp33_ASAP7_75t_L g10807 ( 
.A1(n_10269),
.A2(n_829),
.B(n_827),
.C(n_828),
.Y(n_10807)
);

O2A1O1Ixp33_ASAP7_75t_SL g10808 ( 
.A1(n_10431),
.A2(n_831),
.B(n_828),
.C(n_830),
.Y(n_10808)
);

NOR2xp33_ASAP7_75t_L g10809 ( 
.A(n_9848),
.B(n_830),
.Y(n_10809)
);

INVx4_ASAP7_75t_L g10810 ( 
.A(n_9837),
.Y(n_10810)
);

AOI21xp5_ASAP7_75t_L g10811 ( 
.A1(n_10480),
.A2(n_831),
.B(n_832),
.Y(n_10811)
);

OAI22xp5_ASAP7_75t_L g10812 ( 
.A1(n_10460),
.A2(n_835),
.B1(n_832),
.B2(n_833),
.Y(n_10812)
);

OAI21x1_ASAP7_75t_L g10813 ( 
.A1(n_10529),
.A2(n_833),
.B(n_836),
.Y(n_10813)
);

AOI21xp5_ASAP7_75t_L g10814 ( 
.A1(n_10481),
.A2(n_836),
.B(n_837),
.Y(n_10814)
);

OAI22x1_ASAP7_75t_L g10815 ( 
.A1(n_9937),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.Y(n_10815)
);

AOI21xp5_ASAP7_75t_L g10816 ( 
.A1(n_10483),
.A2(n_838),
.B(n_839),
.Y(n_10816)
);

NAND2xp5_ASAP7_75t_L g10817 ( 
.A(n_9945),
.B(n_840),
.Y(n_10817)
);

BUFx3_ASAP7_75t_L g10818 ( 
.A(n_10241),
.Y(n_10818)
);

NOR2xp33_ASAP7_75t_R g10819 ( 
.A(n_10075),
.B(n_840),
.Y(n_10819)
);

AOI21xp5_ASAP7_75t_L g10820 ( 
.A1(n_10485),
.A2(n_841),
.B(n_842),
.Y(n_10820)
);

INVx1_ASAP7_75t_L g10821 ( 
.A(n_10352),
.Y(n_10821)
);

NAND2xp5_ASAP7_75t_L g10822 ( 
.A(n_9850),
.B(n_841),
.Y(n_10822)
);

O2A1O1Ixp33_ASAP7_75t_L g10823 ( 
.A1(n_10512),
.A2(n_844),
.B(n_842),
.C(n_843),
.Y(n_10823)
);

NAND2xp5_ASAP7_75t_L g10824 ( 
.A(n_9851),
.B(n_843),
.Y(n_10824)
);

O2A1O1Ixp33_ASAP7_75t_L g10825 ( 
.A1(n_10515),
.A2(n_846),
.B(n_844),
.C(n_845),
.Y(n_10825)
);

AOI21xp5_ASAP7_75t_L g10826 ( 
.A1(n_10488),
.A2(n_845),
.B(n_846),
.Y(n_10826)
);

HB1xp67_ASAP7_75t_L g10827 ( 
.A(n_9957),
.Y(n_10827)
);

OAI22xp5_ASAP7_75t_L g10828 ( 
.A1(n_10564),
.A2(n_849),
.B1(n_847),
.B2(n_848),
.Y(n_10828)
);

AOI21xp5_ASAP7_75t_L g10829 ( 
.A1(n_10494),
.A2(n_847),
.B(n_848),
.Y(n_10829)
);

OR2x2_ASAP7_75t_L g10830 ( 
.A(n_10298),
.B(n_849),
.Y(n_10830)
);

NOR2xp33_ASAP7_75t_L g10831 ( 
.A(n_10334),
.B(n_10345),
.Y(n_10831)
);

CKINVDCx8_ASAP7_75t_R g10832 ( 
.A(n_10099),
.Y(n_10832)
);

INVx1_ASAP7_75t_SL g10833 ( 
.A(n_10133),
.Y(n_10833)
);

NAND2xp5_ASAP7_75t_SL g10834 ( 
.A(n_10239),
.B(n_850),
.Y(n_10834)
);

BUFx2_ASAP7_75t_L g10835 ( 
.A(n_10204),
.Y(n_10835)
);

O2A1O1Ixp33_ASAP7_75t_L g10836 ( 
.A1(n_10536),
.A2(n_852),
.B(n_850),
.C(n_851),
.Y(n_10836)
);

AOI21xp5_ASAP7_75t_L g10837 ( 
.A1(n_10496),
.A2(n_851),
.B(n_852),
.Y(n_10837)
);

AOI21xp5_ASAP7_75t_L g10838 ( 
.A1(n_10497),
.A2(n_853),
.B(n_854),
.Y(n_10838)
);

NAND2xp5_ASAP7_75t_L g10839 ( 
.A(n_10389),
.B(n_854),
.Y(n_10839)
);

BUFx2_ASAP7_75t_L g10840 ( 
.A(n_10295),
.Y(n_10840)
);

INVx3_ASAP7_75t_L g10841 ( 
.A(n_9842),
.Y(n_10841)
);

AOI21xp5_ASAP7_75t_L g10842 ( 
.A1(n_10505),
.A2(n_855),
.B(n_856),
.Y(n_10842)
);

INVx4_ASAP7_75t_L g10843 ( 
.A(n_10433),
.Y(n_10843)
);

NAND2xp5_ASAP7_75t_L g10844 ( 
.A(n_10392),
.B(n_855),
.Y(n_10844)
);

BUFx6f_ASAP7_75t_L g10845 ( 
.A(n_9901),
.Y(n_10845)
);

NOR2xp33_ASAP7_75t_L g10846 ( 
.A(n_10457),
.B(n_856),
.Y(n_10846)
);

BUFx2_ASAP7_75t_L g10847 ( 
.A(n_9983),
.Y(n_10847)
);

AOI22xp33_ASAP7_75t_SL g10848 ( 
.A1(n_10364),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_10848)
);

AOI22xp33_ASAP7_75t_L g10849 ( 
.A1(n_10021),
.A2(n_860),
.B1(n_857),
.B2(n_859),
.Y(n_10849)
);

INVx1_ASAP7_75t_L g10850 ( 
.A(n_9894),
.Y(n_10850)
);

BUFx3_ASAP7_75t_L g10851 ( 
.A(n_10562),
.Y(n_10851)
);

AOI21x1_ASAP7_75t_L g10852 ( 
.A1(n_9976),
.A2(n_860),
.B(n_861),
.Y(n_10852)
);

BUFx2_ASAP7_75t_L g10853 ( 
.A(n_10397),
.Y(n_10853)
);

OAI22x1_ASAP7_75t_L g10854 ( 
.A1(n_10135),
.A2(n_864),
.B1(n_862),
.B2(n_863),
.Y(n_10854)
);

BUFx2_ASAP7_75t_L g10855 ( 
.A(n_10406),
.Y(n_10855)
);

NAND2xp5_ASAP7_75t_L g10856 ( 
.A(n_10414),
.B(n_862),
.Y(n_10856)
);

INVx1_ASAP7_75t_L g10857 ( 
.A(n_9902),
.Y(n_10857)
);

NAND2xp33_ASAP7_75t_L g10858 ( 
.A(n_10551),
.B(n_863),
.Y(n_10858)
);

INVxp67_ASAP7_75t_L g10859 ( 
.A(n_10115),
.Y(n_10859)
);

BUFx12f_ASAP7_75t_L g10860 ( 
.A(n_10233),
.Y(n_10860)
);

A2O1A1Ixp33_ASAP7_75t_L g10861 ( 
.A1(n_10113),
.A2(n_866),
.B(n_864),
.C(n_865),
.Y(n_10861)
);

OAI22xp5_ASAP7_75t_L g10862 ( 
.A1(n_10421),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.Y(n_10862)
);

NAND2xp5_ASAP7_75t_SL g10863 ( 
.A(n_10240),
.B(n_10231),
.Y(n_10863)
);

A2O1A1Ixp33_ASAP7_75t_L g10864 ( 
.A1(n_10124),
.A2(n_869),
.B(n_867),
.C(n_868),
.Y(n_10864)
);

AO32x1_ASAP7_75t_L g10865 ( 
.A1(n_10403),
.A2(n_870),
.A3(n_868),
.B1(n_869),
.B2(n_871),
.Y(n_10865)
);

AOI21xp5_ASAP7_75t_L g10866 ( 
.A1(n_10510),
.A2(n_870),
.B(n_872),
.Y(n_10866)
);

A2O1A1Ixp33_ASAP7_75t_L g10867 ( 
.A1(n_9845),
.A2(n_875),
.B(n_873),
.C(n_874),
.Y(n_10867)
);

BUFx4f_ASAP7_75t_SL g10868 ( 
.A(n_9889),
.Y(n_10868)
);

OAI22xp5_ASAP7_75t_L g10869 ( 
.A1(n_10408),
.A2(n_876),
.B1(n_874),
.B2(n_875),
.Y(n_10869)
);

AOI21xp5_ASAP7_75t_L g10870 ( 
.A1(n_10520),
.A2(n_876),
.B(n_877),
.Y(n_10870)
);

AOI21xp5_ASAP7_75t_L g10871 ( 
.A1(n_10521),
.A2(n_877),
.B(n_878),
.Y(n_10871)
);

OAI21xp5_ASAP7_75t_L g10872 ( 
.A1(n_10531),
.A2(n_880),
.B(n_881),
.Y(n_10872)
);

O2A1O1Ixp33_ASAP7_75t_L g10873 ( 
.A1(n_10559),
.A2(n_884),
.B(n_880),
.C(n_883),
.Y(n_10873)
);

NOR2xp33_ASAP7_75t_L g10874 ( 
.A(n_10126),
.B(n_883),
.Y(n_10874)
);

NAND2xp5_ASAP7_75t_L g10875 ( 
.A(n_10428),
.B(n_884),
.Y(n_10875)
);

NAND2xp5_ASAP7_75t_L g10876 ( 
.A(n_10439),
.B(n_885),
.Y(n_10876)
);

INVx3_ASAP7_75t_L g10877 ( 
.A(n_9998),
.Y(n_10877)
);

OAI21x1_ASAP7_75t_L g10878 ( 
.A1(n_10393),
.A2(n_885),
.B(n_886),
.Y(n_10878)
);

OAI22xp5_ASAP7_75t_L g10879 ( 
.A1(n_9892),
.A2(n_888),
.B1(n_886),
.B2(n_887),
.Y(n_10879)
);

NAND2xp5_ASAP7_75t_SL g10880 ( 
.A(n_10186),
.B(n_10189),
.Y(n_10880)
);

AOI21xp5_ASAP7_75t_L g10881 ( 
.A1(n_10540),
.A2(n_888),
.B(n_889),
.Y(n_10881)
);

AND2x4_ASAP7_75t_L g10882 ( 
.A(n_10383),
.B(n_889),
.Y(n_10882)
);

INVx1_ASAP7_75t_L g10883 ( 
.A(n_9915),
.Y(n_10883)
);

A2O1A1Ixp33_ASAP7_75t_L g10884 ( 
.A1(n_10198),
.A2(n_9854),
.B(n_9866),
.C(n_10175),
.Y(n_10884)
);

INVx1_ASAP7_75t_SL g10885 ( 
.A(n_9913),
.Y(n_10885)
);

NAND2xp5_ASAP7_75t_L g10886 ( 
.A(n_10447),
.B(n_890),
.Y(n_10886)
);

INVx2_ASAP7_75t_L g10887 ( 
.A(n_9960),
.Y(n_10887)
);

NOR3xp33_ASAP7_75t_L g10888 ( 
.A(n_10036),
.B(n_890),
.C(n_891),
.Y(n_10888)
);

INVx1_ASAP7_75t_L g10889 ( 
.A(n_9963),
.Y(n_10889)
);

OAI21x1_ASAP7_75t_L g10890 ( 
.A1(n_10396),
.A2(n_891),
.B(n_892),
.Y(n_10890)
);

O2A1O1Ixp33_ASAP7_75t_L g10891 ( 
.A1(n_10250),
.A2(n_894),
.B(n_892),
.C(n_893),
.Y(n_10891)
);

HB1xp67_ASAP7_75t_L g10892 ( 
.A(n_10450),
.Y(n_10892)
);

AND2x2_ASAP7_75t_L g10893 ( 
.A(n_10388),
.B(n_894),
.Y(n_10893)
);

AOI21xp5_ASAP7_75t_L g10894 ( 
.A1(n_10544),
.A2(n_895),
.B(n_896),
.Y(n_10894)
);

AOI22xp5_ASAP7_75t_L g10895 ( 
.A1(n_10259),
.A2(n_897),
.B1(n_895),
.B2(n_896),
.Y(n_10895)
);

NAND2xp5_ASAP7_75t_L g10896 ( 
.A(n_10451),
.B(n_897),
.Y(n_10896)
);

OAI22xp5_ASAP7_75t_L g10897 ( 
.A1(n_10049),
.A2(n_900),
.B1(n_898),
.B2(n_899),
.Y(n_10897)
);

O2A1O1Ixp33_ASAP7_75t_L g10898 ( 
.A1(n_10349),
.A2(n_900),
.B(n_898),
.C(n_899),
.Y(n_10898)
);

NOR2xp33_ASAP7_75t_L g10899 ( 
.A(n_9905),
.B(n_901),
.Y(n_10899)
);

CKINVDCx5p33_ASAP7_75t_R g10900 ( 
.A(n_9925),
.Y(n_10900)
);

BUFx3_ASAP7_75t_L g10901 ( 
.A(n_10207),
.Y(n_10901)
);

AOI21xp5_ASAP7_75t_L g10902 ( 
.A1(n_10545),
.A2(n_901),
.B(n_902),
.Y(n_10902)
);

INVxp67_ASAP7_75t_SL g10903 ( 
.A(n_10444),
.Y(n_10903)
);

NAND2xp5_ASAP7_75t_L g10904 ( 
.A(n_10463),
.B(n_902),
.Y(n_10904)
);

OR2x2_ASAP7_75t_L g10905 ( 
.A(n_10464),
.B(n_903),
.Y(n_10905)
);

AO21x2_ASAP7_75t_L g10906 ( 
.A1(n_10006),
.A2(n_10342),
.B(n_10328),
.Y(n_10906)
);

INVx3_ASAP7_75t_L g10907 ( 
.A(n_10156),
.Y(n_10907)
);

INVx1_ASAP7_75t_L g10908 ( 
.A(n_9991),
.Y(n_10908)
);

NAND2xp5_ASAP7_75t_SL g10909 ( 
.A(n_10193),
.B(n_903),
.Y(n_10909)
);

O2A1O1Ixp33_ASAP7_75t_L g10910 ( 
.A1(n_10356),
.A2(n_906),
.B(n_904),
.C(n_905),
.Y(n_10910)
);

A2O1A1Ixp33_ASAP7_75t_L g10911 ( 
.A1(n_10037),
.A2(n_907),
.B(n_905),
.C(n_906),
.Y(n_10911)
);

OAI22xp5_ASAP7_75t_L g10912 ( 
.A1(n_10324),
.A2(n_909),
.B1(n_907),
.B2(n_908),
.Y(n_10912)
);

AND2x2_ASAP7_75t_L g10913 ( 
.A(n_10434),
.B(n_908),
.Y(n_10913)
);

NAND2xp5_ASAP7_75t_L g10914 ( 
.A(n_10469),
.B(n_910),
.Y(n_10914)
);

BUFx6f_ASAP7_75t_L g10915 ( 
.A(n_10422),
.Y(n_10915)
);

INVx1_ASAP7_75t_L g10916 ( 
.A(n_10039),
.Y(n_10916)
);

NAND2xp5_ASAP7_75t_L g10917 ( 
.A(n_10473),
.B(n_910),
.Y(n_10917)
);

NOR2xp67_ASAP7_75t_L g10918 ( 
.A(n_10210),
.B(n_911),
.Y(n_10918)
);

INVxp67_ASAP7_75t_L g10919 ( 
.A(n_10486),
.Y(n_10919)
);

INVx2_ASAP7_75t_L g10920 ( 
.A(n_10071),
.Y(n_10920)
);

NAND2xp5_ASAP7_75t_SL g10921 ( 
.A(n_10199),
.B(n_911),
.Y(n_10921)
);

OAI21x1_ASAP7_75t_L g10922 ( 
.A1(n_10401),
.A2(n_914),
.B(n_915),
.Y(n_10922)
);

NOR2xp33_ASAP7_75t_L g10923 ( 
.A(n_9940),
.B(n_914),
.Y(n_10923)
);

NAND2xp5_ASAP7_75t_L g10924 ( 
.A(n_10489),
.B(n_915),
.Y(n_10924)
);

NAND2xp5_ASAP7_75t_SL g10925 ( 
.A(n_10206),
.B(n_916),
.Y(n_10925)
);

AOI21xp5_ASAP7_75t_L g10926 ( 
.A1(n_10550),
.A2(n_916),
.B(n_917),
.Y(n_10926)
);

INVx1_ASAP7_75t_L g10927 ( 
.A(n_10106),
.Y(n_10927)
);

INVx1_ASAP7_75t_L g10928 ( 
.A(n_10109),
.Y(n_10928)
);

INVx2_ASAP7_75t_L g10929 ( 
.A(n_10129),
.Y(n_10929)
);

NAND2xp5_ASAP7_75t_L g10930 ( 
.A(n_10490),
.B(n_918),
.Y(n_10930)
);

INVx1_ASAP7_75t_L g10931 ( 
.A(n_10157),
.Y(n_10931)
);

A2O1A1Ixp33_ASAP7_75t_SL g10932 ( 
.A1(n_10554),
.A2(n_921),
.B(n_918),
.C(n_920),
.Y(n_10932)
);

NAND2xp5_ASAP7_75t_L g10933 ( 
.A(n_10501),
.B(n_920),
.Y(n_10933)
);

INVx3_ASAP7_75t_L g10934 ( 
.A(n_10405),
.Y(n_10934)
);

INVx2_ASAP7_75t_L g10935 ( 
.A(n_10195),
.Y(n_10935)
);

BUFx12f_ASAP7_75t_L g10936 ( 
.A(n_10508),
.Y(n_10936)
);

INVx1_ASAP7_75t_L g10937 ( 
.A(n_10200),
.Y(n_10937)
);

INVx1_ASAP7_75t_L g10938 ( 
.A(n_10203),
.Y(n_10938)
);

AOI21xp5_ASAP7_75t_L g10939 ( 
.A1(n_10560),
.A2(n_921),
.B(n_922),
.Y(n_10939)
);

INVx3_ASAP7_75t_L g10940 ( 
.A(n_10336),
.Y(n_10940)
);

BUFx4f_ASAP7_75t_L g10941 ( 
.A(n_10478),
.Y(n_10941)
);

AOI21xp5_ASAP7_75t_L g10942 ( 
.A1(n_10561),
.A2(n_922),
.B(n_923),
.Y(n_10942)
);

AND2x2_ASAP7_75t_L g10943 ( 
.A(n_10513),
.B(n_923),
.Y(n_10943)
);

NAND2xp5_ASAP7_75t_L g10944 ( 
.A(n_10527),
.B(n_10541),
.Y(n_10944)
);

HB1xp67_ASAP7_75t_L g10945 ( 
.A(n_10553),
.Y(n_10945)
);

O2A1O1Ixp33_ASAP7_75t_L g10946 ( 
.A1(n_10286),
.A2(n_927),
.B(n_924),
.C(n_926),
.Y(n_10946)
);

BUFx2_ASAP7_75t_L g10947 ( 
.A(n_10048),
.Y(n_10947)
);

NAND2xp5_ASAP7_75t_L g10948 ( 
.A(n_10056),
.B(n_924),
.Y(n_10948)
);

O2A1O1Ixp33_ASAP7_75t_L g10949 ( 
.A1(n_10367),
.A2(n_928),
.B(n_926),
.C(n_927),
.Y(n_10949)
);

AOI21xp5_ASAP7_75t_L g10950 ( 
.A1(n_10082),
.A2(n_928),
.B(n_929),
.Y(n_10950)
);

NOR2xp33_ASAP7_75t_L g10951 ( 
.A(n_9969),
.B(n_929),
.Y(n_10951)
);

NAND2xp5_ASAP7_75t_SL g10952 ( 
.A(n_10222),
.B(n_930),
.Y(n_10952)
);

NAND2xp5_ASAP7_75t_L g10953 ( 
.A(n_10062),
.B(n_930),
.Y(n_10953)
);

INVx2_ASAP7_75t_L g10954 ( 
.A(n_10221),
.Y(n_10954)
);

NOR2xp33_ASAP7_75t_R g10955 ( 
.A(n_10285),
.B(n_931),
.Y(n_10955)
);

AOI21xp5_ASAP7_75t_L g10956 ( 
.A1(n_10082),
.A2(n_932),
.B(n_933),
.Y(n_10956)
);

CKINVDCx20_ASAP7_75t_R g10957 ( 
.A(n_10122),
.Y(n_10957)
);

AOI21xp5_ASAP7_75t_L g10958 ( 
.A1(n_9880),
.A2(n_932),
.B(n_934),
.Y(n_10958)
);

NOR2xp33_ASAP7_75t_L g10959 ( 
.A(n_9984),
.B(n_934),
.Y(n_10959)
);

NOR2xp33_ASAP7_75t_L g10960 ( 
.A(n_10362),
.B(n_935),
.Y(n_10960)
);

NAND2xp5_ASAP7_75t_SL g10961 ( 
.A(n_9974),
.B(n_936),
.Y(n_10961)
);

INVx2_ASAP7_75t_L g10962 ( 
.A(n_10244),
.Y(n_10962)
);

BUFx3_ASAP7_75t_L g10963 ( 
.A(n_9955),
.Y(n_10963)
);

INVx1_ASAP7_75t_L g10964 ( 
.A(n_10256),
.Y(n_10964)
);

BUFx6f_ASAP7_75t_L g10965 ( 
.A(n_10296),
.Y(n_10965)
);

NAND2xp5_ASAP7_75t_L g10966 ( 
.A(n_10065),
.B(n_937),
.Y(n_10966)
);

CKINVDCx5p33_ASAP7_75t_R g10967 ( 
.A(n_10228),
.Y(n_10967)
);

BUFx3_ASAP7_75t_L g10968 ( 
.A(n_10248),
.Y(n_10968)
);

AOI21xp5_ASAP7_75t_L g10969 ( 
.A1(n_10000),
.A2(n_938),
.B(n_939),
.Y(n_10969)
);

NAND2xp5_ASAP7_75t_SL g10970 ( 
.A(n_10452),
.B(n_938),
.Y(n_10970)
);

NOR2xp33_ASAP7_75t_R g10971 ( 
.A(n_10144),
.B(n_939),
.Y(n_10971)
);

BUFx6f_ASAP7_75t_L g10972 ( 
.A(n_10312),
.Y(n_10972)
);

INVx3_ASAP7_75t_L g10973 ( 
.A(n_10321),
.Y(n_10973)
);

NOR2xp67_ASAP7_75t_SL g10974 ( 
.A(n_10008),
.B(n_940),
.Y(n_10974)
);

AND2x2_ASAP7_75t_L g10975 ( 
.A(n_10003),
.B(n_940),
.Y(n_10975)
);

NOR3xp33_ASAP7_75t_SL g10976 ( 
.A(n_10161),
.B(n_941),
.C(n_942),
.Y(n_10976)
);

NOR2xp33_ASAP7_75t_SL g10977 ( 
.A(n_9944),
.B(n_941),
.Y(n_10977)
);

NAND2xp5_ASAP7_75t_L g10978 ( 
.A(n_10067),
.B(n_943),
.Y(n_10978)
);

NOR2xp33_ASAP7_75t_L g10979 ( 
.A(n_10277),
.B(n_943),
.Y(n_10979)
);

OAI21x1_ASAP7_75t_L g10980 ( 
.A1(n_10459),
.A2(n_944),
.B(n_945),
.Y(n_10980)
);

A2O1A1Ixp33_ASAP7_75t_L g10981 ( 
.A1(n_9959),
.A2(n_947),
.B(n_944),
.C(n_946),
.Y(n_10981)
);

A2O1A1Ixp33_ASAP7_75t_L g10982 ( 
.A1(n_10130),
.A2(n_949),
.B(n_946),
.C(n_948),
.Y(n_10982)
);

AOI21xp5_ASAP7_75t_L g10983 ( 
.A1(n_10000),
.A2(n_10332),
.B(n_9906),
.Y(n_10983)
);

NAND2xp5_ASAP7_75t_L g10984 ( 
.A(n_10072),
.B(n_948),
.Y(n_10984)
);

AOI21xp5_ASAP7_75t_L g10985 ( 
.A1(n_10111),
.A2(n_949),
.B(n_950),
.Y(n_10985)
);

BUFx3_ASAP7_75t_L g10986 ( 
.A(n_10325),
.Y(n_10986)
);

A2O1A1Ixp33_ASAP7_75t_L g10987 ( 
.A1(n_10128),
.A2(n_952),
.B(n_950),
.C(n_951),
.Y(n_10987)
);

NAND2xp5_ASAP7_75t_L g10988 ( 
.A(n_10076),
.B(n_951),
.Y(n_10988)
);

NOR2xp67_ASAP7_75t_SL g10989 ( 
.A(n_10254),
.B(n_952),
.Y(n_10989)
);

INVx1_ASAP7_75t_L g10990 ( 
.A(n_10315),
.Y(n_10990)
);

OAI22xp5_ASAP7_75t_L g10991 ( 
.A1(n_10340),
.A2(n_955),
.B1(n_953),
.B2(n_954),
.Y(n_10991)
);

CKINVDCx20_ASAP7_75t_R g10992 ( 
.A(n_10279),
.Y(n_10992)
);

AOI21xp5_ASAP7_75t_L g10993 ( 
.A1(n_9878),
.A2(n_954),
.B(n_956),
.Y(n_10993)
);

NAND2xp5_ASAP7_75t_SL g10994 ( 
.A(n_10539),
.B(n_956),
.Y(n_10994)
);

AOI21xp5_ASAP7_75t_L g10995 ( 
.A1(n_9989),
.A2(n_957),
.B(n_959),
.Y(n_10995)
);

INVx1_ASAP7_75t_L g10996 ( 
.A(n_10343),
.Y(n_10996)
);

INVx1_ASAP7_75t_SL g10997 ( 
.A(n_10381),
.Y(n_10997)
);

OR2x6_ASAP7_75t_L g10998 ( 
.A(n_9951),
.B(n_957),
.Y(n_10998)
);

INVx2_ASAP7_75t_L g10999 ( 
.A(n_10344),
.Y(n_10999)
);

BUFx6f_ASAP7_75t_L g11000 ( 
.A(n_10359),
.Y(n_11000)
);

BUFx6f_ASAP7_75t_L g11001 ( 
.A(n_10372),
.Y(n_11001)
);

BUFx3_ASAP7_75t_L g11002 ( 
.A(n_10271),
.Y(n_11002)
);

INVx1_ASAP7_75t_L g11003 ( 
.A(n_10399),
.Y(n_11003)
);

BUFx2_ASAP7_75t_L g11004 ( 
.A(n_10086),
.Y(n_11004)
);

OAI22xp5_ASAP7_75t_L g11005 ( 
.A1(n_9859),
.A2(n_961),
.B1(n_959),
.B2(n_960),
.Y(n_11005)
);

NAND2xp5_ASAP7_75t_SL g11006 ( 
.A(n_10171),
.B(n_960),
.Y(n_11006)
);

OAI22xp5_ASAP7_75t_L g11007 ( 
.A1(n_9975),
.A2(n_963),
.B1(n_961),
.B2(n_962),
.Y(n_11007)
);

NOR3xp33_ASAP7_75t_SL g11008 ( 
.A(n_10073),
.B(n_962),
.C(n_963),
.Y(n_11008)
);

OAI22xp5_ASAP7_75t_L g11009 ( 
.A1(n_10079),
.A2(n_966),
.B1(n_964),
.B2(n_965),
.Y(n_11009)
);

INVx1_ASAP7_75t_L g11010 ( 
.A(n_10416),
.Y(n_11010)
);

NOR2xp33_ASAP7_75t_L g11011 ( 
.A(n_10060),
.B(n_964),
.Y(n_11011)
);

AOI21xp5_ASAP7_75t_L g11012 ( 
.A1(n_10050),
.A2(n_966),
.B(n_967),
.Y(n_11012)
);

INVxp67_ASAP7_75t_L g11013 ( 
.A(n_10227),
.Y(n_11013)
);

A2O1A1Ixp33_ASAP7_75t_L g11014 ( 
.A1(n_10017),
.A2(n_10176),
.B(n_10319),
.C(n_10280),
.Y(n_11014)
);

AOI21xp5_ASAP7_75t_L g11015 ( 
.A1(n_9903),
.A2(n_967),
.B(n_968),
.Y(n_11015)
);

NAND2x1p5_ASAP7_75t_L g11016 ( 
.A(n_9891),
.B(n_9900),
.Y(n_11016)
);

OAI22xp5_ASAP7_75t_L g11017 ( 
.A1(n_9923),
.A2(n_971),
.B1(n_968),
.B2(n_969),
.Y(n_11017)
);

AOI22xp33_ASAP7_75t_L g11018 ( 
.A1(n_10030),
.A2(n_972),
.B1(n_969),
.B2(n_971),
.Y(n_11018)
);

NAND2xp5_ASAP7_75t_L g11019 ( 
.A(n_10088),
.B(n_972),
.Y(n_11019)
);

NAND2xp5_ASAP7_75t_L g11020 ( 
.A(n_10090),
.B(n_973),
.Y(n_11020)
);

NOR2xp67_ASAP7_75t_SL g11021 ( 
.A(n_10238),
.B(n_973),
.Y(n_11021)
);

BUFx12f_ASAP7_75t_L g11022 ( 
.A(n_10095),
.Y(n_11022)
);

AOI21xp5_ASAP7_75t_L g11023 ( 
.A1(n_9911),
.A2(n_974),
.B(n_975),
.Y(n_11023)
);

AOI221xp5_ASAP7_75t_L g11024 ( 
.A1(n_10419),
.A2(n_976),
.B1(n_974),
.B2(n_975),
.C(n_977),
.Y(n_11024)
);

A2O1A1Ixp33_ASAP7_75t_SL g11025 ( 
.A1(n_9855),
.A2(n_978),
.B(n_976),
.C(n_977),
.Y(n_11025)
);

AOI21xp5_ASAP7_75t_L g11026 ( 
.A1(n_9916),
.A2(n_978),
.B(n_979),
.Y(n_11026)
);

INVx2_ASAP7_75t_L g11027 ( 
.A(n_10436),
.Y(n_11027)
);

AOI21xp5_ASAP7_75t_L g11028 ( 
.A1(n_10410),
.A2(n_979),
.B(n_980),
.Y(n_11028)
);

NOR2xp67_ASAP7_75t_L g11029 ( 
.A(n_10232),
.B(n_980),
.Y(n_11029)
);

AND2x2_ASAP7_75t_L g11030 ( 
.A(n_10134),
.B(n_981),
.Y(n_11030)
);

NAND2xp5_ASAP7_75t_SL g11031 ( 
.A(n_10158),
.B(n_981),
.Y(n_11031)
);

NAND2xp5_ASAP7_75t_SL g11032 ( 
.A(n_9934),
.B(n_982),
.Y(n_11032)
);

CKINVDCx5p33_ASAP7_75t_R g11033 ( 
.A(n_10185),
.Y(n_11033)
);

O2A1O1Ixp33_ASAP7_75t_L g11034 ( 
.A1(n_10376),
.A2(n_984),
.B(n_982),
.C(n_983),
.Y(n_11034)
);

INVx1_ASAP7_75t_L g11035 ( 
.A(n_10441),
.Y(n_11035)
);

AOI21xp5_ASAP7_75t_L g11036 ( 
.A1(n_10444),
.A2(n_983),
.B(n_984),
.Y(n_11036)
);

AOI22xp5_ASAP7_75t_L g11037 ( 
.A1(n_10263),
.A2(n_987),
.B1(n_985),
.B2(n_986),
.Y(n_11037)
);

AOI21xp5_ASAP7_75t_L g11038 ( 
.A1(n_9968),
.A2(n_986),
.B(n_987),
.Y(n_11038)
);

NAND2xp5_ASAP7_75t_L g11039 ( 
.A(n_10091),
.B(n_989),
.Y(n_11039)
);

NAND2xp5_ASAP7_75t_L g11040 ( 
.A(n_9985),
.B(n_989),
.Y(n_11040)
);

O2A1O1Ixp33_ASAP7_75t_L g11041 ( 
.A1(n_10293),
.A2(n_992),
.B(n_990),
.C(n_991),
.Y(n_11041)
);

NAND2xp5_ASAP7_75t_L g11042 ( 
.A(n_9987),
.B(n_9992),
.Y(n_11042)
);

NOR2xp33_ASAP7_75t_L g11043 ( 
.A(n_10080),
.B(n_991),
.Y(n_11043)
);

AND2x2_ASAP7_75t_L g11044 ( 
.A(n_10187),
.B(n_992),
.Y(n_11044)
);

NOR3xp33_ASAP7_75t_SL g11045 ( 
.A(n_9867),
.B(n_993),
.C(n_994),
.Y(n_11045)
);

NAND2xp5_ASAP7_75t_L g11046 ( 
.A(n_9997),
.B(n_993),
.Y(n_11046)
);

INVx3_ASAP7_75t_L g11047 ( 
.A(n_10320),
.Y(n_11047)
);

AOI21xp5_ASAP7_75t_L g11048 ( 
.A1(n_10074),
.A2(n_994),
.B(n_995),
.Y(n_11048)
);

INVx2_ASAP7_75t_L g11049 ( 
.A(n_10454),
.Y(n_11049)
);

AOI21xp5_ASAP7_75t_L g11050 ( 
.A1(n_9952),
.A2(n_995),
.B(n_996),
.Y(n_11050)
);

A2O1A1Ixp33_ASAP7_75t_L g11051 ( 
.A1(n_10289),
.A2(n_998),
.B(n_996),
.C(n_997),
.Y(n_11051)
);

AOI21xp5_ASAP7_75t_L g11052 ( 
.A1(n_9961),
.A2(n_10147),
.B(n_10146),
.Y(n_11052)
);

NOR2xp33_ASAP7_75t_L g11053 ( 
.A(n_10120),
.B(n_997),
.Y(n_11053)
);

INVx1_ASAP7_75t_L g11054 ( 
.A(n_10491),
.Y(n_11054)
);

BUFx12f_ASAP7_75t_L g11055 ( 
.A(n_10194),
.Y(n_11055)
);

INVx1_ASAP7_75t_L g11056 ( 
.A(n_10504),
.Y(n_11056)
);

INVx1_ASAP7_75t_SL g11057 ( 
.A(n_10202),
.Y(n_11057)
);

AOI21xp5_ASAP7_75t_L g11058 ( 
.A1(n_9967),
.A2(n_998),
.B(n_999),
.Y(n_11058)
);

A2O1A1Ixp33_ASAP7_75t_L g11059 ( 
.A1(n_10291),
.A2(n_1001),
.B(n_999),
.C(n_1000),
.Y(n_11059)
);

INVx5_ASAP7_75t_L g11060 ( 
.A(n_10384),
.Y(n_11060)
);

INVx3_ASAP7_75t_L g11061 ( 
.A(n_10211),
.Y(n_11061)
);

INVx4_ASAP7_75t_L g11062 ( 
.A(n_10507),
.Y(n_11062)
);

AND2x2_ASAP7_75t_L g11063 ( 
.A(n_10224),
.B(n_1000),
.Y(n_11063)
);

OR2x6_ASAP7_75t_L g11064 ( 
.A(n_10305),
.B(n_1001),
.Y(n_11064)
);

NAND2xp5_ASAP7_75t_L g11065 ( 
.A(n_9999),
.B(n_1002),
.Y(n_11065)
);

NOR3xp33_ASAP7_75t_L g11066 ( 
.A(n_10253),
.B(n_1002),
.C(n_1003),
.Y(n_11066)
);

NAND2xp5_ASAP7_75t_L g11067 ( 
.A(n_10011),
.B(n_1003),
.Y(n_11067)
);

INVx1_ASAP7_75t_L g11068 ( 
.A(n_10514),
.Y(n_11068)
);

AND2x4_ASAP7_75t_L g11069 ( 
.A(n_10517),
.B(n_1004),
.Y(n_11069)
);

NAND2xp5_ASAP7_75t_SL g11070 ( 
.A(n_10306),
.B(n_1005),
.Y(n_11070)
);

OAI22xp5_ASAP7_75t_L g11071 ( 
.A1(n_10353),
.A2(n_1007),
.B1(n_1005),
.B2(n_1006),
.Y(n_11071)
);

INVx1_ASAP7_75t_L g11072 ( 
.A(n_10528),
.Y(n_11072)
);

AOI22xp5_ASAP7_75t_L g11073 ( 
.A1(n_10404),
.A2(n_1008),
.B1(n_1006),
.B2(n_1007),
.Y(n_11073)
);

INVx1_ASAP7_75t_L g11074 ( 
.A(n_10012),
.Y(n_11074)
);

AOI21xp5_ASAP7_75t_L g11075 ( 
.A1(n_9847),
.A2(n_1008),
.B(n_1009),
.Y(n_11075)
);

NAND2xp5_ASAP7_75t_L g11076 ( 
.A(n_10013),
.B(n_1009),
.Y(n_11076)
);

AOI21xp5_ASAP7_75t_L g11077 ( 
.A1(n_10101),
.A2(n_1011),
.B(n_1012),
.Y(n_11077)
);

BUFx6f_ASAP7_75t_L g11078 ( 
.A(n_10346),
.Y(n_11078)
);

NOR2xp33_ASAP7_75t_L g11079 ( 
.A(n_10251),
.B(n_1012),
.Y(n_11079)
);

INVx5_ASAP7_75t_L g11080 ( 
.A(n_10276),
.Y(n_11080)
);

INVx1_ASAP7_75t_SL g11081 ( 
.A(n_10267),
.Y(n_11081)
);

NAND3xp33_ASAP7_75t_SL g11082 ( 
.A(n_10347),
.B(n_1013),
.C(n_1014),
.Y(n_11082)
);

NAND2xp5_ASAP7_75t_L g11083 ( 
.A(n_10020),
.B(n_1014),
.Y(n_11083)
);

A2O1A1Ixp33_ASAP7_75t_L g11084 ( 
.A1(n_10304),
.A2(n_1017),
.B(n_1015),
.C(n_1016),
.Y(n_11084)
);

OAI22xp5_ASAP7_75t_L g11085 ( 
.A1(n_10307),
.A2(n_1017),
.B1(n_1015),
.B2(n_1016),
.Y(n_11085)
);

AO21x2_ASAP7_75t_L g11086 ( 
.A1(n_10357),
.A2(n_1018),
.B(n_1019),
.Y(n_11086)
);

OAI22xp5_ASAP7_75t_L g11087 ( 
.A1(n_10018),
.A2(n_1021),
.B1(n_1018),
.B2(n_1019),
.Y(n_11087)
);

AOI21xp5_ASAP7_75t_L g11088 ( 
.A1(n_9986),
.A2(n_1021),
.B(n_1022),
.Y(n_11088)
);

AOI21xp5_ASAP7_75t_L g11089 ( 
.A1(n_9877),
.A2(n_1023),
.B(n_1024),
.Y(n_11089)
);

BUFx3_ASAP7_75t_L g11090 ( 
.A(n_10159),
.Y(n_11090)
);

INVx2_ASAP7_75t_SL g11091 ( 
.A(n_9865),
.Y(n_11091)
);

INVx2_ASAP7_75t_L g11092 ( 
.A(n_10363),
.Y(n_11092)
);

AOI21xp5_ASAP7_75t_L g11093 ( 
.A1(n_10354),
.A2(n_1023),
.B(n_1024),
.Y(n_11093)
);

BUFx6f_ASAP7_75t_L g11094 ( 
.A(n_10366),
.Y(n_11094)
);

CKINVDCx20_ASAP7_75t_R g11095 ( 
.A(n_10378),
.Y(n_11095)
);

INVx1_ASAP7_75t_L g11096 ( 
.A(n_10031),
.Y(n_11096)
);

AOI21xp5_ASAP7_75t_L g11097 ( 
.A1(n_10246),
.A2(n_1025),
.B(n_1026),
.Y(n_11097)
);

AND2x6_ASAP7_75t_L g11098 ( 
.A(n_10042),
.B(n_1027),
.Y(n_11098)
);

INVx2_ASAP7_75t_L g11099 ( 
.A(n_10368),
.Y(n_11099)
);

INVx2_ASAP7_75t_L g11100 ( 
.A(n_10369),
.Y(n_11100)
);

NOR2xp33_ASAP7_75t_L g11101 ( 
.A(n_10264),
.B(n_1027),
.Y(n_11101)
);

BUFx6f_ASAP7_75t_L g11102 ( 
.A(n_10373),
.Y(n_11102)
);

INVx2_ASAP7_75t_L g11103 ( 
.A(n_10033),
.Y(n_11103)
);

BUFx6f_ASAP7_75t_L g11104 ( 
.A(n_10301),
.Y(n_11104)
);

AO21x1_ASAP7_75t_L g11105 ( 
.A1(n_9994),
.A2(n_1028),
.B(n_1029),
.Y(n_11105)
);

A2O1A1Ixp33_ASAP7_75t_L g11106 ( 
.A1(n_10358),
.A2(n_1030),
.B(n_1028),
.C(n_1029),
.Y(n_11106)
);

INVx3_ASAP7_75t_L g11107 ( 
.A(n_10116),
.Y(n_11107)
);

OA22x2_ASAP7_75t_L g11108 ( 
.A1(n_10022),
.A2(n_1033),
.B1(n_1030),
.B2(n_1032),
.Y(n_11108)
);

NAND2xp33_ASAP7_75t_SL g11109 ( 
.A(n_10164),
.B(n_1032),
.Y(n_11109)
);

NOR3xp33_ASAP7_75t_SL g11110 ( 
.A(n_10093),
.B(n_1033),
.C(n_1034),
.Y(n_11110)
);

NOR2xp67_ASAP7_75t_L g11111 ( 
.A(n_10107),
.B(n_10108),
.Y(n_11111)
);

BUFx6f_ASAP7_75t_L g11112 ( 
.A(n_10302),
.Y(n_11112)
);

OR2x2_ASAP7_75t_L g11113 ( 
.A(n_10163),
.B(n_1034),
.Y(n_11113)
);

INVx1_ASAP7_75t_L g11114 ( 
.A(n_10448),
.Y(n_11114)
);

INVx1_ASAP7_75t_L g11115 ( 
.A(n_10448),
.Y(n_11115)
);

O2A1O1Ixp33_ASAP7_75t_L g11116 ( 
.A1(n_10310),
.A2(n_10313),
.B(n_9943),
.C(n_10355),
.Y(n_11116)
);

A2O1A1Ixp33_ASAP7_75t_L g11117 ( 
.A1(n_10154),
.A2(n_1037),
.B(n_1035),
.C(n_1036),
.Y(n_11117)
);

AND2x2_ASAP7_75t_L g11118 ( 
.A(n_10299),
.B(n_1035),
.Y(n_11118)
);

AO21x1_ASAP7_75t_L g11119 ( 
.A1(n_10089),
.A2(n_1036),
.B(n_1037),
.Y(n_11119)
);

AOI21x1_ASAP7_75t_L g11120 ( 
.A1(n_10182),
.A2(n_1038),
.B(n_1039),
.Y(n_11120)
);

OAI22xp5_ASAP7_75t_L g11121 ( 
.A1(n_10425),
.A2(n_1041),
.B1(n_1038),
.B2(n_1040),
.Y(n_11121)
);

INVx2_ASAP7_75t_L g11122 ( 
.A(n_10448),
.Y(n_11122)
);

NAND2xp5_ASAP7_75t_SL g11123 ( 
.A(n_10174),
.B(n_1040),
.Y(n_11123)
);

INVx2_ASAP7_75t_L g11124 ( 
.A(n_9860),
.Y(n_11124)
);

HB1xp67_ASAP7_75t_L g11125 ( 
.A(n_9861),
.Y(n_11125)
);

NOR2xp33_ASAP7_75t_L g11126 ( 
.A(n_10300),
.B(n_1041),
.Y(n_11126)
);

INVx3_ASAP7_75t_L g11127 ( 
.A(n_10191),
.Y(n_11127)
);

INVx1_ASAP7_75t_L g11128 ( 
.A(n_9871),
.Y(n_11128)
);

NAND2xp5_ASAP7_75t_L g11129 ( 
.A(n_9884),
.B(n_1042),
.Y(n_11129)
);

INVx2_ASAP7_75t_L g11130 ( 
.A(n_9886),
.Y(n_11130)
);

INVx1_ASAP7_75t_L g11131 ( 
.A(n_9898),
.Y(n_11131)
);

O2A1O1Ixp33_ASAP7_75t_L g11132 ( 
.A1(n_10261),
.A2(n_1044),
.B(n_1042),
.C(n_1043),
.Y(n_11132)
);

INVx1_ASAP7_75t_L g11133 ( 
.A(n_9904),
.Y(n_11133)
);

INVx2_ASAP7_75t_L g11134 ( 
.A(n_9907),
.Y(n_11134)
);

A2O1A1Ixp33_ASAP7_75t_L g11135 ( 
.A1(n_10155),
.A2(n_1046),
.B(n_1043),
.C(n_1045),
.Y(n_11135)
);

NAND2xp5_ASAP7_75t_L g11136 ( 
.A(n_9919),
.B(n_1045),
.Y(n_11136)
);

NAND2xp5_ASAP7_75t_SL g11137 ( 
.A(n_9927),
.B(n_1047),
.Y(n_11137)
);

BUFx10_ASAP7_75t_L g11138 ( 
.A(n_10140),
.Y(n_11138)
);

INVx1_ASAP7_75t_SL g11139 ( 
.A(n_10245),
.Y(n_11139)
);

BUFx2_ASAP7_75t_L g11140 ( 
.A(n_9920),
.Y(n_11140)
);

INVx2_ASAP7_75t_L g11141 ( 
.A(n_9928),
.Y(n_11141)
);

NOR2xp33_ASAP7_75t_L g11142 ( 
.A(n_10247),
.B(n_1047),
.Y(n_11142)
);

NAND2xp5_ASAP7_75t_SL g11143 ( 
.A(n_10257),
.B(n_10112),
.Y(n_11143)
);

BUFx2_ASAP7_75t_L g11144 ( 
.A(n_9935),
.Y(n_11144)
);

BUFx2_ASAP7_75t_L g11145 ( 
.A(n_9936),
.Y(n_11145)
);

NAND2xp5_ASAP7_75t_L g11146 ( 
.A(n_9941),
.B(n_1048),
.Y(n_11146)
);

INVx3_ASAP7_75t_SL g11147 ( 
.A(n_10322),
.Y(n_11147)
);

INVx1_ASAP7_75t_L g11148 ( 
.A(n_9942),
.Y(n_11148)
);

INVx1_ASAP7_75t_L g11149 ( 
.A(n_9981),
.Y(n_11149)
);

NAND2xp5_ASAP7_75t_L g11150 ( 
.A(n_10169),
.B(n_1048),
.Y(n_11150)
);

NAND2xp33_ASAP7_75t_SL g11151 ( 
.A(n_10438),
.B(n_1049),
.Y(n_11151)
);

INVx2_ASAP7_75t_L g11152 ( 
.A(n_10400),
.Y(n_11152)
);

NOR2xp33_ASAP7_75t_L g11153 ( 
.A(n_10117),
.B(n_1049),
.Y(n_11153)
);

AOI22xp5_ASAP7_75t_L g11154 ( 
.A1(n_10449),
.A2(n_1052),
.B1(n_1050),
.B2(n_1051),
.Y(n_11154)
);

O2A1O1Ixp5_ASAP7_75t_L g11155 ( 
.A1(n_10465),
.A2(n_1052),
.B(n_1050),
.C(n_1051),
.Y(n_11155)
);

HB1xp67_ASAP7_75t_L g11156 ( 
.A(n_10525),
.Y(n_11156)
);

NOR2xp33_ASAP7_75t_L g11157 ( 
.A(n_10236),
.B(n_1053),
.Y(n_11157)
);

OAI22xp5_ASAP7_75t_L g11158 ( 
.A1(n_10503),
.A2(n_1055),
.B1(n_1053),
.B2(n_1054),
.Y(n_11158)
);

AOI21xp33_ASAP7_75t_L g11159 ( 
.A1(n_10509),
.A2(n_1054),
.B(n_1055),
.Y(n_11159)
);

AOI22xp5_ASAP7_75t_L g11160 ( 
.A1(n_10537),
.A2(n_9996),
.B1(n_10290),
.B2(n_10258),
.Y(n_11160)
);

INVx2_ASAP7_75t_L g11161 ( 
.A(n_10400),
.Y(n_11161)
);

BUFx6f_ASAP7_75t_L g11162 ( 
.A(n_10149),
.Y(n_11162)
);

AOI21xp5_ASAP7_75t_L g11163 ( 
.A1(n_10148),
.A2(n_1056),
.B(n_1057),
.Y(n_11163)
);

AOI21xp5_ASAP7_75t_L g11164 ( 
.A1(n_10150),
.A2(n_1057),
.B(n_1058),
.Y(n_11164)
);

NOR2xp33_ASAP7_75t_L g11165 ( 
.A(n_10181),
.B(n_10172),
.Y(n_11165)
);

AOI21xp5_ASAP7_75t_L g11166 ( 
.A1(n_10170),
.A2(n_1058),
.B(n_1059),
.Y(n_11166)
);

O2A1O1Ixp33_ASAP7_75t_L g11167 ( 
.A1(n_10217),
.A2(n_1061),
.B(n_1059),
.C(n_1060),
.Y(n_11167)
);

NOR2xp67_ASAP7_75t_L g11168 ( 
.A(n_10167),
.B(n_1061),
.Y(n_11168)
);

AOI21xp5_ASAP7_75t_L g11169 ( 
.A1(n_9841),
.A2(n_1062),
.B(n_1063),
.Y(n_11169)
);

NAND2xp5_ASAP7_75t_L g11170 ( 
.A(n_10069),
.B(n_1062),
.Y(n_11170)
);

AOI21xp5_ASAP7_75t_L g11171 ( 
.A1(n_10061),
.A2(n_1063),
.B(n_1064),
.Y(n_11171)
);

AO22x1_ASAP7_75t_L g11172 ( 
.A1(n_10255),
.A2(n_1066),
.B1(n_1064),
.B2(n_1065),
.Y(n_11172)
);

NAND2xp5_ASAP7_75t_SL g11173 ( 
.A(n_10374),
.B(n_1065),
.Y(n_11173)
);

INVx5_ASAP7_75t_L g11174 ( 
.A(n_10411),
.Y(n_11174)
);

A2O1A1Ixp33_ASAP7_75t_L g11175 ( 
.A1(n_10272),
.A2(n_1068),
.B(n_1066),
.C(n_1067),
.Y(n_11175)
);

O2A1O1Ixp33_ASAP7_75t_L g11176 ( 
.A1(n_9965),
.A2(n_1070),
.B(n_1068),
.C(n_1069),
.Y(n_11176)
);

NAND2xp5_ASAP7_75t_L g11177 ( 
.A(n_10094),
.B(n_1070),
.Y(n_11177)
);

INVx1_ASAP7_75t_L g11178 ( 
.A(n_10400),
.Y(n_11178)
);

BUFx6f_ASAP7_75t_L g11179 ( 
.A(n_10215),
.Y(n_11179)
);

AND2x4_ASAP7_75t_L g11180 ( 
.A(n_10027),
.B(n_1071),
.Y(n_11180)
);

A2O1A1Ixp33_ASAP7_75t_L g11181 ( 
.A1(n_10273),
.A2(n_1073),
.B(n_1071),
.C(n_1072),
.Y(n_11181)
);

A2O1A1Ixp33_ASAP7_75t_L g11182 ( 
.A1(n_9993),
.A2(n_10016),
.B(n_10025),
.C(n_10019),
.Y(n_11182)
);

BUFx6f_ASAP7_75t_L g11183 ( 
.A(n_10226),
.Y(n_11183)
);

AOI21xp5_ASAP7_75t_L g11184 ( 
.A1(n_10064),
.A2(n_9964),
.B(n_10119),
.Y(n_11184)
);

BUFx4f_ASAP7_75t_SL g11185 ( 
.A(n_10068),
.Y(n_11185)
);

AOI21xp5_ASAP7_75t_L g11186 ( 
.A1(n_10123),
.A2(n_1072),
.B(n_1074),
.Y(n_11186)
);

NAND2xp5_ASAP7_75t_L g11187 ( 
.A(n_10029),
.B(n_1074),
.Y(n_11187)
);

BUFx12f_ASAP7_75t_L g11188 ( 
.A(n_10380),
.Y(n_11188)
);

NAND2xp5_ASAP7_75t_L g11189 ( 
.A(n_10032),
.B(n_1075),
.Y(n_11189)
);

AO21x1_ASAP7_75t_L g11190 ( 
.A1(n_10375),
.A2(n_1075),
.B(n_1076),
.Y(n_11190)
);

AND2x4_ASAP7_75t_L g11191 ( 
.A(n_10311),
.B(n_1076),
.Y(n_11191)
);

OAI21x1_ASAP7_75t_L g11192 ( 
.A1(n_10532),
.A2(n_1077),
.B(n_1078),
.Y(n_11192)
);

AO21x1_ASAP7_75t_L g11193 ( 
.A1(n_10043),
.A2(n_1078),
.B(n_1079),
.Y(n_11193)
);

AOI21xp5_ASAP7_75t_L g11194 ( 
.A1(n_10213),
.A2(n_1079),
.B(n_1080),
.Y(n_11194)
);

INVx2_ASAP7_75t_L g11195 ( 
.A(n_10040),
.Y(n_11195)
);

NOR2xp67_ASAP7_75t_SL g11196 ( 
.A(n_9870),
.B(n_1080),
.Y(n_11196)
);

BUFx6f_ASAP7_75t_L g11197 ( 
.A(n_10098),
.Y(n_11197)
);

OAI22xp5_ASAP7_75t_L g11198 ( 
.A1(n_9899),
.A2(n_1084),
.B1(n_1082),
.B2(n_1083),
.Y(n_11198)
);

AND2x4_ASAP7_75t_L g11199 ( 
.A(n_10168),
.B(n_1083),
.Y(n_11199)
);

NAND2xp5_ASAP7_75t_L g11200 ( 
.A(n_10047),
.B(n_1084),
.Y(n_11200)
);

NAND3xp33_ASAP7_75t_L g11201 ( 
.A(n_10052),
.B(n_10053),
.C(n_10066),
.Y(n_11201)
);

AOI21xp5_ASAP7_75t_L g11202 ( 
.A1(n_10288),
.A2(n_1085),
.B(n_1086),
.Y(n_11202)
);

NOR2xp33_ASAP7_75t_L g11203 ( 
.A(n_10386),
.B(n_1085),
.Y(n_11203)
);

NAND3xp33_ASAP7_75t_L g11204 ( 
.A(n_10104),
.B(n_1086),
.C(n_1087),
.Y(n_11204)
);

CKINVDCx16_ASAP7_75t_R g11205 ( 
.A(n_10377),
.Y(n_11205)
);

INVxp67_ASAP7_75t_SL g11206 ( 
.A(n_10054),
.Y(n_11206)
);

HB1xp67_ASAP7_75t_L g11207 ( 
.A(n_10023),
.Y(n_11207)
);

INVx5_ASAP7_75t_L g11208 ( 
.A(n_10382),
.Y(n_11208)
);

NAND2xp5_ASAP7_75t_SL g11209 ( 
.A(n_10118),
.B(n_1087),
.Y(n_11209)
);

NOR2xp33_ASAP7_75t_L g11210 ( 
.A(n_10266),
.B(n_1088),
.Y(n_11210)
);

AOI33xp33_ASAP7_75t_L g11211 ( 
.A1(n_10268),
.A2(n_1091),
.A3(n_1093),
.B1(n_1089),
.B2(n_1090),
.B3(n_1092),
.Y(n_11211)
);

HB1xp67_ASAP7_75t_L g11212 ( 
.A(n_10166),
.Y(n_11212)
);

NOR2xp33_ASAP7_75t_L g11213 ( 
.A(n_10121),
.B(n_1089),
.Y(n_11213)
);

NAND2xp5_ASAP7_75t_L g11214 ( 
.A(n_10125),
.B(n_1090),
.Y(n_11214)
);

AOI21xp5_ASAP7_75t_L g11215 ( 
.A1(n_10294),
.A2(n_10308),
.B(n_10303),
.Y(n_11215)
);

NAND2xp5_ASAP7_75t_L g11216 ( 
.A(n_10131),
.B(n_10137),
.Y(n_11216)
);

AOI22xp33_ASAP7_75t_L g11217 ( 
.A1(n_9909),
.A2(n_1094),
.B1(n_1092),
.B2(n_1093),
.Y(n_11217)
);

NAND2xp5_ASAP7_75t_L g11218 ( 
.A(n_10292),
.B(n_1094),
.Y(n_11218)
);

BUFx2_ASAP7_75t_L g11219 ( 
.A(n_10151),
.Y(n_11219)
);

OAI22xp5_ASAP7_75t_L g11220 ( 
.A1(n_9885),
.A2(n_1097),
.B1(n_1095),
.B2(n_1096),
.Y(n_11220)
);

NAND2xp5_ASAP7_75t_L g11221 ( 
.A(n_10223),
.B(n_1095),
.Y(n_11221)
);

BUFx2_ASAP7_75t_L g11222 ( 
.A(n_10327),
.Y(n_11222)
);

NAND2xp5_ASAP7_75t_SL g11223 ( 
.A(n_10178),
.B(n_1096),
.Y(n_11223)
);

NOR3xp33_ASAP7_75t_SL g11224 ( 
.A(n_10234),
.B(n_1097),
.C(n_1098),
.Y(n_11224)
);

NAND3xp33_ASAP7_75t_L g11225 ( 
.A(n_10180),
.B(n_10190),
.C(n_10183),
.Y(n_11225)
);

AND2x4_ASAP7_75t_L g11226 ( 
.A(n_10329),
.B(n_1098),
.Y(n_11226)
);

OAI22xp5_ASAP7_75t_L g11227 ( 
.A1(n_9857),
.A2(n_1101),
.B1(n_1099),
.B2(n_1100),
.Y(n_11227)
);

NAND2xp5_ASAP7_75t_SL g11228 ( 
.A(n_10197),
.B(n_1100),
.Y(n_11228)
);

INVx1_ASAP7_75t_L g11229 ( 
.A(n_10309),
.Y(n_11229)
);

INVx1_ASAP7_75t_L g11230 ( 
.A(n_10326),
.Y(n_11230)
);

O2A1O1Ixp33_ASAP7_75t_L g11231 ( 
.A1(n_10034),
.A2(n_10152),
.B(n_9896),
.C(n_10216),
.Y(n_11231)
);

NAND2xp33_ASAP7_75t_R g11232 ( 
.A(n_10218),
.B(n_1101),
.Y(n_11232)
);

AOI21xp5_ASAP7_75t_L g11233 ( 
.A1(n_9858),
.A2(n_1102),
.B(n_1103),
.Y(n_11233)
);

CKINVDCx20_ASAP7_75t_R g11234 ( 
.A(n_10335),
.Y(n_11234)
);

A2O1A1Ixp33_ASAP7_75t_L g11235 ( 
.A1(n_10348),
.A2(n_10360),
.B(n_10370),
.C(n_10365),
.Y(n_11235)
);

A2O1A1Ixp33_ASAP7_75t_L g11236 ( 
.A1(n_10371),
.A2(n_1107),
.B(n_1105),
.C(n_1106),
.Y(n_11236)
);

OAI22xp5_ASAP7_75t_L g11237 ( 
.A1(n_9868),
.A2(n_1108),
.B1(n_1105),
.B2(n_1106),
.Y(n_11237)
);

OAI22xp5_ASAP7_75t_L g11238 ( 
.A1(n_10423),
.A2(n_1110),
.B1(n_1108),
.B2(n_1109),
.Y(n_11238)
);

INVx4_ASAP7_75t_L g11239 ( 
.A(n_10205),
.Y(n_11239)
);

NAND2xp5_ASAP7_75t_L g11240 ( 
.A(n_10432),
.B(n_1109),
.Y(n_11240)
);

A2O1A1Ixp33_ASAP7_75t_L g11241 ( 
.A1(n_9966),
.A2(n_1113),
.B(n_1111),
.C(n_1112),
.Y(n_11241)
);

OAI22xp5_ASAP7_75t_L g11242 ( 
.A1(n_10423),
.A2(n_1114),
.B1(n_1112),
.B2(n_1113),
.Y(n_11242)
);

AOI21xp5_ASAP7_75t_L g11243 ( 
.A1(n_9912),
.A2(n_1114),
.B(n_1115),
.Y(n_11243)
);

AOI21x1_ASAP7_75t_L g11244 ( 
.A1(n_10078),
.A2(n_1115),
.B(n_1116),
.Y(n_11244)
);

AOI21xp5_ASAP7_75t_L g11245 ( 
.A1(n_9912),
.A2(n_1116),
.B(n_1117),
.Y(n_11245)
);

AOI21xp5_ASAP7_75t_L g11246 ( 
.A1(n_9912),
.A2(n_1117),
.B(n_1118),
.Y(n_11246)
);

BUFx3_ASAP7_75t_L g11247 ( 
.A(n_10230),
.Y(n_11247)
);

CKINVDCx5p33_ASAP7_75t_R g11248 ( 
.A(n_10051),
.Y(n_11248)
);

BUFx4_ASAP7_75t_SL g11249 ( 
.A(n_10420),
.Y(n_11249)
);

INVx1_ASAP7_75t_SL g11250 ( 
.A(n_10230),
.Y(n_11250)
);

AOI22xp33_ASAP7_75t_L g11251 ( 
.A1(n_9950),
.A2(n_1122),
.B1(n_1118),
.B2(n_1121),
.Y(n_11251)
);

NOR2xp33_ASAP7_75t_L g11252 ( 
.A(n_10281),
.B(n_1121),
.Y(n_11252)
);

AOI21xp5_ASAP7_75t_L g11253 ( 
.A1(n_9912),
.A2(n_1122),
.B(n_1123),
.Y(n_11253)
);

INVx2_ASAP7_75t_L g11254 ( 
.A(n_10235),
.Y(n_11254)
);

NAND3xp33_ASAP7_75t_L g11255 ( 
.A(n_10423),
.B(n_1123),
.C(n_1124),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_10010),
.Y(n_11256)
);

OAI22xp5_ASAP7_75t_L g11257 ( 
.A1(n_10423),
.A2(n_1126),
.B1(n_1124),
.B2(n_1125),
.Y(n_11257)
);

AOI21xp5_ASAP7_75t_L g11258 ( 
.A1(n_9912),
.A2(n_1125),
.B(n_1126),
.Y(n_11258)
);

A2O1A1Ixp33_ASAP7_75t_L g11259 ( 
.A1(n_9966),
.A2(n_1129),
.B(n_1127),
.C(n_1128),
.Y(n_11259)
);

NAND2xp5_ASAP7_75t_SL g11260 ( 
.A(n_9949),
.B(n_1127),
.Y(n_11260)
);

OAI221xp5_ASAP7_75t_L g11261 ( 
.A1(n_9883),
.A2(n_1131),
.B1(n_1128),
.B2(n_1130),
.C(n_1132),
.Y(n_11261)
);

O2A1O1Ixp33_ASAP7_75t_L g11262 ( 
.A1(n_9966),
.A2(n_1133),
.B(n_1130),
.C(n_1131),
.Y(n_11262)
);

CKINVDCx16_ASAP7_75t_R g11263 ( 
.A(n_10051),
.Y(n_11263)
);

BUFx6f_ASAP7_75t_L g11264 ( 
.A(n_10114),
.Y(n_11264)
);

INVx2_ASAP7_75t_L g11265 ( 
.A(n_10235),
.Y(n_11265)
);

AOI21xp5_ASAP7_75t_L g11266 ( 
.A1(n_9912),
.A2(n_1133),
.B(n_1134),
.Y(n_11266)
);

NAND2xp5_ASAP7_75t_L g11267 ( 
.A(n_10432),
.B(n_1134),
.Y(n_11267)
);

NAND2xp5_ASAP7_75t_L g11268 ( 
.A(n_10432),
.B(n_1135),
.Y(n_11268)
);

AOI21xp5_ASAP7_75t_L g11269 ( 
.A1(n_9912),
.A2(n_1136),
.B(n_1137),
.Y(n_11269)
);

AOI21xp5_ASAP7_75t_L g11270 ( 
.A1(n_9912),
.A2(n_1138),
.B(n_1139),
.Y(n_11270)
);

OAI21xp33_ASAP7_75t_SL g11271 ( 
.A1(n_10423),
.A2(n_1139),
.B(n_1140),
.Y(n_11271)
);

NAND2xp5_ASAP7_75t_L g11272 ( 
.A(n_10432),
.B(n_1140),
.Y(n_11272)
);

A2O1A1Ixp33_ASAP7_75t_L g11273 ( 
.A1(n_9966),
.A2(n_1143),
.B(n_1141),
.C(n_1142),
.Y(n_11273)
);

BUFx6f_ASAP7_75t_L g11274 ( 
.A(n_10114),
.Y(n_11274)
);

OAI22xp5_ASAP7_75t_L g11275 ( 
.A1(n_10423),
.A2(n_1144),
.B1(n_1142),
.B2(n_1143),
.Y(n_11275)
);

BUFx8_ASAP7_75t_L g11276 ( 
.A(n_10051),
.Y(n_11276)
);

O2A1O1Ixp33_ASAP7_75t_L g11277 ( 
.A1(n_9966),
.A2(n_1146),
.B(n_1144),
.C(n_1145),
.Y(n_11277)
);

NAND2xp5_ASAP7_75t_SL g11278 ( 
.A(n_9949),
.B(n_1145),
.Y(n_11278)
);

CKINVDCx14_ASAP7_75t_R g11279 ( 
.A(n_10051),
.Y(n_11279)
);

CKINVDCx6p67_ASAP7_75t_R g11280 ( 
.A(n_10087),
.Y(n_11280)
);

NOR2xp33_ASAP7_75t_L g11281 ( 
.A(n_10281),
.B(n_1146),
.Y(n_11281)
);

NAND2xp5_ASAP7_75t_SL g11282 ( 
.A(n_9949),
.B(n_1147),
.Y(n_11282)
);

AND2x4_ASAP7_75t_L g11283 ( 
.A(n_10252),
.B(n_1148),
.Y(n_11283)
);

BUFx3_ASAP7_75t_L g11284 ( 
.A(n_10230),
.Y(n_11284)
);

NAND2xp5_ASAP7_75t_L g11285 ( 
.A(n_10432),
.B(n_1148),
.Y(n_11285)
);

INVx3_ASAP7_75t_L g11286 ( 
.A(n_9980),
.Y(n_11286)
);

INVx1_ASAP7_75t_L g11287 ( 
.A(n_10010),
.Y(n_11287)
);

INVx2_ASAP7_75t_L g11288 ( 
.A(n_10235),
.Y(n_11288)
);

OAI22xp5_ASAP7_75t_L g11289 ( 
.A1(n_10566),
.A2(n_1151),
.B1(n_1149),
.B2(n_1150),
.Y(n_11289)
);

AOI21xp5_ASAP7_75t_L g11290 ( 
.A1(n_10586),
.A2(n_1150),
.B(n_1151),
.Y(n_11290)
);

NOR2x1_ASAP7_75t_L g11291 ( 
.A(n_10783),
.B(n_1152),
.Y(n_11291)
);

OAI21x1_ASAP7_75t_L g11292 ( 
.A1(n_11122),
.A2(n_1152),
.B(n_1153),
.Y(n_11292)
);

OAI21x1_ASAP7_75t_L g11293 ( 
.A1(n_11127),
.A2(n_1153),
.B(n_1154),
.Y(n_11293)
);

O2A1O1Ixp5_ASAP7_75t_L g11294 ( 
.A1(n_10719),
.A2(n_1156),
.B(n_1154),
.C(n_1155),
.Y(n_11294)
);

AOI21xp5_ASAP7_75t_L g11295 ( 
.A1(n_11215),
.A2(n_1155),
.B(n_1157),
.Y(n_11295)
);

OAI21x1_ASAP7_75t_L g11296 ( 
.A1(n_11107),
.A2(n_1157),
.B(n_1158),
.Y(n_11296)
);

BUFx12f_ASAP7_75t_L g11297 ( 
.A(n_11276),
.Y(n_11297)
);

CKINVDCx11_ASAP7_75t_R g11298 ( 
.A(n_11280),
.Y(n_11298)
);

OA21x2_ASAP7_75t_L g11299 ( 
.A1(n_10863),
.A2(n_1158),
.B(n_1159),
.Y(n_11299)
);

NAND2xp5_ASAP7_75t_L g11300 ( 
.A(n_10654),
.B(n_1159),
.Y(n_11300)
);

AO31x2_ASAP7_75t_L g11301 ( 
.A1(n_11152),
.A2(n_1162),
.A3(n_1160),
.B(n_1161),
.Y(n_11301)
);

OAI21x1_ASAP7_75t_L g11302 ( 
.A1(n_10973),
.A2(n_1160),
.B(n_1161),
.Y(n_11302)
);

O2A1O1Ixp5_ASAP7_75t_SL g11303 ( 
.A1(n_11047),
.A2(n_1165),
.B(n_1162),
.C(n_1163),
.Y(n_11303)
);

AOI22xp33_ASAP7_75t_L g11304 ( 
.A1(n_11234),
.A2(n_1167),
.B1(n_1163),
.B2(n_1166),
.Y(n_11304)
);

NAND2xp5_ASAP7_75t_L g11305 ( 
.A(n_10615),
.B(n_1167),
.Y(n_11305)
);

NAND2xp5_ASAP7_75t_L g11306 ( 
.A(n_10627),
.B(n_1168),
.Y(n_11306)
);

BUFx3_ASAP7_75t_L g11307 ( 
.A(n_10612),
.Y(n_11307)
);

AO21x2_ASAP7_75t_L g11308 ( 
.A1(n_10903),
.A2(n_1168),
.B(n_1169),
.Y(n_11308)
);

AOI21xp5_ASAP7_75t_L g11309 ( 
.A1(n_11052),
.A2(n_1169),
.B(n_1170),
.Y(n_11309)
);

NAND3xp33_ASAP7_75t_L g11310 ( 
.A(n_11255),
.B(n_1170),
.C(n_1171),
.Y(n_11310)
);

AOI21xp5_ASAP7_75t_SL g11311 ( 
.A1(n_10585),
.A2(n_1171),
.B(n_1172),
.Y(n_11311)
);

AOI31xp67_ASAP7_75t_L g11312 ( 
.A1(n_11161),
.A2(n_1174),
.A3(n_1172),
.B(n_1173),
.Y(n_11312)
);

INVx2_ASAP7_75t_L g11313 ( 
.A(n_10965),
.Y(n_11313)
);

OA22x2_ASAP7_75t_L g11314 ( 
.A1(n_10698),
.A2(n_1175),
.B1(n_1173),
.B2(n_1174),
.Y(n_11314)
);

AOI21xp5_ASAP7_75t_L g11315 ( 
.A1(n_10703),
.A2(n_10858),
.B(n_10644),
.Y(n_11315)
);

NAND2xp5_ASAP7_75t_L g11316 ( 
.A(n_10569),
.B(n_1176),
.Y(n_11316)
);

BUFx2_ASAP7_75t_L g11317 ( 
.A(n_10717),
.Y(n_11317)
);

AND2x2_ASAP7_75t_L g11318 ( 
.A(n_10708),
.B(n_1176),
.Y(n_11318)
);

NAND2xp5_ASAP7_75t_L g11319 ( 
.A(n_11256),
.B(n_11287),
.Y(n_11319)
);

OAI21x1_ASAP7_75t_L g11320 ( 
.A1(n_10608),
.A2(n_1177),
.B(n_1178),
.Y(n_11320)
);

OAI21x1_ASAP7_75t_L g11321 ( 
.A1(n_11114),
.A2(n_1178),
.B(n_1179),
.Y(n_11321)
);

INVx1_ASAP7_75t_SL g11322 ( 
.A(n_10818),
.Y(n_11322)
);

A2O1A1Ixp33_ASAP7_75t_L g11323 ( 
.A1(n_10602),
.A2(n_1181),
.B(n_1179),
.C(n_1180),
.Y(n_11323)
);

OAI22xp5_ASAP7_75t_L g11324 ( 
.A1(n_11205),
.A2(n_1182),
.B1(n_1180),
.B2(n_1181),
.Y(n_11324)
);

INVx2_ASAP7_75t_L g11325 ( 
.A(n_10965),
.Y(n_11325)
);

NAND2xp5_ASAP7_75t_L g11326 ( 
.A(n_10781),
.B(n_1182),
.Y(n_11326)
);

NAND2xp5_ASAP7_75t_L g11327 ( 
.A(n_10587),
.B(n_1183),
.Y(n_11327)
);

OAI22xp5_ASAP7_75t_SL g11328 ( 
.A1(n_10628),
.A2(n_1185),
.B1(n_1183),
.B2(n_1184),
.Y(n_11328)
);

AO31x2_ASAP7_75t_L g11329 ( 
.A1(n_11115),
.A2(n_1186),
.A3(n_1184),
.B(n_1185),
.Y(n_11329)
);

OAI21x1_ASAP7_75t_L g11330 ( 
.A1(n_11036),
.A2(n_1186),
.B(n_1187),
.Y(n_11330)
);

AO31x2_ASAP7_75t_L g11331 ( 
.A1(n_11178),
.A2(n_1190),
.A3(n_1188),
.B(n_1189),
.Y(n_11331)
);

OAI21xp5_ASAP7_75t_L g11332 ( 
.A1(n_10575),
.A2(n_1189),
.B(n_1190),
.Y(n_11332)
);

AND2x6_ASAP7_75t_L g11333 ( 
.A(n_11229),
.B(n_1191),
.Y(n_11333)
);

INVx2_ASAP7_75t_L g11334 ( 
.A(n_10972),
.Y(n_11334)
);

BUFx6f_ASAP7_75t_L g11335 ( 
.A(n_10804),
.Y(n_11335)
);

OAI22xp5_ASAP7_75t_L g11336 ( 
.A1(n_11014),
.A2(n_1193),
.B1(n_1191),
.B2(n_1192),
.Y(n_11336)
);

INVxp67_ASAP7_75t_L g11337 ( 
.A(n_10578),
.Y(n_11337)
);

OAI21x1_ASAP7_75t_L g11338 ( 
.A1(n_11206),
.A2(n_1192),
.B(n_1193),
.Y(n_11338)
);

HB1xp67_ASAP7_75t_L g11339 ( 
.A(n_10735),
.Y(n_11339)
);

OAI21x1_ASAP7_75t_L g11340 ( 
.A1(n_10570),
.A2(n_1194),
.B(n_1195),
.Y(n_11340)
);

NAND2xp33_ASAP7_75t_L g11341 ( 
.A(n_10819),
.B(n_1196),
.Y(n_11341)
);

OAI21x1_ASAP7_75t_L g11342 ( 
.A1(n_11244),
.A2(n_1196),
.B(n_1197),
.Y(n_11342)
);

O2A1O1Ixp33_ASAP7_75t_L g11343 ( 
.A1(n_11123),
.A2(n_1199),
.B(n_1197),
.C(n_1198),
.Y(n_11343)
);

NAND2xp5_ASAP7_75t_L g11344 ( 
.A(n_10892),
.B(n_10945),
.Y(n_11344)
);

OAI21xp5_ASAP7_75t_L g11345 ( 
.A1(n_11243),
.A2(n_1198),
.B(n_1200),
.Y(n_11345)
);

AND2x2_ASAP7_75t_L g11346 ( 
.A(n_11061),
.B(n_1200),
.Y(n_11346)
);

BUFx2_ASAP7_75t_L g11347 ( 
.A(n_10847),
.Y(n_11347)
);

INVx2_ASAP7_75t_SL g11348 ( 
.A(n_11247),
.Y(n_11348)
);

OAI21x1_ASAP7_75t_L g11349 ( 
.A1(n_11195),
.A2(n_1201),
.B(n_1202),
.Y(n_11349)
);

OAI21x1_ASAP7_75t_L g11350 ( 
.A1(n_10582),
.A2(n_1201),
.B(n_1202),
.Y(n_11350)
);

AND2x4_ASAP7_75t_L g11351 ( 
.A(n_10748),
.B(n_1203),
.Y(n_11351)
);

AO21x1_ASAP7_75t_L g11352 ( 
.A1(n_10710),
.A2(n_1204),
.B(n_1205),
.Y(n_11352)
);

AO21x1_ASAP7_75t_L g11353 ( 
.A1(n_10593),
.A2(n_1205),
.B(n_1206),
.Y(n_11353)
);

INVx1_ASAP7_75t_L g11354 ( 
.A(n_10780),
.Y(n_11354)
);

NAND2x1p5_ASAP7_75t_L g11355 ( 
.A(n_10628),
.B(n_1206),
.Y(n_11355)
);

NAND2xp5_ASAP7_75t_L g11356 ( 
.A(n_11125),
.B(n_1207),
.Y(n_11356)
);

NAND2xp5_ASAP7_75t_SL g11357 ( 
.A(n_11060),
.B(n_1207),
.Y(n_11357)
);

OAI21x1_ASAP7_75t_L g11358 ( 
.A1(n_10880),
.A2(n_1208),
.B(n_1209),
.Y(n_11358)
);

AO31x2_ASAP7_75t_L g11359 ( 
.A1(n_10647),
.A2(n_11222),
.A3(n_11119),
.B(n_11105),
.Y(n_11359)
);

INVx2_ASAP7_75t_L g11360 ( 
.A(n_10972),
.Y(n_11360)
);

AOI21xp5_ASAP7_75t_L g11361 ( 
.A1(n_11260),
.A2(n_1208),
.B(n_1210),
.Y(n_11361)
);

OAI21x1_ASAP7_75t_L g11362 ( 
.A1(n_11120),
.A2(n_1210),
.B(n_1211),
.Y(n_11362)
);

AO21x2_ASAP7_75t_L g11363 ( 
.A1(n_10756),
.A2(n_1211),
.B(n_1212),
.Y(n_11363)
);

AOI21xp5_ASAP7_75t_L g11364 ( 
.A1(n_11278),
.A2(n_1212),
.B(n_1213),
.Y(n_11364)
);

OAI21xp5_ASAP7_75t_L g11365 ( 
.A1(n_11245),
.A2(n_1214),
.B(n_1215),
.Y(n_11365)
);

NOR4xp25_ASAP7_75t_L g11366 ( 
.A(n_11106),
.B(n_1217),
.C(n_1214),
.D(n_1216),
.Y(n_11366)
);

BUFx6f_ASAP7_75t_L g11367 ( 
.A(n_10804),
.Y(n_11367)
);

OAI21xp5_ASAP7_75t_L g11368 ( 
.A1(n_11246),
.A2(n_1217),
.B(n_1218),
.Y(n_11368)
);

O2A1O1Ixp33_ASAP7_75t_L g11369 ( 
.A1(n_10643),
.A2(n_1222),
.B(n_1219),
.C(n_1220),
.Y(n_11369)
);

OAI21xp5_ASAP7_75t_L g11370 ( 
.A1(n_11253),
.A2(n_1220),
.B(n_1222),
.Y(n_11370)
);

AND2x2_ASAP7_75t_L g11371 ( 
.A(n_11060),
.B(n_1223),
.Y(n_11371)
);

INVx2_ASAP7_75t_L g11372 ( 
.A(n_11000),
.Y(n_11372)
);

NOR2xp67_ASAP7_75t_L g11373 ( 
.A(n_10702),
.B(n_10787),
.Y(n_11373)
);

OAI21x1_ASAP7_75t_L g11374 ( 
.A1(n_10695),
.A2(n_1224),
.B(n_1225),
.Y(n_11374)
);

NAND2xp5_ASAP7_75t_L g11375 ( 
.A(n_10947),
.B(n_1224),
.Y(n_11375)
);

AOI21xp33_ASAP7_75t_L g11376 ( 
.A1(n_11232),
.A2(n_1225),
.B(n_1226),
.Y(n_11376)
);

AOI21xp5_ASAP7_75t_L g11377 ( 
.A1(n_11282),
.A2(n_1226),
.B(n_1227),
.Y(n_11377)
);

NAND2xp33_ASAP7_75t_L g11378 ( 
.A(n_10633),
.B(n_10955),
.Y(n_11378)
);

NAND2xp5_ASAP7_75t_SL g11379 ( 
.A(n_11162),
.B(n_1227),
.Y(n_11379)
);

BUFx3_ASAP7_75t_L g11380 ( 
.A(n_10669),
.Y(n_11380)
);

INVx1_ASAP7_75t_L g11381 ( 
.A(n_10766),
.Y(n_11381)
);

AOI21x1_ASAP7_75t_L g11382 ( 
.A1(n_11212),
.A2(n_1228),
.B(n_1229),
.Y(n_11382)
);

NAND2xp5_ASAP7_75t_SL g11383 ( 
.A(n_11162),
.B(n_1228),
.Y(n_11383)
);

OAI21x1_ASAP7_75t_SL g11384 ( 
.A1(n_11258),
.A2(n_1229),
.B(n_1230),
.Y(n_11384)
);

AND2x2_ASAP7_75t_L g11385 ( 
.A(n_10986),
.B(n_10968),
.Y(n_11385)
);

AOI221xp5_ASAP7_75t_L g11386 ( 
.A1(n_11210),
.A2(n_1232),
.B1(n_1230),
.B2(n_1231),
.C(n_1233),
.Y(n_11386)
);

AND2x2_ASAP7_75t_L g11387 ( 
.A(n_11057),
.B(n_1231),
.Y(n_11387)
);

NAND2xp5_ASAP7_75t_L g11388 ( 
.A(n_11004),
.B(n_1232),
.Y(n_11388)
);

OAI21x1_ASAP7_75t_L g11389 ( 
.A1(n_11230),
.A2(n_1233),
.B(n_1234),
.Y(n_11389)
);

NAND2xp5_ASAP7_75t_L g11390 ( 
.A(n_10827),
.B(n_1234),
.Y(n_11390)
);

AOI21x1_ASAP7_75t_L g11391 ( 
.A1(n_11156),
.A2(n_1235),
.B(n_1236),
.Y(n_11391)
);

CKINVDCx11_ASAP7_75t_R g11392 ( 
.A(n_10832),
.Y(n_11392)
);

O2A1O1Ixp5_ASAP7_75t_L g11393 ( 
.A1(n_11031),
.A2(n_1238),
.B(n_1235),
.C(n_1236),
.Y(n_11393)
);

NAND2x1p5_ASAP7_75t_L g11394 ( 
.A(n_10652),
.B(n_1238),
.Y(n_11394)
);

AO22x2_ASAP7_75t_L g11395 ( 
.A1(n_10799),
.A2(n_1241),
.B1(n_1239),
.B2(n_1240),
.Y(n_11395)
);

OAI21xp5_ASAP7_75t_L g11396 ( 
.A1(n_11266),
.A2(n_1239),
.B(n_1240),
.Y(n_11396)
);

AOI21x1_ASAP7_75t_SL g11397 ( 
.A1(n_11216),
.A2(n_1241),
.B(n_1242),
.Y(n_11397)
);

OAI21xp5_ASAP7_75t_L g11398 ( 
.A1(n_11269),
.A2(n_1242),
.B(n_1243),
.Y(n_11398)
);

AOI21x1_ASAP7_75t_SL g11399 ( 
.A1(n_11285),
.A2(n_1243),
.B(n_1244),
.Y(n_11399)
);

OAI21x1_ASAP7_75t_L g11400 ( 
.A1(n_11184),
.A2(n_1244),
.B(n_1245),
.Y(n_11400)
);

AOI21xp5_ASAP7_75t_L g11401 ( 
.A1(n_10730),
.A2(n_1246),
.B(n_1247),
.Y(n_11401)
);

INVx2_ASAP7_75t_L g11402 ( 
.A(n_11000),
.Y(n_11402)
);

OAI21x1_ASAP7_75t_L g11403 ( 
.A1(n_10852),
.A2(n_1246),
.B(n_1247),
.Y(n_11403)
);

BUFx6f_ASAP7_75t_L g11404 ( 
.A(n_10691),
.Y(n_11404)
);

AOI22xp5_ASAP7_75t_L g11405 ( 
.A1(n_10686),
.A2(n_1250),
.B1(n_1248),
.B2(n_1249),
.Y(n_11405)
);

NAND2xp5_ASAP7_75t_L g11406 ( 
.A(n_11074),
.B(n_1248),
.Y(n_11406)
);

OAI21x1_ASAP7_75t_L g11407 ( 
.A1(n_11207),
.A2(n_1250),
.B(n_1251),
.Y(n_11407)
);

OAI21x1_ASAP7_75t_L g11408 ( 
.A1(n_10577),
.A2(n_11267),
.B(n_11240),
.Y(n_11408)
);

OAI21x1_ASAP7_75t_L g11409 ( 
.A1(n_11268),
.A2(n_1252),
.B(n_1253),
.Y(n_11409)
);

A2O1A1Ixp33_ASAP7_75t_L g11410 ( 
.A1(n_10727),
.A2(n_1254),
.B(n_1252),
.C(n_1253),
.Y(n_11410)
);

BUFx6f_ASAP7_75t_L g11411 ( 
.A(n_10691),
.Y(n_11411)
);

OAI21x1_ASAP7_75t_L g11412 ( 
.A1(n_11272),
.A2(n_1254),
.B(n_1255),
.Y(n_11412)
);

INVx2_ASAP7_75t_L g11413 ( 
.A(n_11001),
.Y(n_11413)
);

AO21x2_ASAP7_75t_L g11414 ( 
.A1(n_11111),
.A2(n_1255),
.B(n_1256),
.Y(n_11414)
);

OAI21x1_ASAP7_75t_SL g11415 ( 
.A1(n_11270),
.A2(n_1256),
.B(n_1257),
.Y(n_11415)
);

NAND2x1p5_ASAP7_75t_L g11416 ( 
.A(n_10652),
.B(n_1257),
.Y(n_11416)
);

NAND3xp33_ASAP7_75t_SL g11417 ( 
.A(n_10977),
.B(n_1258),
.C(n_1259),
.Y(n_11417)
);

NAND2xp5_ASAP7_75t_L g11418 ( 
.A(n_11096),
.B(n_1259),
.Y(n_11418)
);

BUFx2_ASAP7_75t_L g11419 ( 
.A(n_10853),
.Y(n_11419)
);

BUFx3_ASAP7_75t_L g11420 ( 
.A(n_10588),
.Y(n_11420)
);

NAND2xp5_ASAP7_75t_L g11421 ( 
.A(n_10855),
.B(n_1260),
.Y(n_11421)
);

INVx1_ASAP7_75t_L g11422 ( 
.A(n_10773),
.Y(n_11422)
);

OAI21xp5_ASAP7_75t_L g11423 ( 
.A1(n_10731),
.A2(n_1260),
.B(n_1262),
.Y(n_11423)
);

OAI21x1_ASAP7_75t_L g11424 ( 
.A1(n_10813),
.A2(n_1263),
.B(n_1264),
.Y(n_11424)
);

OAI21x1_ASAP7_75t_SL g11425 ( 
.A1(n_10692),
.A2(n_1263),
.B(n_1265),
.Y(n_11425)
);

NAND3xp33_ASAP7_75t_L g11426 ( 
.A(n_11201),
.B(n_1265),
.C(n_1266),
.Y(n_11426)
);

OAI21xp5_ASAP7_75t_L g11427 ( 
.A1(n_10676),
.A2(n_1266),
.B(n_1267),
.Y(n_11427)
);

AND2x2_ASAP7_75t_L g11428 ( 
.A(n_10885),
.B(n_1267),
.Y(n_11428)
);

NAND2xp5_ASAP7_75t_L g11429 ( 
.A(n_11128),
.B(n_1268),
.Y(n_11429)
);

A2O1A1Ixp33_ASAP7_75t_L g11430 ( 
.A1(n_10737),
.A2(n_1270),
.B(n_1268),
.C(n_1269),
.Y(n_11430)
);

OAI21x1_ASAP7_75t_L g11431 ( 
.A1(n_10878),
.A2(n_1269),
.B(n_1271),
.Y(n_11431)
);

INVx1_ASAP7_75t_L g11432 ( 
.A(n_10775),
.Y(n_11432)
);

OAI22x1_ASAP7_75t_L g11433 ( 
.A1(n_10702),
.A2(n_1273),
.B1(n_1271),
.B2(n_1272),
.Y(n_11433)
);

BUFx3_ASAP7_75t_L g11434 ( 
.A(n_11284),
.Y(n_11434)
);

OAI21x1_ASAP7_75t_L g11435 ( 
.A1(n_10890),
.A2(n_1272),
.B(n_1273),
.Y(n_11435)
);

OAI21x1_ASAP7_75t_L g11436 ( 
.A1(n_10922),
.A2(n_1274),
.B(n_1275),
.Y(n_11436)
);

AND2x4_ASAP7_75t_L g11437 ( 
.A(n_10666),
.B(n_1275),
.Y(n_11437)
);

NAND2xp5_ASAP7_75t_L g11438 ( 
.A(n_11131),
.B(n_1276),
.Y(n_11438)
);

OAI21xp5_ASAP7_75t_L g11439 ( 
.A1(n_11241),
.A2(n_1276),
.B(n_1277),
.Y(n_11439)
);

NAND2xp5_ASAP7_75t_L g11440 ( 
.A(n_11133),
.B(n_1277),
.Y(n_11440)
);

NAND2xp5_ASAP7_75t_L g11441 ( 
.A(n_11148),
.B(n_1278),
.Y(n_11441)
);

NAND2xp5_ASAP7_75t_SL g11442 ( 
.A(n_10967),
.B(n_1278),
.Y(n_11442)
);

AOI21xp5_ASAP7_75t_L g11443 ( 
.A1(n_11143),
.A2(n_1279),
.B(n_1280),
.Y(n_11443)
);

OA22x2_ASAP7_75t_L g11444 ( 
.A1(n_10585),
.A2(n_11147),
.B1(n_11091),
.B2(n_10596),
.Y(n_11444)
);

INVx4_ASAP7_75t_L g11445 ( 
.A(n_10761),
.Y(n_11445)
);

INVx2_ASAP7_75t_L g11446 ( 
.A(n_11001),
.Y(n_11446)
);

OAI21x1_ASAP7_75t_L g11447 ( 
.A1(n_10980),
.A2(n_1279),
.B(n_1280),
.Y(n_11447)
);

INVx1_ASAP7_75t_L g11448 ( 
.A(n_10685),
.Y(n_11448)
);

NAND2xp5_ASAP7_75t_L g11449 ( 
.A(n_11149),
.B(n_1281),
.Y(n_11449)
);

BUFx2_ASAP7_75t_L g11450 ( 
.A(n_10797),
.Y(n_11450)
);

OAI21x1_ASAP7_75t_L g11451 ( 
.A1(n_11192),
.A2(n_1281),
.B(n_1282),
.Y(n_11451)
);

AO31x2_ASAP7_75t_L g11452 ( 
.A1(n_11219),
.A2(n_1284),
.A3(n_1282),
.B(n_1283),
.Y(n_11452)
);

INVx2_ASAP7_75t_L g11453 ( 
.A(n_10701),
.Y(n_11453)
);

AO21x2_ASAP7_75t_L g11454 ( 
.A1(n_10771),
.A2(n_1283),
.B(n_1284),
.Y(n_11454)
);

AO31x2_ASAP7_75t_L g11455 ( 
.A1(n_11190),
.A2(n_11193),
.A3(n_11099),
.B(n_11100),
.Y(n_11455)
);

OAI21xp5_ASAP7_75t_L g11456 ( 
.A1(n_11259),
.A2(n_1285),
.B(n_1287),
.Y(n_11456)
);

OAI21xp5_ASAP7_75t_L g11457 ( 
.A1(n_11273),
.A2(n_10918),
.B(n_10600),
.Y(n_11457)
);

AO31x2_ASAP7_75t_L g11458 ( 
.A1(n_11092),
.A2(n_1290),
.A3(n_1287),
.B(n_1289),
.Y(n_11458)
);

NAND2xp5_ASAP7_75t_L g11459 ( 
.A(n_11103),
.B(n_1289),
.Y(n_11459)
);

AOI21xp5_ASAP7_75t_L g11460 ( 
.A1(n_10638),
.A2(n_1290),
.B(n_1291),
.Y(n_11460)
);

BUFx6f_ASAP7_75t_L g11461 ( 
.A(n_10629),
.Y(n_11461)
);

INVx2_ASAP7_75t_L g11462 ( 
.A(n_10779),
.Y(n_11462)
);

OR2x2_ASAP7_75t_L g11463 ( 
.A(n_10746),
.B(n_1291),
.Y(n_11463)
);

INVx4_ASAP7_75t_L g11464 ( 
.A(n_10610),
.Y(n_11464)
);

INVx5_ASAP7_75t_L g11465 ( 
.A(n_11263),
.Y(n_11465)
);

BUFx12f_ASAP7_75t_L g11466 ( 
.A(n_11248),
.Y(n_11466)
);

OAI21x1_ASAP7_75t_L g11467 ( 
.A1(n_10803),
.A2(n_1292),
.B(n_1293),
.Y(n_11467)
);

AO31x2_ASAP7_75t_L g11468 ( 
.A1(n_11062),
.A2(n_1294),
.A3(n_1292),
.B(n_1293),
.Y(n_11468)
);

OA21x2_ASAP7_75t_L g11469 ( 
.A1(n_11013),
.A2(n_1294),
.B(n_1295),
.Y(n_11469)
);

NAND2xp5_ASAP7_75t_L g11470 ( 
.A(n_10649),
.B(n_10655),
.Y(n_11470)
);

OAI21x1_ASAP7_75t_L g11471 ( 
.A1(n_11050),
.A2(n_1295),
.B(n_1296),
.Y(n_11471)
);

OAI21x1_ASAP7_75t_L g11472 ( 
.A1(n_11093),
.A2(n_1296),
.B(n_1297),
.Y(n_11472)
);

OAI21x1_ASAP7_75t_L g11473 ( 
.A1(n_10744),
.A2(n_11028),
.B(n_10605),
.Y(n_11473)
);

AOI21xp5_ASAP7_75t_L g11474 ( 
.A1(n_10884),
.A2(n_1297),
.B(n_1298),
.Y(n_11474)
);

NAND2xp5_ASAP7_75t_SL g11475 ( 
.A(n_11080),
.B(n_1298),
.Y(n_11475)
);

NAND2x1_ASAP7_75t_L g11476 ( 
.A(n_10573),
.B(n_1300),
.Y(n_11476)
);

NAND2xp5_ASAP7_75t_L g11477 ( 
.A(n_10687),
.B(n_1300),
.Y(n_11477)
);

NAND2xp5_ASAP7_75t_L g11478 ( 
.A(n_10726),
.B(n_10859),
.Y(n_11478)
);

INVx1_ASAP7_75t_L g11479 ( 
.A(n_11265),
.Y(n_11479)
);

INVx2_ASAP7_75t_L g11480 ( 
.A(n_11288),
.Y(n_11480)
);

INVx5_ASAP7_75t_L g11481 ( 
.A(n_10601),
.Y(n_11481)
);

AO21x1_ASAP7_75t_L g11482 ( 
.A1(n_11011),
.A2(n_1301),
.B(n_1302),
.Y(n_11482)
);

INVx1_ASAP7_75t_L g11483 ( 
.A(n_10571),
.Y(n_11483)
);

OAI21x1_ASAP7_75t_L g11484 ( 
.A1(n_10594),
.A2(n_1301),
.B(n_1303),
.Y(n_11484)
);

AND2x2_ASAP7_75t_L g11485 ( 
.A(n_10835),
.B(n_1304),
.Y(n_11485)
);

AO31x2_ASAP7_75t_L g11486 ( 
.A1(n_10815),
.A2(n_1306),
.A3(n_1304),
.B(n_1305),
.Y(n_11486)
);

AO21x2_ASAP7_75t_L g11487 ( 
.A1(n_10614),
.A2(n_1305),
.B(n_1307),
.Y(n_11487)
);

OAI21x1_ASAP7_75t_L g11488 ( 
.A1(n_10607),
.A2(n_1308),
.B(n_1309),
.Y(n_11488)
);

AOI21xp5_ASAP7_75t_L g11489 ( 
.A1(n_10597),
.A2(n_1308),
.B(n_1309),
.Y(n_11489)
);

NOR2xp33_ASAP7_75t_L g11490 ( 
.A(n_10721),
.B(n_1310),
.Y(n_11490)
);

A2O1A1Ixp33_ASAP7_75t_L g11491 ( 
.A1(n_11213),
.A2(n_1312),
.B(n_1310),
.C(n_1311),
.Y(n_11491)
);

NOR2xp67_ASAP7_75t_L g11492 ( 
.A(n_10787),
.B(n_1312),
.Y(n_11492)
);

NOR2xp67_ASAP7_75t_L g11493 ( 
.A(n_11080),
.B(n_1313),
.Y(n_11493)
);

AND2x2_ASAP7_75t_L g11494 ( 
.A(n_10840),
.B(n_1313),
.Y(n_11494)
);

INVx3_ASAP7_75t_L g11495 ( 
.A(n_10603),
.Y(n_11495)
);

CKINVDCx8_ASAP7_75t_R g11496 ( 
.A(n_10620),
.Y(n_11496)
);

INVx3_ASAP7_75t_L g11497 ( 
.A(n_10609),
.Y(n_11497)
);

BUFx2_ASAP7_75t_L g11498 ( 
.A(n_10618),
.Y(n_11498)
);

BUFx3_ASAP7_75t_L g11499 ( 
.A(n_10630),
.Y(n_11499)
);

AOI21xp5_ASAP7_75t_L g11500 ( 
.A1(n_10983),
.A2(n_1315),
.B(n_1316),
.Y(n_11500)
);

OAI21x1_ASAP7_75t_L g11501 ( 
.A1(n_10621),
.A2(n_1315),
.B(n_1316),
.Y(n_11501)
);

A2O1A1Ixp33_ASAP7_75t_L g11502 ( 
.A1(n_11109),
.A2(n_1319),
.B(n_1317),
.C(n_1318),
.Y(n_11502)
);

NOR2x1_ASAP7_75t_L g11503 ( 
.A(n_11002),
.B(n_1317),
.Y(n_11503)
);

OAI21x1_ASAP7_75t_L g11504 ( 
.A1(n_10668),
.A2(n_1319),
.B(n_1320),
.Y(n_11504)
);

AOI21xp5_ASAP7_75t_L g11505 ( 
.A1(n_11235),
.A2(n_1320),
.B(n_1321),
.Y(n_11505)
);

O2A1O1Ixp5_ASAP7_75t_SL g11506 ( 
.A1(n_10919),
.A2(n_1323),
.B(n_1321),
.C(n_1322),
.Y(n_11506)
);

AO31x2_ASAP7_75t_L g11507 ( 
.A1(n_10854),
.A2(n_1325),
.A3(n_1322),
.B(n_1324),
.Y(n_11507)
);

INVx3_ASAP7_75t_L g11508 ( 
.A(n_10851),
.Y(n_11508)
);

NAND2xp5_ASAP7_75t_L g11509 ( 
.A(n_11140),
.B(n_1324),
.Y(n_11509)
);

NOR2xp67_ASAP7_75t_L g11510 ( 
.A(n_10810),
.B(n_10843),
.Y(n_11510)
);

AOI21xp5_ASAP7_75t_L g11511 ( 
.A1(n_10646),
.A2(n_1325),
.B(n_1326),
.Y(n_11511)
);

AOI21x1_ASAP7_75t_L g11512 ( 
.A1(n_10624),
.A2(n_1326),
.B(n_1327),
.Y(n_11512)
);

OAI21x1_ASAP7_75t_SL g11513 ( 
.A1(n_10747),
.A2(n_1327),
.B(n_1328),
.Y(n_11513)
);

OAI21x1_ASAP7_75t_L g11514 ( 
.A1(n_10674),
.A2(n_1329),
.B(n_1330),
.Y(n_11514)
);

AOI21xp5_ASAP7_75t_L g11515 ( 
.A1(n_10648),
.A2(n_1329),
.B(n_1330),
.Y(n_11515)
);

NAND2xp5_ASAP7_75t_L g11516 ( 
.A(n_11144),
.B(n_1331),
.Y(n_11516)
);

NOR2xp33_ASAP7_75t_R g11517 ( 
.A(n_11279),
.B(n_1331),
.Y(n_11517)
);

OR2x2_ASAP7_75t_L g11518 ( 
.A(n_10581),
.B(n_1332),
.Y(n_11518)
);

CKINVDCx20_ASAP7_75t_R g11519 ( 
.A(n_10667),
.Y(n_11519)
);

OAI21x1_ASAP7_75t_L g11520 ( 
.A1(n_10683),
.A2(n_1332),
.B(n_1333),
.Y(n_11520)
);

AOI21xp5_ASAP7_75t_L g11521 ( 
.A1(n_11182),
.A2(n_1334),
.B(n_1335),
.Y(n_11521)
);

NAND2xp5_ASAP7_75t_SL g11522 ( 
.A(n_11078),
.B(n_1334),
.Y(n_11522)
);

AND2x4_ASAP7_75t_L g11523 ( 
.A(n_10745),
.B(n_1335),
.Y(n_11523)
);

OAI21x1_ASAP7_75t_L g11524 ( 
.A1(n_10697),
.A2(n_10716),
.B(n_10715),
.Y(n_11524)
);

OAI22xp5_ASAP7_75t_L g11525 ( 
.A1(n_11160),
.A2(n_1339),
.B1(n_1336),
.B2(n_1337),
.Y(n_11525)
);

NAND2xp5_ASAP7_75t_L g11526 ( 
.A(n_11145),
.B(n_1336),
.Y(n_11526)
);

OAI21x1_ASAP7_75t_L g11527 ( 
.A1(n_10728),
.A2(n_1339),
.B(n_1340),
.Y(n_11527)
);

CKINVDCx6p67_ASAP7_75t_R g11528 ( 
.A(n_10693),
.Y(n_11528)
);

AOI31xp67_ASAP7_75t_L g11529 ( 
.A1(n_11006),
.A2(n_1342),
.A3(n_1340),
.B(n_1341),
.Y(n_11529)
);

OAI21x1_ASAP7_75t_L g11530 ( 
.A1(n_10732),
.A2(n_1342),
.B(n_1343),
.Y(n_11530)
);

OAI21x1_ASAP7_75t_L g11531 ( 
.A1(n_10738),
.A2(n_1343),
.B(n_1344),
.Y(n_11531)
);

NAND2xp5_ASAP7_75t_SL g11532 ( 
.A(n_11078),
.B(n_1344),
.Y(n_11532)
);

AO31x2_ASAP7_75t_L g11533 ( 
.A1(n_10635),
.A2(n_1347),
.A3(n_1345),
.B(n_1346),
.Y(n_11533)
);

AND2x4_ASAP7_75t_L g11534 ( 
.A(n_10651),
.B(n_1345),
.Y(n_11534)
);

OAI21xp5_ASAP7_75t_L g11535 ( 
.A1(n_10795),
.A2(n_1346),
.B(n_1347),
.Y(n_11535)
);

AO31x2_ASAP7_75t_L g11536 ( 
.A1(n_10636),
.A2(n_1350),
.A3(n_1348),
.B(n_1349),
.Y(n_11536)
);

OAI21x1_ASAP7_75t_L g11537 ( 
.A1(n_10758),
.A2(n_1348),
.B(n_1349),
.Y(n_11537)
);

OAI21x1_ASAP7_75t_L g11538 ( 
.A1(n_11016),
.A2(n_1350),
.B(n_1351),
.Y(n_11538)
);

OAI21x1_ASAP7_75t_SL g11539 ( 
.A1(n_10634),
.A2(n_1351),
.B(n_1352),
.Y(n_11539)
);

NAND2xp5_ASAP7_75t_L g11540 ( 
.A(n_11042),
.B(n_1353),
.Y(n_11540)
);

NAND2xp5_ASAP7_75t_L g11541 ( 
.A(n_11124),
.B(n_1353),
.Y(n_11541)
);

AND2x2_ASAP7_75t_L g11542 ( 
.A(n_10963),
.B(n_1354),
.Y(n_11542)
);

AOI21xp5_ASAP7_75t_L g11543 ( 
.A1(n_10767),
.A2(n_1354),
.B(n_1355),
.Y(n_11543)
);

CKINVDCx5p33_ASAP7_75t_R g11544 ( 
.A(n_10725),
.Y(n_11544)
);

AOI21xp5_ASAP7_75t_SL g11545 ( 
.A1(n_10982),
.A2(n_1355),
.B(n_1356),
.Y(n_11545)
);

NOR2xp33_ASAP7_75t_L g11546 ( 
.A(n_10900),
.B(n_1356),
.Y(n_11546)
);

OAI21x1_ASAP7_75t_L g11547 ( 
.A1(n_10763),
.A2(n_1357),
.B(n_1358),
.Y(n_11547)
);

AOI21xp5_ASAP7_75t_L g11548 ( 
.A1(n_10802),
.A2(n_1357),
.B(n_1358),
.Y(n_11548)
);

AO31x2_ASAP7_75t_L g11549 ( 
.A1(n_10642),
.A2(n_1362),
.A3(n_1359),
.B(n_1360),
.Y(n_11549)
);

AOI211x1_ASAP7_75t_L g11550 ( 
.A1(n_10711),
.A2(n_1364),
.B(n_1360),
.C(n_1363),
.Y(n_11550)
);

OR2x2_ASAP7_75t_L g11551 ( 
.A(n_11254),
.B(n_1363),
.Y(n_11551)
);

OAI22xp5_ASAP7_75t_L g11552 ( 
.A1(n_10987),
.A2(n_1367),
.B1(n_1365),
.B2(n_1366),
.Y(n_11552)
);

NAND2xp5_ASAP7_75t_L g11553 ( 
.A(n_11130),
.B(n_1365),
.Y(n_11553)
);

OAI21x1_ASAP7_75t_L g11554 ( 
.A1(n_10764),
.A2(n_1366),
.B(n_1367),
.Y(n_11554)
);

AND2x2_ASAP7_75t_SL g11555 ( 
.A(n_10805),
.B(n_1368),
.Y(n_11555)
);

OAI21x1_ASAP7_75t_L g11556 ( 
.A1(n_10772),
.A2(n_10789),
.B(n_10786),
.Y(n_11556)
);

INVx5_ASAP7_75t_L g11557 ( 
.A(n_10601),
.Y(n_11557)
);

INVx1_ASAP7_75t_L g11558 ( 
.A(n_10821),
.Y(n_11558)
);

OAI21x1_ASAP7_75t_L g11559 ( 
.A1(n_10796),
.A2(n_1368),
.B(n_1369),
.Y(n_11559)
);

NAND2x1p5_ASAP7_75t_L g11560 ( 
.A(n_10709),
.B(n_1371),
.Y(n_11560)
);

OAI21x1_ASAP7_75t_L g11561 ( 
.A1(n_10811),
.A2(n_1371),
.B(n_1372),
.Y(n_11561)
);

INVx2_ASAP7_75t_L g11562 ( 
.A(n_10800),
.Y(n_11562)
);

AOI21x1_ASAP7_75t_L g11563 ( 
.A1(n_10944),
.A2(n_1373),
.B(n_1374),
.Y(n_11563)
);

AOI21xp5_ASAP7_75t_L g11564 ( 
.A1(n_10823),
.A2(n_10836),
.B(n_10825),
.Y(n_11564)
);

NAND2xp5_ASAP7_75t_L g11565 ( 
.A(n_11134),
.B(n_11141),
.Y(n_11565)
);

AO31x2_ASAP7_75t_L g11566 ( 
.A1(n_10565),
.A2(n_10580),
.A3(n_11242),
.B(n_11238),
.Y(n_11566)
);

INVx3_ASAP7_75t_SL g11567 ( 
.A(n_10616),
.Y(n_11567)
);

AND2x2_ASAP7_75t_L g11568 ( 
.A(n_10941),
.B(n_1373),
.Y(n_11568)
);

AOI21xp5_ASAP7_75t_L g11569 ( 
.A1(n_10873),
.A2(n_1374),
.B(n_1376),
.Y(n_11569)
);

NAND2xp5_ASAP7_75t_L g11570 ( 
.A(n_11139),
.B(n_10997),
.Y(n_11570)
);

BUFx3_ASAP7_75t_L g11571 ( 
.A(n_10792),
.Y(n_11571)
);

OAI21xp5_ASAP7_75t_L g11572 ( 
.A1(n_10995),
.A2(n_1376),
.B(n_1377),
.Y(n_11572)
);

OAI21xp5_ASAP7_75t_L g11573 ( 
.A1(n_10741),
.A2(n_1377),
.B(n_1378),
.Y(n_11573)
);

NAND2xp5_ASAP7_75t_SL g11574 ( 
.A(n_11094),
.B(n_1378),
.Y(n_11574)
);

NAND2xp5_ASAP7_75t_L g11575 ( 
.A(n_11081),
.B(n_1379),
.Y(n_11575)
);

AOI21xp5_ASAP7_75t_L g11576 ( 
.A1(n_10584),
.A2(n_10808),
.B(n_10718),
.Y(n_11576)
);

NAND2xp5_ASAP7_75t_L g11577 ( 
.A(n_10788),
.B(n_1380),
.Y(n_11577)
);

OAI21xp33_ASAP7_75t_L g11578 ( 
.A1(n_10640),
.A2(n_1380),
.B(n_1381),
.Y(n_11578)
);

OAI22xp5_ASAP7_75t_L g11579 ( 
.A1(n_10807),
.A2(n_1383),
.B1(n_1381),
.B2(n_1382),
.Y(n_11579)
);

NAND2xp33_ASAP7_75t_SL g11580 ( 
.A(n_10613),
.B(n_1383),
.Y(n_11580)
);

NAND2xp5_ASAP7_75t_L g11581 ( 
.A(n_10617),
.B(n_1384),
.Y(n_11581)
);

AND2x2_ASAP7_75t_L g11582 ( 
.A(n_10572),
.B(n_1384),
.Y(n_11582)
);

OAI21x1_ASAP7_75t_L g11583 ( 
.A1(n_10814),
.A2(n_1385),
.B(n_1386),
.Y(n_11583)
);

INVx1_ASAP7_75t_L g11584 ( 
.A(n_10850),
.Y(n_11584)
);

AND2x4_ASAP7_75t_L g11585 ( 
.A(n_10704),
.B(n_1385),
.Y(n_11585)
);

AOI21xp5_ASAP7_75t_SL g11586 ( 
.A1(n_11051),
.A2(n_1386),
.B(n_1387),
.Y(n_11586)
);

NAND2xp5_ASAP7_75t_L g11587 ( 
.A(n_11090),
.B(n_1387),
.Y(n_11587)
);

INVx2_ASAP7_75t_L g11588 ( 
.A(n_10801),
.Y(n_11588)
);

OAI21xp5_ASAP7_75t_L g11589 ( 
.A1(n_10653),
.A2(n_1388),
.B(n_1389),
.Y(n_11589)
);

OA21x2_ASAP7_75t_L g11590 ( 
.A1(n_10622),
.A2(n_1388),
.B(n_1389),
.Y(n_11590)
);

AOI21xp5_ASAP7_75t_L g11591 ( 
.A1(n_10623),
.A2(n_1390),
.B(n_1392),
.Y(n_11591)
);

AO31x2_ASAP7_75t_L g11592 ( 
.A1(n_11257),
.A2(n_1393),
.A3(n_1390),
.B(n_1392),
.Y(n_11592)
);

OA22x2_ASAP7_75t_L g11593 ( 
.A1(n_10599),
.A2(n_1395),
.B1(n_1393),
.B2(n_1394),
.Y(n_11593)
);

AOI22xp5_ASAP7_75t_L g11594 ( 
.A1(n_11151),
.A2(n_1396),
.B1(n_1394),
.B2(n_1395),
.Y(n_11594)
);

AOI211x1_ASAP7_75t_L g11595 ( 
.A1(n_11261),
.A2(n_11172),
.B(n_10985),
.C(n_11275),
.Y(n_11595)
);

NAND2xp5_ASAP7_75t_L g11596 ( 
.A(n_10736),
.B(n_1396),
.Y(n_11596)
);

NAND2xp5_ASAP7_75t_L g11597 ( 
.A(n_10650),
.B(n_1397),
.Y(n_11597)
);

OAI21x1_ASAP7_75t_L g11598 ( 
.A1(n_10816),
.A2(n_1397),
.B(n_1398),
.Y(n_11598)
);

AND2x2_ASAP7_75t_L g11599 ( 
.A(n_11250),
.B(n_1398),
.Y(n_11599)
);

AOI21xp5_ASAP7_75t_L g11600 ( 
.A1(n_10872),
.A2(n_1399),
.B(n_1400),
.Y(n_11600)
);

OAI22xp5_ASAP7_75t_L g11601 ( 
.A1(n_11059),
.A2(n_1401),
.B1(n_1399),
.B2(n_1400),
.Y(n_11601)
);

NAND2x1p5_ASAP7_75t_L g11602 ( 
.A(n_10693),
.B(n_1402),
.Y(n_11602)
);

AOI21xp5_ASAP7_75t_L g11603 ( 
.A1(n_11262),
.A2(n_1402),
.B(n_1403),
.Y(n_11603)
);

INVx1_ASAP7_75t_L g11604 ( 
.A(n_10857),
.Y(n_11604)
);

A2O1A1Ixp33_ASAP7_75t_L g11605 ( 
.A1(n_11211),
.A2(n_1406),
.B(n_1404),
.C(n_1405),
.Y(n_11605)
);

NAND2xp5_ASAP7_75t_L g11606 ( 
.A(n_10650),
.B(n_1405),
.Y(n_11606)
);

OAI21x1_ASAP7_75t_L g11607 ( 
.A1(n_10820),
.A2(n_10829),
.B(n_10826),
.Y(n_11607)
);

AOI21x1_ASAP7_75t_L g11608 ( 
.A1(n_10661),
.A2(n_1407),
.B(n_1408),
.Y(n_11608)
);

NAND2xp5_ASAP7_75t_SL g11609 ( 
.A(n_11094),
.B(n_1407),
.Y(n_11609)
);

AO31x2_ASAP7_75t_L g11610 ( 
.A1(n_11085),
.A2(n_11009),
.A3(n_10576),
.B(n_10864),
.Y(n_11610)
);

AND2x2_ASAP7_75t_L g11611 ( 
.A(n_10901),
.B(n_1408),
.Y(n_11611)
);

AO21x2_ASAP7_75t_L g11612 ( 
.A1(n_10971),
.A2(n_1409),
.B(n_1410),
.Y(n_11612)
);

AOI21xp5_ASAP7_75t_L g11613 ( 
.A1(n_11277),
.A2(n_1409),
.B(n_1410),
.Y(n_11613)
);

NAND3xp33_ASAP7_75t_SL g11614 ( 
.A(n_10662),
.B(n_1411),
.C(n_1412),
.Y(n_11614)
);

NAND2xp5_ASAP7_75t_L g11615 ( 
.A(n_10650),
.B(n_1411),
.Y(n_11615)
);

AO31x2_ASAP7_75t_L g11616 ( 
.A1(n_10861),
.A2(n_1414),
.A3(n_1412),
.B(n_1413),
.Y(n_11616)
);

OAI21xp5_ASAP7_75t_L g11617 ( 
.A1(n_11271),
.A2(n_11053),
.B(n_11043),
.Y(n_11617)
);

NAND2xp5_ASAP7_75t_L g11618 ( 
.A(n_11102),
.B(n_1413),
.Y(n_11618)
);

OAI22xp5_ASAP7_75t_L g11619 ( 
.A1(n_11084),
.A2(n_1416),
.B1(n_1414),
.B2(n_1415),
.Y(n_11619)
);

INVx2_ASAP7_75t_L g11620 ( 
.A(n_10887),
.Y(n_11620)
);

NAND2xp5_ASAP7_75t_L g11621 ( 
.A(n_11102),
.B(n_1415),
.Y(n_11621)
);

NOR2xp33_ASAP7_75t_L g11622 ( 
.A(n_10574),
.B(n_1416),
.Y(n_11622)
);

AOI21xp5_ASAP7_75t_L g11623 ( 
.A1(n_10619),
.A2(n_1417),
.B(n_1418),
.Y(n_11623)
);

AOI21xp5_ASAP7_75t_L g11624 ( 
.A1(n_10639),
.A2(n_1418),
.B(n_1419),
.Y(n_11624)
);

NAND2xp5_ASAP7_75t_L g11625 ( 
.A(n_10906),
.B(n_1419),
.Y(n_11625)
);

NAND3xp33_ASAP7_75t_SL g11626 ( 
.A(n_10753),
.B(n_10959),
.C(n_10951),
.Y(n_11626)
);

NAND2xp5_ASAP7_75t_SL g11627 ( 
.A(n_11104),
.B(n_1420),
.Y(n_11627)
);

BUFx6f_ASAP7_75t_L g11628 ( 
.A(n_10629),
.Y(n_11628)
);

OAI21x1_ASAP7_75t_L g11629 ( 
.A1(n_10837),
.A2(n_1421),
.B(n_1422),
.Y(n_11629)
);

OAI22x1_ASAP7_75t_L g11630 ( 
.A1(n_11033),
.A2(n_1423),
.B1(n_1421),
.B2(n_1422),
.Y(n_11630)
);

OAI21xp5_ASAP7_75t_SL g11631 ( 
.A1(n_10895),
.A2(n_1424),
.B(n_1425),
.Y(n_11631)
);

INVx1_ASAP7_75t_L g11632 ( 
.A(n_10883),
.Y(n_11632)
);

NAND2xp5_ASAP7_75t_L g11633 ( 
.A(n_10637),
.B(n_1425),
.Y(n_11633)
);

A2O1A1Ixp33_ASAP7_75t_L g11634 ( 
.A1(n_10712),
.A2(n_11116),
.B(n_10734),
.C(n_10626),
.Y(n_11634)
);

OAI21xp5_ASAP7_75t_L g11635 ( 
.A1(n_10606),
.A2(n_1426),
.B(n_1427),
.Y(n_11635)
);

NAND2xp5_ASAP7_75t_L g11636 ( 
.A(n_10833),
.B(n_1426),
.Y(n_11636)
);

AOI221xp5_ASAP7_75t_L g11637 ( 
.A1(n_10675),
.A2(n_11087),
.B1(n_11024),
.B2(n_10888),
.C(n_10680),
.Y(n_11637)
);

AOI21xp5_ASAP7_75t_L g11638 ( 
.A1(n_10932),
.A2(n_1428),
.B(n_1429),
.Y(n_11638)
);

NAND3xp33_ASAP7_75t_L g11639 ( 
.A(n_11225),
.B(n_1428),
.C(n_1429),
.Y(n_11639)
);

INVx1_ASAP7_75t_L g11640 ( 
.A(n_10889),
.Y(n_11640)
);

AOI21xp5_ASAP7_75t_L g11641 ( 
.A1(n_10946),
.A2(n_1430),
.B(n_1431),
.Y(n_11641)
);

INVx1_ASAP7_75t_L g11642 ( 
.A(n_10908),
.Y(n_11642)
);

AO21x2_ASAP7_75t_L g11643 ( 
.A1(n_11029),
.A2(n_1430),
.B(n_1431),
.Y(n_11643)
);

AOI21xp5_ASAP7_75t_L g11644 ( 
.A1(n_11012),
.A2(n_1432),
.B(n_1433),
.Y(n_11644)
);

AND2x2_ASAP7_75t_L g11645 ( 
.A(n_10591),
.B(n_1432),
.Y(n_11645)
);

OAI21x1_ASAP7_75t_L g11646 ( 
.A1(n_10838),
.A2(n_1433),
.B(n_1434),
.Y(n_11646)
);

INVx3_ASAP7_75t_L g11647 ( 
.A(n_10845),
.Y(n_11647)
);

AND2x2_ASAP7_75t_L g11648 ( 
.A(n_11138),
.B(n_1435),
.Y(n_11648)
);

OAI21x1_ASAP7_75t_L g11649 ( 
.A1(n_10842),
.A2(n_1436),
.B(n_1437),
.Y(n_11649)
);

INVx1_ASAP7_75t_L g11650 ( 
.A(n_10916),
.Y(n_11650)
);

AOI21xp5_ASAP7_75t_L g11651 ( 
.A1(n_10891),
.A2(n_1436),
.B(n_1437),
.Y(n_11651)
);

BUFx10_ASAP7_75t_L g11652 ( 
.A(n_10699),
.Y(n_11652)
);

NAND2xp5_ASAP7_75t_L g11653 ( 
.A(n_11165),
.B(n_1438),
.Y(n_11653)
);

INVx1_ASAP7_75t_L g11654 ( 
.A(n_10927),
.Y(n_11654)
);

NAND2xp5_ASAP7_75t_L g11655 ( 
.A(n_10830),
.B(n_1438),
.Y(n_11655)
);

OAI21x1_ASAP7_75t_L g11656 ( 
.A1(n_10866),
.A2(n_1439),
.B(n_1440),
.Y(n_11656)
);

OAI21x1_ASAP7_75t_L g11657 ( 
.A1(n_10870),
.A2(n_1439),
.B(n_1440),
.Y(n_11657)
);

NAND3xp33_ASAP7_75t_SL g11658 ( 
.A(n_10899),
.B(n_1441),
.C(n_1442),
.Y(n_11658)
);

OAI21x1_ASAP7_75t_L g11659 ( 
.A1(n_10871),
.A2(n_1441),
.B(n_1442),
.Y(n_11659)
);

AOI21xp5_ASAP7_75t_L g11660 ( 
.A1(n_10898),
.A2(n_1443),
.B(n_1444),
.Y(n_11660)
);

BUFx2_ASAP7_75t_L g11661 ( 
.A(n_10660),
.Y(n_11661)
);

INVx3_ASAP7_75t_L g11662 ( 
.A(n_10845),
.Y(n_11662)
);

BUFx4f_ASAP7_75t_L g11663 ( 
.A(n_10671),
.Y(n_11663)
);

OAI22xp5_ASAP7_75t_L g11664 ( 
.A1(n_10790),
.A2(n_1445),
.B1(n_1443),
.B2(n_1444),
.Y(n_11664)
);

AOI21x1_ASAP7_75t_L g11665 ( 
.A1(n_10834),
.A2(n_1445),
.B(n_1446),
.Y(n_11665)
);

HB1xp67_ASAP7_75t_L g11666 ( 
.A(n_11086),
.Y(n_11666)
);

OAI21x1_ASAP7_75t_L g11667 ( 
.A1(n_10881),
.A2(n_1446),
.B(n_1447),
.Y(n_11667)
);

INVx1_ASAP7_75t_L g11668 ( 
.A(n_10928),
.Y(n_11668)
);

AOI21xp5_ASAP7_75t_L g11669 ( 
.A1(n_10910),
.A2(n_1447),
.B(n_1448),
.Y(n_11669)
);

OAI22xp5_ASAP7_75t_L g11670 ( 
.A1(n_10706),
.A2(n_1450),
.B1(n_1448),
.B2(n_1449),
.Y(n_11670)
);

NAND2xp5_ASAP7_75t_L g11671 ( 
.A(n_10765),
.B(n_1449),
.Y(n_11671)
);

OAI21x1_ASAP7_75t_L g11672 ( 
.A1(n_10894),
.A2(n_1450),
.B(n_1451),
.Y(n_11672)
);

AND2x2_ASAP7_75t_L g11673 ( 
.A(n_10589),
.B(n_1451),
.Y(n_11673)
);

OAI22xp5_ASAP7_75t_L g11674 ( 
.A1(n_10998),
.A2(n_1454),
.B1(n_1452),
.B2(n_1453),
.Y(n_11674)
);

NOR2xp33_ASAP7_75t_L g11675 ( 
.A(n_10574),
.B(n_1453),
.Y(n_11675)
);

AO31x2_ASAP7_75t_L g11676 ( 
.A1(n_10911),
.A2(n_1456),
.A3(n_1454),
.B(n_1455),
.Y(n_11676)
);

OAI21xp33_ASAP7_75t_L g11677 ( 
.A1(n_10848),
.A2(n_1455),
.B(n_1456),
.Y(n_11677)
);

NAND2x1p5_ASAP7_75t_L g11678 ( 
.A(n_11239),
.B(n_1457),
.Y(n_11678)
);

AO31x2_ASAP7_75t_L g11679 ( 
.A1(n_10931),
.A2(n_1460),
.A3(n_1458),
.B(n_1459),
.Y(n_11679)
);

OA22x2_ASAP7_75t_L g11680 ( 
.A1(n_11064),
.A2(n_1460),
.B1(n_1458),
.B2(n_1459),
.Y(n_11680)
);

OAI22xp5_ASAP7_75t_L g11681 ( 
.A1(n_10998),
.A2(n_1463),
.B1(n_1461),
.B2(n_1462),
.Y(n_11681)
);

AOI21xp5_ASAP7_75t_L g11682 ( 
.A1(n_11034),
.A2(n_1462),
.B(n_1463),
.Y(n_11682)
);

NAND2xp5_ASAP7_75t_L g11683 ( 
.A(n_10770),
.B(n_1464),
.Y(n_11683)
);

NAND2xp5_ASAP7_75t_L g11684 ( 
.A(n_10739),
.B(n_1465),
.Y(n_11684)
);

OAI21x1_ASAP7_75t_L g11685 ( 
.A1(n_10902),
.A2(n_1465),
.B(n_1466),
.Y(n_11685)
);

NAND2xp5_ASAP7_75t_SL g11686 ( 
.A(n_11104),
.B(n_1466),
.Y(n_11686)
);

AOI21x1_ASAP7_75t_SL g11687 ( 
.A1(n_10948),
.A2(n_1467),
.B(n_1468),
.Y(n_11687)
);

BUFx6f_ASAP7_75t_SL g11688 ( 
.A(n_10689),
.Y(n_11688)
);

INVx1_ASAP7_75t_L g11689 ( 
.A(n_10937),
.Y(n_11689)
);

OAI21x1_ASAP7_75t_L g11690 ( 
.A1(n_10926),
.A2(n_1468),
.B(n_1469),
.Y(n_11690)
);

OAI21x1_ASAP7_75t_L g11691 ( 
.A1(n_10939),
.A2(n_1469),
.B(n_1470),
.Y(n_11691)
);

CKINVDCx8_ASAP7_75t_R g11692 ( 
.A(n_10595),
.Y(n_11692)
);

AO32x2_ASAP7_75t_L g11693 ( 
.A1(n_10592),
.A2(n_11071),
.A3(n_10665),
.B1(n_10659),
.B2(n_10991),
.Y(n_11693)
);

NAND2xp5_ASAP7_75t_SL g11694 ( 
.A(n_11112),
.B(n_1470),
.Y(n_11694)
);

INVx1_ASAP7_75t_L g11695 ( 
.A(n_10938),
.Y(n_11695)
);

NAND2xp5_ASAP7_75t_L g11696 ( 
.A(n_10791),
.B(n_1471),
.Y(n_11696)
);

INVx1_ASAP7_75t_L g11697 ( 
.A(n_10964),
.Y(n_11697)
);

AOI22xp5_ASAP7_75t_L g11698 ( 
.A1(n_11082),
.A2(n_1473),
.B1(n_1471),
.B2(n_1472),
.Y(n_11698)
);

AND2x4_ASAP7_75t_L g11699 ( 
.A(n_10700),
.B(n_1472),
.Y(n_11699)
);

AO22x2_ASAP7_75t_L g11700 ( 
.A1(n_10990),
.A2(n_1475),
.B1(n_1473),
.B2(n_1474),
.Y(n_11700)
);

BUFx6f_ASAP7_75t_L g11701 ( 
.A(n_10724),
.Y(n_11701)
);

AOI21xp5_ASAP7_75t_L g11702 ( 
.A1(n_11041),
.A2(n_1475),
.B(n_1476),
.Y(n_11702)
);

OAI21x1_ASAP7_75t_L g11703 ( 
.A1(n_10942),
.A2(n_1476),
.B(n_1477),
.Y(n_11703)
);

INVx1_ASAP7_75t_L g11704 ( 
.A(n_10996),
.Y(n_11704)
);

OAI21x1_ASAP7_75t_L g11705 ( 
.A1(n_11038),
.A2(n_1477),
.B(n_1478),
.Y(n_11705)
);

NOR2xp33_ASAP7_75t_L g11706 ( 
.A(n_10595),
.B(n_11264),
.Y(n_11706)
);

NAND2xp5_ASAP7_75t_SL g11707 ( 
.A(n_11112),
.B(n_1478),
.Y(n_11707)
);

NAND2xp5_ASAP7_75t_SL g11708 ( 
.A(n_11174),
.B(n_11208),
.Y(n_11708)
);

NAND2xp5_ASAP7_75t_L g11709 ( 
.A(n_10841),
.B(n_1479),
.Y(n_11709)
);

AOI21xp5_ASAP7_75t_L g11710 ( 
.A1(n_10949),
.A2(n_1479),
.B(n_1480),
.Y(n_11710)
);

NOR2xp67_ASAP7_75t_SL g11711 ( 
.A(n_11208),
.B(n_1480),
.Y(n_11711)
);

NAND2xp5_ASAP7_75t_L g11712 ( 
.A(n_10567),
.B(n_11283),
.Y(n_11712)
);

OAI21x1_ASAP7_75t_L g11713 ( 
.A1(n_10604),
.A2(n_1481),
.B(n_1482),
.Y(n_11713)
);

INVx2_ASAP7_75t_SL g11714 ( 
.A(n_11286),
.Y(n_11714)
);

AOI21xp5_ASAP7_75t_L g11715 ( 
.A1(n_10993),
.A2(n_1481),
.B(n_1482),
.Y(n_11715)
);

NAND2xp5_ASAP7_75t_L g11716 ( 
.A(n_10782),
.B(n_1483),
.Y(n_11716)
);

AOI21x1_ASAP7_75t_L g11717 ( 
.A1(n_10909),
.A2(n_1483),
.B(n_1484),
.Y(n_11717)
);

AO31x2_ASAP7_75t_L g11718 ( 
.A1(n_11003),
.A2(n_11035),
.A3(n_11054),
.B(n_11010),
.Y(n_11718)
);

OAI21xp5_ASAP7_75t_L g11719 ( 
.A1(n_11204),
.A2(n_1484),
.B(n_1485),
.Y(n_11719)
);

OAI21x1_ASAP7_75t_L g11720 ( 
.A1(n_10958),
.A2(n_1485),
.B(n_1486),
.Y(n_11720)
);

OAI22xp5_ASAP7_75t_L g11721 ( 
.A1(n_10694),
.A2(n_1488),
.B1(n_1486),
.B2(n_1487),
.Y(n_11721)
);

OAI21x1_ASAP7_75t_L g11722 ( 
.A1(n_11097),
.A2(n_1487),
.B(n_1489),
.Y(n_11722)
);

BUFx4_ASAP7_75t_SL g11723 ( 
.A(n_10699),
.Y(n_11723)
);

OAI21x1_ASAP7_75t_L g11724 ( 
.A1(n_10720),
.A2(n_1489),
.B(n_1491),
.Y(n_11724)
);

OAI21x1_ASAP7_75t_L g11725 ( 
.A1(n_10723),
.A2(n_1491),
.B(n_1492),
.Y(n_11725)
);

NAND2xp5_ASAP7_75t_L g11726 ( 
.A(n_10934),
.B(n_10678),
.Y(n_11726)
);

BUFx2_ASAP7_75t_L g11727 ( 
.A(n_10681),
.Y(n_11727)
);

AOI21xp5_ASAP7_75t_L g11728 ( 
.A1(n_11015),
.A2(n_1492),
.B(n_1493),
.Y(n_11728)
);

AOI21xp5_ASAP7_75t_L g11729 ( 
.A1(n_10579),
.A2(n_1493),
.B(n_1494),
.Y(n_11729)
);

HB1xp67_ASAP7_75t_L g11730 ( 
.A(n_11197),
.Y(n_11730)
);

INVx1_ASAP7_75t_L g11731 ( 
.A(n_11056),
.Y(n_11731)
);

NOR2xp33_ASAP7_75t_L g11732 ( 
.A(n_11264),
.B(n_1494),
.Y(n_11732)
);

OAI21xp5_ASAP7_75t_L g11733 ( 
.A1(n_10757),
.A2(n_1495),
.B(n_1496),
.Y(n_11733)
);

AOI21x1_ASAP7_75t_L g11734 ( 
.A1(n_10921),
.A2(n_1495),
.B(n_1496),
.Y(n_11734)
);

NAND2x1p5_ASAP7_75t_L g11735 ( 
.A(n_10794),
.B(n_1497),
.Y(n_11735)
);

AO22x2_ASAP7_75t_L g11736 ( 
.A1(n_11068),
.A2(n_1499),
.B1(n_1497),
.B2(n_1498),
.Y(n_11736)
);

AOI21xp5_ASAP7_75t_L g11737 ( 
.A1(n_10631),
.A2(n_1500),
.B(n_1501),
.Y(n_11737)
);

AOI21xp5_ASAP7_75t_L g11738 ( 
.A1(n_10645),
.A2(n_1500),
.B(n_1501),
.Y(n_11738)
);

NAND3xp33_ASAP7_75t_L g11739 ( 
.A(n_10743),
.B(n_1502),
.C(n_1503),
.Y(n_11739)
);

AND2x6_ASAP7_75t_L g11740 ( 
.A(n_10877),
.B(n_10907),
.Y(n_11740)
);

INVx1_ASAP7_75t_L g11741 ( 
.A(n_11072),
.Y(n_11741)
);

INVx2_ASAP7_75t_L g11742 ( 
.A(n_10920),
.Y(n_11742)
);

NAND2xp5_ASAP7_75t_L g11743 ( 
.A(n_10905),
.B(n_1502),
.Y(n_11743)
);

AO31x2_ASAP7_75t_L g11744 ( 
.A1(n_10950),
.A2(n_1505),
.A3(n_1503),
.B(n_1504),
.Y(n_11744)
);

AO31x2_ASAP7_75t_L g11745 ( 
.A1(n_10956),
.A2(n_1506),
.A3(n_1504),
.B(n_1505),
.Y(n_11745)
);

BUFx6f_ASAP7_75t_L g11746 ( 
.A(n_10724),
.Y(n_11746)
);

OR2x2_ASAP7_75t_L g11747 ( 
.A(n_10929),
.B(n_1507),
.Y(n_11747)
);

NAND2xp5_ASAP7_75t_L g11748 ( 
.A(n_11064),
.B(n_1508),
.Y(n_11748)
);

NOR2xp33_ASAP7_75t_L g11749 ( 
.A(n_11274),
.B(n_1508),
.Y(n_11749)
);

INVx1_ASAP7_75t_SL g11750 ( 
.A(n_11249),
.Y(n_11750)
);

OAI21x1_ASAP7_75t_L g11751 ( 
.A1(n_11231),
.A2(n_1509),
.B(n_1510),
.Y(n_11751)
);

BUFx2_ASAP7_75t_L g11752 ( 
.A(n_10762),
.Y(n_11752)
);

AOI211x1_ASAP7_75t_L g11753 ( 
.A1(n_10742),
.A2(n_1511),
.B(n_1509),
.C(n_1510),
.Y(n_11753)
);

AOI21x1_ASAP7_75t_SL g11754 ( 
.A1(n_10953),
.A2(n_1511),
.B(n_1512),
.Y(n_11754)
);

INVx1_ASAP7_75t_L g11755 ( 
.A(n_10935),
.Y(n_11755)
);

CKINVDCx8_ASAP7_75t_R g11756 ( 
.A(n_11274),
.Y(n_11756)
);

INVx1_ASAP7_75t_L g11757 ( 
.A(n_10954),
.Y(n_11757)
);

NOR2x1_ASAP7_75t_L g11758 ( 
.A(n_10831),
.B(n_1513),
.Y(n_11758)
);

AOI21xp33_ASAP7_75t_L g11759 ( 
.A1(n_11108),
.A2(n_1513),
.B(n_1514),
.Y(n_11759)
);

BUFx3_ASAP7_75t_L g11760 ( 
.A(n_11022),
.Y(n_11760)
);

NAND2xp5_ASAP7_75t_L g11761 ( 
.A(n_10690),
.B(n_1514),
.Y(n_11761)
);

NAND2xp5_ASAP7_75t_L g11762 ( 
.A(n_10696),
.B(n_1515),
.Y(n_11762)
);

A2O1A1Ixp33_ASAP7_75t_L g11763 ( 
.A1(n_11203),
.A2(n_1517),
.B(n_1515),
.C(n_1516),
.Y(n_11763)
);

OAI21xp5_ASAP7_75t_L g11764 ( 
.A1(n_10611),
.A2(n_1517),
.B(n_1518),
.Y(n_11764)
);

AOI21x1_ASAP7_75t_L g11765 ( 
.A1(n_10925),
.A2(n_1518),
.B(n_1519),
.Y(n_11765)
);

AO31x2_ASAP7_75t_L g11766 ( 
.A1(n_10733),
.A2(n_1521),
.A3(n_1519),
.B(n_1520),
.Y(n_11766)
);

NAND2xp33_ASAP7_75t_L g11767 ( 
.A(n_10684),
.B(n_1523),
.Y(n_11767)
);

AND2x2_ASAP7_75t_L g11768 ( 
.A(n_11055),
.B(n_1524),
.Y(n_11768)
);

NAND2xp5_ASAP7_75t_L g11769 ( 
.A(n_11040),
.B(n_1524),
.Y(n_11769)
);

OAI22x1_ASAP7_75t_L g11770 ( 
.A1(n_10923),
.A2(n_1527),
.B1(n_1525),
.B2(n_1526),
.Y(n_11770)
);

OAI21xp33_ASAP7_75t_SL g11771 ( 
.A1(n_10874),
.A2(n_1526),
.B(n_1528),
.Y(n_11771)
);

OAI21xp5_ASAP7_75t_L g11772 ( 
.A1(n_11168),
.A2(n_1530),
.B(n_1531),
.Y(n_11772)
);

NAND2xp5_ASAP7_75t_L g11773 ( 
.A(n_11046),
.B(n_1530),
.Y(n_11773)
);

OAI21x1_ASAP7_75t_L g11774 ( 
.A1(n_11058),
.A2(n_1532),
.B(n_1533),
.Y(n_11774)
);

OAI21x1_ASAP7_75t_L g11775 ( 
.A1(n_11048),
.A2(n_1532),
.B(n_1533),
.Y(n_11775)
);

A2O1A1Ixp33_ASAP7_75t_L g11776 ( 
.A1(n_11176),
.A2(n_1536),
.B(n_1534),
.C(n_1535),
.Y(n_11776)
);

OAI21x1_ASAP7_75t_L g11777 ( 
.A1(n_11088),
.A2(n_1534),
.B(n_1535),
.Y(n_11777)
);

OAI21x1_ASAP7_75t_L g11778 ( 
.A1(n_11166),
.A2(n_11202),
.B(n_11163),
.Y(n_11778)
);

NAND2xp5_ASAP7_75t_SL g11779 ( 
.A(n_11174),
.B(n_1536),
.Y(n_11779)
);

NAND2x1p5_ASAP7_75t_L g11780 ( 
.A(n_10705),
.B(n_1537),
.Y(n_11780)
);

OAI33xp33_ASAP7_75t_L g11781 ( 
.A1(n_10869),
.A2(n_1539),
.A3(n_1541),
.B1(n_1537),
.B2(n_1538),
.B3(n_1540),
.Y(n_11781)
);

AOI21x1_ASAP7_75t_L g11782 ( 
.A1(n_10952),
.A2(n_1538),
.B(n_1539),
.Y(n_11782)
);

OAI21xp33_ASAP7_75t_L g11783 ( 
.A1(n_10976),
.A2(n_1540),
.B(n_1541),
.Y(n_11783)
);

A2O1A1Ixp33_ASAP7_75t_L g11784 ( 
.A1(n_11045),
.A2(n_1544),
.B(n_1542),
.C(n_1543),
.Y(n_11784)
);

AOI21xp5_ASAP7_75t_L g11785 ( 
.A1(n_11173),
.A2(n_1543),
.B(n_1544),
.Y(n_11785)
);

AND2x2_ASAP7_75t_L g11786 ( 
.A(n_10798),
.B(n_1545),
.Y(n_11786)
);

NAND2xp5_ASAP7_75t_L g11787 ( 
.A(n_11065),
.B(n_1545),
.Y(n_11787)
);

OAI21xp5_ASAP7_75t_L g11788 ( 
.A1(n_11075),
.A2(n_1546),
.B(n_1547),
.Y(n_11788)
);

AND2x4_ASAP7_75t_L g11789 ( 
.A(n_10752),
.B(n_1546),
.Y(n_11789)
);

OAI22xp5_ASAP7_75t_L g11790 ( 
.A1(n_10598),
.A2(n_1549),
.B1(n_1547),
.B2(n_1548),
.Y(n_11790)
);

INVx2_ASAP7_75t_SL g11791 ( 
.A(n_10759),
.Y(n_11791)
);

OAI21x1_ASAP7_75t_L g11792 ( 
.A1(n_11077),
.A2(n_1548),
.B(n_1549),
.Y(n_11792)
);

OAI21x1_ASAP7_75t_L g11793 ( 
.A1(n_11164),
.A2(n_11171),
.B(n_11155),
.Y(n_11793)
);

AOI221xp5_ASAP7_75t_L g11794 ( 
.A1(n_11170),
.A2(n_1552),
.B1(n_1550),
.B2(n_1551),
.C(n_1553),
.Y(n_11794)
);

AOI21xp5_ASAP7_75t_L g11795 ( 
.A1(n_11025),
.A2(n_1550),
.B(n_1551),
.Y(n_11795)
);

OAI21x1_ASAP7_75t_L g11796 ( 
.A1(n_10749),
.A2(n_1552),
.B(n_1554),
.Y(n_11796)
);

AO31x2_ASAP7_75t_L g11797 ( 
.A1(n_10750),
.A2(n_1556),
.A3(n_1554),
.B(n_1555),
.Y(n_11797)
);

NAND2xp5_ASAP7_75t_L g11798 ( 
.A(n_11067),
.B(n_1555),
.Y(n_11798)
);

INVxp67_ASAP7_75t_SL g11799 ( 
.A(n_11197),
.Y(n_11799)
);

AOI22xp5_ASAP7_75t_L g11800 ( 
.A1(n_10897),
.A2(n_1558),
.B1(n_1556),
.B2(n_1557),
.Y(n_11800)
);

AND2x2_ASAP7_75t_L g11801 ( 
.A(n_10893),
.B(n_10913),
.Y(n_11801)
);

AOI21xp5_ASAP7_75t_L g11802 ( 
.A1(n_11223),
.A2(n_1557),
.B(n_1558),
.Y(n_11802)
);

OAI21x1_ASAP7_75t_L g11803 ( 
.A1(n_11070),
.A2(n_1559),
.B(n_1560),
.Y(n_11803)
);

AOI21x1_ASAP7_75t_L g11804 ( 
.A1(n_10970),
.A2(n_1559),
.B(n_1561),
.Y(n_11804)
);

OAI21xp5_ASAP7_75t_L g11805 ( 
.A1(n_11117),
.A2(n_1561),
.B(n_1562),
.Y(n_11805)
);

AOI21xp5_ASAP7_75t_SL g11806 ( 
.A1(n_10777),
.A2(n_10806),
.B(n_11175),
.Y(n_11806)
);

OAI22xp5_ASAP7_75t_L g11807 ( 
.A1(n_10583),
.A2(n_1565),
.B1(n_1562),
.B2(n_1564),
.Y(n_11807)
);

OAI21x1_ASAP7_75t_L g11808 ( 
.A1(n_10969),
.A2(n_1566),
.B(n_1567),
.Y(n_11808)
);

OAI22xp5_ASAP7_75t_L g11809 ( 
.A1(n_11037),
.A2(n_11185),
.B1(n_10849),
.B2(n_11018),
.Y(n_11809)
);

INVx2_ASAP7_75t_L g11810 ( 
.A(n_10962),
.Y(n_11810)
);

AOI21xp5_ASAP7_75t_L g11811 ( 
.A1(n_11228),
.A2(n_1568),
.B(n_1569),
.Y(n_11811)
);

INVx3_ASAP7_75t_L g11812 ( 
.A(n_10759),
.Y(n_11812)
);

AND2x4_ASAP7_75t_L g11813 ( 
.A(n_10776),
.B(n_1568),
.Y(n_11813)
);

INVx1_ASAP7_75t_L g11814 ( 
.A(n_10999),
.Y(n_11814)
);

AO21x2_ASAP7_75t_L g11815 ( 
.A1(n_11076),
.A2(n_1569),
.B(n_1570),
.Y(n_11815)
);

NAND2x1_ASAP7_75t_L g11816 ( 
.A(n_10793),
.B(n_1570),
.Y(n_11816)
);

INVx1_ASAP7_75t_L g11817 ( 
.A(n_11027),
.Y(n_11817)
);

AOI21xp5_ASAP7_75t_L g11818 ( 
.A1(n_10865),
.A2(n_11167),
.B(n_11209),
.Y(n_11818)
);

BUFx3_ASAP7_75t_L g11819 ( 
.A(n_10755),
.Y(n_11819)
);

AOI21x1_ASAP7_75t_L g11820 ( 
.A1(n_10994),
.A2(n_1571),
.B(n_1572),
.Y(n_11820)
);

BUFx4f_ASAP7_75t_L g11821 ( 
.A(n_10860),
.Y(n_11821)
);

NAND2xp5_ASAP7_75t_L g11822 ( 
.A(n_11083),
.B(n_1571),
.Y(n_11822)
);

NAND2x1p5_ASAP7_75t_L g11823 ( 
.A(n_10760),
.B(n_1572),
.Y(n_11823)
);

OAI21xp5_ASAP7_75t_L g11824 ( 
.A1(n_11135),
.A2(n_1573),
.B(n_1575),
.Y(n_11824)
);

AO31x2_ASAP7_75t_L g11825 ( 
.A1(n_11049),
.A2(n_1577),
.A3(n_1575),
.B(n_1576),
.Y(n_11825)
);

OAI21x1_ASAP7_75t_SL g11826 ( 
.A1(n_10966),
.A2(n_1577),
.B(n_1578),
.Y(n_11826)
);

INVx4_ASAP7_75t_L g11827 ( 
.A(n_10760),
.Y(n_11827)
);

NAND2xp5_ASAP7_75t_L g11828 ( 
.A(n_10817),
.B(n_1578),
.Y(n_11828)
);

OR2x2_ASAP7_75t_L g11829 ( 
.A(n_11113),
.B(n_1579),
.Y(n_11829)
);

BUFx2_ASAP7_75t_L g11830 ( 
.A(n_10785),
.Y(n_11830)
);

NAND2xp5_ASAP7_75t_L g11831 ( 
.A(n_10978),
.B(n_1579),
.Y(n_11831)
);

NAND2xp5_ASAP7_75t_L g11832 ( 
.A(n_10984),
.B(n_1580),
.Y(n_11832)
);

OAI21x1_ASAP7_75t_L g11833 ( 
.A1(n_11169),
.A2(n_1581),
.B(n_1582),
.Y(n_11833)
);

A2O1A1Ixp33_ASAP7_75t_L g11834 ( 
.A1(n_10714),
.A2(n_1583),
.B(n_1581),
.C(n_1582),
.Y(n_11834)
);

AOI21xp5_ASAP7_75t_L g11835 ( 
.A1(n_10865),
.A2(n_1583),
.B(n_1584),
.Y(n_11835)
);

INVx1_ASAP7_75t_L g11836 ( 
.A(n_11069),
.Y(n_11836)
);

NAND2x1p5_ASAP7_75t_L g11837 ( 
.A(n_10785),
.B(n_10882),
.Y(n_11837)
);

OAI21xp5_ASAP7_75t_SL g11838 ( 
.A1(n_11073),
.A2(n_1584),
.B(n_1585),
.Y(n_11838)
);

AND2x2_ASAP7_75t_L g11839 ( 
.A(n_10943),
.B(n_1585),
.Y(n_11839)
);

NAND2xp33_ASAP7_75t_L g11840 ( 
.A(n_11008),
.B(n_1586),
.Y(n_11840)
);

NOR2xp33_ASAP7_75t_L g11841 ( 
.A(n_10784),
.B(n_1586),
.Y(n_11841)
);

INVx1_ASAP7_75t_L g11842 ( 
.A(n_10751),
.Y(n_11842)
);

INVx1_ASAP7_75t_L g11843 ( 
.A(n_10751),
.Y(n_11843)
);

A2O1A1Ixp33_ASAP7_75t_L g11844 ( 
.A1(n_11110),
.A2(n_1589),
.B(n_1587),
.C(n_1588),
.Y(n_11844)
);

AO31x2_ASAP7_75t_L g11845 ( 
.A1(n_10912),
.A2(n_1589),
.A3(n_1587),
.B(n_1588),
.Y(n_11845)
);

INVxp67_ASAP7_75t_L g11846 ( 
.A(n_10839),
.Y(n_11846)
);

OAI21xp33_ASAP7_75t_L g11847 ( 
.A1(n_11177),
.A2(n_1590),
.B(n_1591),
.Y(n_11847)
);

AOI22x1_ASAP7_75t_L g11848 ( 
.A1(n_10656),
.A2(n_10657),
.B1(n_10670),
.B2(n_10664),
.Y(n_11848)
);

OAI22xp5_ASAP7_75t_L g11849 ( 
.A1(n_10568),
.A2(n_1592),
.B1(n_1590),
.B2(n_1591),
.Y(n_11849)
);

NAND2xp5_ASAP7_75t_L g11850 ( 
.A(n_10988),
.B(n_1592),
.Y(n_11850)
);

INVx1_ASAP7_75t_L g11851 ( 
.A(n_11199),
.Y(n_11851)
);

AOI21xp5_ASAP7_75t_L g11852 ( 
.A1(n_10867),
.A2(n_10682),
.B(n_10768),
.Y(n_11852)
);

OAI21x1_ASAP7_75t_L g11853 ( 
.A1(n_11233),
.A2(n_1593),
.B(n_1594),
.Y(n_11853)
);

AOI21xp5_ASAP7_75t_L g11854 ( 
.A1(n_10774),
.A2(n_1593),
.B(n_1594),
.Y(n_11854)
);

NAND2xp5_ASAP7_75t_L g11855 ( 
.A(n_11019),
.B(n_1595),
.Y(n_11855)
);

OAI21xp5_ASAP7_75t_L g11856 ( 
.A1(n_11181),
.A2(n_1595),
.B(n_1597),
.Y(n_11856)
);

INVx1_ASAP7_75t_L g11857 ( 
.A(n_11020),
.Y(n_11857)
);

OAI21x1_ASAP7_75t_L g11858 ( 
.A1(n_11089),
.A2(n_1598),
.B(n_1599),
.Y(n_11858)
);

OAI21x1_ASAP7_75t_L g11859 ( 
.A1(n_10673),
.A2(n_1598),
.B(n_1599),
.Y(n_11859)
);

OAI21x1_ASAP7_75t_L g11860 ( 
.A1(n_11023),
.A2(n_1600),
.B(n_1601),
.Y(n_11860)
);

A2O1A1Ixp33_ASAP7_75t_L g11861 ( 
.A1(n_11224),
.A2(n_1603),
.B(n_1601),
.C(n_1602),
.Y(n_11861)
);

AOI21xp5_ASAP7_75t_L g11862 ( 
.A1(n_10812),
.A2(n_10828),
.B(n_11137),
.Y(n_11862)
);

AOI221xp5_ASAP7_75t_L g11863 ( 
.A1(n_11187),
.A2(n_1605),
.B1(n_1603),
.B2(n_1604),
.C(n_1606),
.Y(n_11863)
);

AO31x2_ASAP7_75t_L g11864 ( 
.A1(n_11198),
.A2(n_1607),
.A3(n_1604),
.B(n_1605),
.Y(n_11864)
);

HB1xp67_ASAP7_75t_L g11865 ( 
.A(n_11039),
.Y(n_11865)
);

OR2x2_ASAP7_75t_L g11866 ( 
.A(n_10822),
.B(n_1607),
.Y(n_11866)
);

OAI21xp5_ASAP7_75t_L g11867 ( 
.A1(n_11026),
.A2(n_1608),
.B(n_1609),
.Y(n_11867)
);

AND2x4_ASAP7_75t_L g11868 ( 
.A(n_10658),
.B(n_1608),
.Y(n_11868)
);

NAND2xp5_ASAP7_75t_L g11869 ( 
.A(n_10824),
.B(n_1609),
.Y(n_11869)
);

OAI21x1_ASAP7_75t_L g11870 ( 
.A1(n_11186),
.A2(n_1610),
.B(n_1611),
.Y(n_11870)
);

OAI21x1_ASAP7_75t_L g11871 ( 
.A1(n_11194),
.A2(n_1610),
.B(n_1611),
.Y(n_11871)
);

AOI21x1_ASAP7_75t_L g11872 ( 
.A1(n_10729),
.A2(n_1612),
.B(n_1613),
.Y(n_11872)
);

INVx1_ASAP7_75t_L g11873 ( 
.A(n_11129),
.Y(n_11873)
);

OAI21x1_ASAP7_75t_L g11874 ( 
.A1(n_10769),
.A2(n_1612),
.B(n_1614),
.Y(n_11874)
);

OAI21x1_ASAP7_75t_L g11875 ( 
.A1(n_11221),
.A2(n_1615),
.B(n_1616),
.Y(n_11875)
);

AND2x2_ASAP7_75t_L g11876 ( 
.A(n_10975),
.B(n_1615),
.Y(n_11876)
);

AND2x2_ASAP7_75t_L g11877 ( 
.A(n_11030),
.B(n_1616),
.Y(n_11877)
);

OAI21x1_ASAP7_75t_L g11878 ( 
.A1(n_11214),
.A2(n_1617),
.B(n_1618),
.Y(n_11878)
);

NAND2x1_ASAP7_75t_L g11879 ( 
.A(n_10601),
.B(n_1618),
.Y(n_11879)
);

NOR2xp33_ASAP7_75t_L g11880 ( 
.A(n_10809),
.B(n_1619),
.Y(n_11880)
);

AO32x2_ASAP7_75t_L g11881 ( 
.A1(n_10688),
.A2(n_1621),
.A3(n_1619),
.B1(n_1620),
.B2(n_1622),
.Y(n_11881)
);

NAND2xp5_ASAP7_75t_L g11882 ( 
.A(n_10844),
.B(n_1620),
.Y(n_11882)
);

AND2x2_ASAP7_75t_L g11883 ( 
.A(n_11044),
.B(n_1621),
.Y(n_11883)
);

INVx3_ASAP7_75t_L g11884 ( 
.A(n_10641),
.Y(n_11884)
);

OAI22xp5_ASAP7_75t_L g11885 ( 
.A1(n_11251),
.A2(n_1624),
.B1(n_1622),
.B2(n_1623),
.Y(n_11885)
);

NAND2xp5_ASAP7_75t_L g11886 ( 
.A(n_11842),
.B(n_10856),
.Y(n_11886)
);

BUFx2_ASAP7_75t_L g11887 ( 
.A(n_11465),
.Y(n_11887)
);

INVx2_ASAP7_75t_L g11888 ( 
.A(n_11718),
.Y(n_11888)
);

BUFx3_ASAP7_75t_L g11889 ( 
.A(n_11297),
.Y(n_11889)
);

BUFx3_ASAP7_75t_L g11890 ( 
.A(n_11298),
.Y(n_11890)
);

OAI21x1_ASAP7_75t_L g11891 ( 
.A1(n_11315),
.A2(n_11032),
.B(n_10876),
.Y(n_11891)
);

AOI21x1_ASAP7_75t_L g11892 ( 
.A1(n_11625),
.A2(n_10886),
.B(n_10875),
.Y(n_11892)
);

OAI21xp5_ASAP7_75t_L g11893 ( 
.A1(n_11617),
.A2(n_11153),
.B(n_10979),
.Y(n_11893)
);

INVx1_ASAP7_75t_L g11894 ( 
.A(n_11718),
.Y(n_11894)
);

BUFx12f_ASAP7_75t_L g11895 ( 
.A(n_11392),
.Y(n_11895)
);

BUFx4f_ASAP7_75t_SL g11896 ( 
.A(n_11466),
.Y(n_11896)
);

AO21x2_ASAP7_75t_L g11897 ( 
.A1(n_11666),
.A2(n_10904),
.B(n_10896),
.Y(n_11897)
);

OR2x2_ASAP7_75t_L g11898 ( 
.A(n_11344),
.B(n_11136),
.Y(n_11898)
);

BUFx10_ASAP7_75t_L g11899 ( 
.A(n_11688),
.Y(n_11899)
);

INVx1_ASAP7_75t_L g11900 ( 
.A(n_11558),
.Y(n_11900)
);

OAI21x1_ASAP7_75t_L g11901 ( 
.A1(n_11444),
.A2(n_10917),
.B(n_10914),
.Y(n_11901)
);

AOI21xp5_ASAP7_75t_L g11902 ( 
.A1(n_11806),
.A2(n_11236),
.B(n_10981),
.Y(n_11902)
);

BUFx3_ASAP7_75t_L g11903 ( 
.A(n_11465),
.Y(n_11903)
);

OAI21x1_ASAP7_75t_L g11904 ( 
.A1(n_11708),
.A2(n_10930),
.B(n_10924),
.Y(n_11904)
);

OAI21x1_ASAP7_75t_L g11905 ( 
.A1(n_11408),
.A2(n_10933),
.B(n_11146),
.Y(n_11905)
);

OAI21x1_ASAP7_75t_L g11906 ( 
.A1(n_11391),
.A2(n_10961),
.B(n_11189),
.Y(n_11906)
);

AOI22x1_ASAP7_75t_L g11907 ( 
.A1(n_11521),
.A2(n_10936),
.B1(n_11188),
.B2(n_10940),
.Y(n_11907)
);

AND2x2_ASAP7_75t_L g11908 ( 
.A(n_11317),
.B(n_11063),
.Y(n_11908)
);

AND2x4_ASAP7_75t_L g11909 ( 
.A(n_11347),
.B(n_11179),
.Y(n_11909)
);

INVx2_ASAP7_75t_L g11910 ( 
.A(n_11453),
.Y(n_11910)
);

BUFx2_ASAP7_75t_SL g11911 ( 
.A(n_11496),
.Y(n_11911)
);

INVx2_ASAP7_75t_L g11912 ( 
.A(n_11462),
.Y(n_11912)
);

INVx2_ASAP7_75t_L g11913 ( 
.A(n_11480),
.Y(n_11913)
);

AO21x2_ASAP7_75t_L g11914 ( 
.A1(n_11373),
.A2(n_11150),
.B(n_11066),
.Y(n_11914)
);

OAI21xp5_ASAP7_75t_L g11915 ( 
.A1(n_11291),
.A2(n_11142),
.B(n_11126),
.Y(n_11915)
);

INVx1_ASAP7_75t_SL g11916 ( 
.A(n_11322),
.Y(n_11916)
);

AOI22xp5_ASAP7_75t_L g11917 ( 
.A1(n_11341),
.A2(n_11098),
.B1(n_11021),
.B2(n_10974),
.Y(n_11917)
);

OAI21x1_ASAP7_75t_L g11918 ( 
.A1(n_11473),
.A2(n_11200),
.B(n_11218),
.Y(n_11918)
);

AND2x2_ASAP7_75t_L g11919 ( 
.A(n_11419),
.B(n_11118),
.Y(n_11919)
);

AO21x2_ASAP7_75t_L g11920 ( 
.A1(n_11843),
.A2(n_11159),
.B(n_11101),
.Y(n_11920)
);

CKINVDCx5p33_ASAP7_75t_R g11921 ( 
.A(n_11380),
.Y(n_11921)
);

OAI21x1_ASAP7_75t_L g11922 ( 
.A1(n_11524),
.A2(n_10677),
.B(n_10672),
.Y(n_11922)
);

OAI21x1_ASAP7_75t_L g11923 ( 
.A1(n_11382),
.A2(n_11132),
.B(n_10778),
.Y(n_11923)
);

AOI22x1_ASAP7_75t_L g11924 ( 
.A1(n_11630),
.A2(n_10915),
.B1(n_11183),
.B2(n_11179),
.Y(n_11924)
);

OAI21x1_ASAP7_75t_L g11925 ( 
.A1(n_11799),
.A2(n_10663),
.B(n_11227),
.Y(n_11925)
);

CKINVDCx16_ASAP7_75t_R g11926 ( 
.A(n_11517),
.Y(n_11926)
);

OAI21x1_ASAP7_75t_L g11927 ( 
.A1(n_11563),
.A2(n_11237),
.B(n_11220),
.Y(n_11927)
);

INVx1_ASAP7_75t_L g11928 ( 
.A(n_11319),
.Y(n_11928)
);

OAI21x1_ASAP7_75t_L g11929 ( 
.A1(n_11570),
.A2(n_11326),
.B(n_11399),
.Y(n_11929)
);

AO21x2_ASAP7_75t_L g11930 ( 
.A1(n_11857),
.A2(n_11157),
.B(n_11079),
.Y(n_11930)
);

AOI21xp5_ASAP7_75t_L g11931 ( 
.A1(n_11564),
.A2(n_11158),
.B(n_11121),
.Y(n_11931)
);

INVx3_ASAP7_75t_L g11932 ( 
.A(n_11420),
.Y(n_11932)
);

BUFx6f_ASAP7_75t_L g11933 ( 
.A(n_11307),
.Y(n_11933)
);

INVx1_ASAP7_75t_L g11934 ( 
.A(n_11381),
.Y(n_11934)
);

INVx3_ASAP7_75t_L g11935 ( 
.A(n_11434),
.Y(n_11935)
);

OAI21x1_ASAP7_75t_L g11936 ( 
.A1(n_11730),
.A2(n_10632),
.B(n_10625),
.Y(n_11936)
);

INVx1_ASAP7_75t_L g11937 ( 
.A(n_11422),
.Y(n_11937)
);

AOI22xp33_ASAP7_75t_L g11938 ( 
.A1(n_11593),
.A2(n_11098),
.B1(n_11226),
.B2(n_10989),
.Y(n_11938)
);

INVx1_ASAP7_75t_L g11939 ( 
.A(n_11432),
.Y(n_11939)
);

AND2x2_ASAP7_75t_L g11940 ( 
.A(n_11450),
.B(n_10992),
.Y(n_11940)
);

CKINVDCx5p33_ASAP7_75t_R g11941 ( 
.A(n_11544),
.Y(n_11941)
);

OA21x2_ASAP7_75t_L g11942 ( 
.A1(n_11470),
.A2(n_11252),
.B(n_10590),
.Y(n_11942)
);

NOR2xp33_ASAP7_75t_SL g11943 ( 
.A(n_11750),
.B(n_10868),
.Y(n_11943)
);

INVx3_ASAP7_75t_L g11944 ( 
.A(n_11571),
.Y(n_11944)
);

INVx1_ASAP7_75t_L g11945 ( 
.A(n_11448),
.Y(n_11945)
);

NAND2x1p5_ASAP7_75t_L g11946 ( 
.A(n_11481),
.B(n_11183),
.Y(n_11946)
);

BUFx3_ASAP7_75t_L g11947 ( 
.A(n_11519),
.Y(n_11947)
);

OAI21x1_ASAP7_75t_L g11948 ( 
.A1(n_11425),
.A2(n_10846),
.B(n_11005),
.Y(n_11948)
);

HB1xp67_ASAP7_75t_L g11949 ( 
.A(n_11339),
.Y(n_11949)
);

CKINVDCx16_ASAP7_75t_R g11950 ( 
.A(n_11760),
.Y(n_11950)
);

BUFx3_ASAP7_75t_L g11951 ( 
.A(n_11498),
.Y(n_11951)
);

INVx1_ASAP7_75t_L g11952 ( 
.A(n_11479),
.Y(n_11952)
);

AO21x1_ASAP7_75t_L g11953 ( 
.A1(n_11580),
.A2(n_11442),
.B(n_11357),
.Y(n_11953)
);

INVx1_ASAP7_75t_L g11954 ( 
.A(n_11483),
.Y(n_11954)
);

OR2x2_ASAP7_75t_L g11955 ( 
.A(n_11337),
.B(n_10960),
.Y(n_11955)
);

OAI21x1_ASAP7_75t_L g11956 ( 
.A1(n_11513),
.A2(n_11508),
.B(n_11397),
.Y(n_11956)
);

BUFx6f_ASAP7_75t_L g11957 ( 
.A(n_11461),
.Y(n_11957)
);

INVx2_ASAP7_75t_L g11958 ( 
.A(n_11562),
.Y(n_11958)
);

OAI21x1_ASAP7_75t_L g11959 ( 
.A1(n_11687),
.A2(n_11281),
.B(n_10707),
.Y(n_11959)
);

BUFx3_ASAP7_75t_L g11960 ( 
.A(n_11821),
.Y(n_11960)
);

INVx1_ASAP7_75t_L g11961 ( 
.A(n_11584),
.Y(n_11961)
);

INVx1_ASAP7_75t_L g11962 ( 
.A(n_11604),
.Y(n_11962)
);

BUFx2_ASAP7_75t_SL g11963 ( 
.A(n_11464),
.Y(n_11963)
);

OA21x2_ASAP7_75t_L g11964 ( 
.A1(n_11478),
.A2(n_10713),
.B(n_10679),
.Y(n_11964)
);

AOI21xp5_ASAP7_75t_L g11965 ( 
.A1(n_11505),
.A2(n_10722),
.B(n_10862),
.Y(n_11965)
);

AOI21x1_ASAP7_75t_L g11966 ( 
.A1(n_11865),
.A2(n_11196),
.B(n_11180),
.Y(n_11966)
);

INVx1_ASAP7_75t_L g11967 ( 
.A(n_11632),
.Y(n_11967)
);

CKINVDCx20_ASAP7_75t_R g11968 ( 
.A(n_11692),
.Y(n_11968)
);

BUFx8_ASAP7_75t_L g11969 ( 
.A(n_11768),
.Y(n_11969)
);

CKINVDCx20_ASAP7_75t_R g11970 ( 
.A(n_11756),
.Y(n_11970)
);

BUFx6f_ASAP7_75t_L g11971 ( 
.A(n_11461),
.Y(n_11971)
);

INVx1_ASAP7_75t_L g11972 ( 
.A(n_11640),
.Y(n_11972)
);

BUFx4f_ASAP7_75t_L g11973 ( 
.A(n_11555),
.Y(n_11973)
);

INVx5_ASAP7_75t_L g11974 ( 
.A(n_11333),
.Y(n_11974)
);

INVx1_ASAP7_75t_L g11975 ( 
.A(n_11642),
.Y(n_11975)
);

INVx1_ASAP7_75t_L g11976 ( 
.A(n_11650),
.Y(n_11976)
);

NAND2xp5_ASAP7_75t_L g11977 ( 
.A(n_11354),
.B(n_11098),
.Y(n_11977)
);

NAND2x1p5_ASAP7_75t_L g11978 ( 
.A(n_11481),
.B(n_10915),
.Y(n_11978)
);

INVx3_ASAP7_75t_L g11979 ( 
.A(n_11499),
.Y(n_11979)
);

BUFx2_ASAP7_75t_SL g11980 ( 
.A(n_11445),
.Y(n_11980)
);

BUFx12f_ASAP7_75t_L g11981 ( 
.A(n_11404),
.Y(n_11981)
);

BUFx3_ASAP7_75t_L g11982 ( 
.A(n_11495),
.Y(n_11982)
);

BUFx8_ASAP7_75t_SL g11983 ( 
.A(n_11404),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_11654),
.Y(n_11984)
);

AND2x4_ASAP7_75t_L g11985 ( 
.A(n_11385),
.B(n_10740),
.Y(n_11985)
);

INVx2_ASAP7_75t_L g11986 ( 
.A(n_11588),
.Y(n_11986)
);

INVx1_ASAP7_75t_L g11987 ( 
.A(n_11668),
.Y(n_11987)
);

INVx2_ASAP7_75t_SL g11988 ( 
.A(n_11652),
.Y(n_11988)
);

INVx1_ASAP7_75t_L g11989 ( 
.A(n_11689),
.Y(n_11989)
);

AOI21x1_ASAP7_75t_L g11990 ( 
.A1(n_11510),
.A2(n_11191),
.B(n_11007),
.Y(n_11990)
);

INVx1_ASAP7_75t_L g11991 ( 
.A(n_11695),
.Y(n_11991)
);

OAI21x1_ASAP7_75t_L g11992 ( 
.A1(n_11754),
.A2(n_11217),
.B(n_10754),
.Y(n_11992)
);

BUFx2_ASAP7_75t_L g11993 ( 
.A(n_11752),
.Y(n_11993)
);

INVx1_ASAP7_75t_L g11994 ( 
.A(n_11697),
.Y(n_11994)
);

INVx1_ASAP7_75t_L g11995 ( 
.A(n_11704),
.Y(n_11995)
);

AND2x4_ASAP7_75t_L g11996 ( 
.A(n_11661),
.B(n_11095),
.Y(n_11996)
);

CKINVDCx20_ASAP7_75t_R g11997 ( 
.A(n_11819),
.Y(n_11997)
);

INVx1_ASAP7_75t_L g11998 ( 
.A(n_11731),
.Y(n_11998)
);

INVx1_ASAP7_75t_L g11999 ( 
.A(n_11741),
.Y(n_11999)
);

INVx5_ASAP7_75t_L g12000 ( 
.A(n_11333),
.Y(n_12000)
);

NOR2xp33_ASAP7_75t_L g12001 ( 
.A(n_11626),
.B(n_10957),
.Y(n_12001)
);

OAI21x1_ASAP7_75t_L g12002 ( 
.A1(n_11316),
.A2(n_11154),
.B(n_11017),
.Y(n_12002)
);

BUFx2_ASAP7_75t_L g12003 ( 
.A(n_11727),
.Y(n_12003)
);

INVx2_ASAP7_75t_SL g12004 ( 
.A(n_11497),
.Y(n_12004)
);

NAND2x1p5_ASAP7_75t_L g12005 ( 
.A(n_11557),
.B(n_1623),
.Y(n_12005)
);

HB1xp67_ASAP7_75t_L g12006 ( 
.A(n_11873),
.Y(n_12006)
);

INVx1_ASAP7_75t_L g12007 ( 
.A(n_11565),
.Y(n_12007)
);

NOR2xp33_ASAP7_75t_L g12008 ( 
.A(n_11567),
.B(n_10879),
.Y(n_12008)
);

INVx2_ASAP7_75t_SL g12009 ( 
.A(n_11348),
.Y(n_12009)
);

INVx4_ASAP7_75t_L g12010 ( 
.A(n_11411),
.Y(n_12010)
);

NAND2xp5_ASAP7_75t_L g12011 ( 
.A(n_11846),
.B(n_1624),
.Y(n_12011)
);

NAND2x1p5_ASAP7_75t_L g12012 ( 
.A(n_11557),
.B(n_1625),
.Y(n_12012)
);

OR2x2_ASAP7_75t_L g12013 ( 
.A(n_11851),
.B(n_11726),
.Y(n_12013)
);

OAI21x1_ASAP7_75t_L g12014 ( 
.A1(n_11503),
.A2(n_1626),
.B(n_1627),
.Y(n_12014)
);

INVxp67_ASAP7_75t_SL g12015 ( 
.A(n_11463),
.Y(n_12015)
);

CKINVDCx16_ASAP7_75t_R g12016 ( 
.A(n_11568),
.Y(n_12016)
);

AND2x2_ASAP7_75t_L g12017 ( 
.A(n_11801),
.B(n_1626),
.Y(n_12017)
);

CKINVDCx16_ASAP7_75t_R g12018 ( 
.A(n_11490),
.Y(n_12018)
);

BUFx2_ASAP7_75t_L g12019 ( 
.A(n_11830),
.Y(n_12019)
);

NOR2xp67_ASAP7_75t_SL g12020 ( 
.A(n_11311),
.B(n_1628),
.Y(n_12020)
);

INVx3_ASAP7_75t_L g12021 ( 
.A(n_11528),
.Y(n_12021)
);

OAI21x1_ASAP7_75t_L g12022 ( 
.A1(n_11477),
.A2(n_1628),
.B(n_1629),
.Y(n_12022)
);

OR2x6_ASAP7_75t_L g12023 ( 
.A(n_11411),
.B(n_1630),
.Y(n_12023)
);

INVx2_ASAP7_75t_L g12024 ( 
.A(n_11620),
.Y(n_12024)
);

OAI21xp5_ASAP7_75t_L g12025 ( 
.A1(n_11634),
.A2(n_1631),
.B(n_1632),
.Y(n_12025)
);

NAND2xp5_ASAP7_75t_SL g12026 ( 
.A(n_11628),
.B(n_1631),
.Y(n_12026)
);

BUFx6f_ASAP7_75t_L g12027 ( 
.A(n_11628),
.Y(n_12027)
);

INVx1_ASAP7_75t_L g12028 ( 
.A(n_11755),
.Y(n_12028)
);

NOR2xp33_ASAP7_75t_L g12029 ( 
.A(n_11653),
.B(n_1632),
.Y(n_12029)
);

INVx1_ASAP7_75t_L g12030 ( 
.A(n_11757),
.Y(n_12030)
);

OAI21x1_ASAP7_75t_L g12031 ( 
.A1(n_11407),
.A2(n_1633),
.B(n_1634),
.Y(n_12031)
);

INVx3_ASAP7_75t_L g12032 ( 
.A(n_11647),
.Y(n_12032)
);

AND2x4_ASAP7_75t_L g12033 ( 
.A(n_11313),
.B(n_1633),
.Y(n_12033)
);

INVx1_ASAP7_75t_L g12034 ( 
.A(n_11814),
.Y(n_12034)
);

OAI21x1_ASAP7_75t_L g12035 ( 
.A1(n_11758),
.A2(n_1634),
.B(n_1635),
.Y(n_12035)
);

INVx3_ASAP7_75t_SL g12036 ( 
.A(n_11523),
.Y(n_12036)
);

BUFx6f_ASAP7_75t_SL g12037 ( 
.A(n_11868),
.Y(n_12037)
);

HB1xp67_ASAP7_75t_L g12038 ( 
.A(n_11305),
.Y(n_12038)
);

INVx1_ASAP7_75t_L g12039 ( 
.A(n_11817),
.Y(n_12039)
);

INVx1_ASAP7_75t_L g12040 ( 
.A(n_11742),
.Y(n_12040)
);

INVxp67_ASAP7_75t_SL g12041 ( 
.A(n_11306),
.Y(n_12041)
);

OAI21x1_ASAP7_75t_L g12042 ( 
.A1(n_11327),
.A2(n_1635),
.B(n_1636),
.Y(n_12042)
);

BUFx6f_ASAP7_75t_L g12043 ( 
.A(n_11701),
.Y(n_12043)
);

HB1xp67_ASAP7_75t_L g12044 ( 
.A(n_11518),
.Y(n_12044)
);

AO21x2_ASAP7_75t_L g12045 ( 
.A1(n_11300),
.A2(n_1637),
.B(n_1638),
.Y(n_12045)
);

INVx2_ASAP7_75t_L g12046 ( 
.A(n_11810),
.Y(n_12046)
);

BUFx3_ASAP7_75t_L g12047 ( 
.A(n_11335),
.Y(n_12047)
);

BUFx3_ASAP7_75t_L g12048 ( 
.A(n_11335),
.Y(n_12048)
);

INVx3_ASAP7_75t_L g12049 ( 
.A(n_11662),
.Y(n_12049)
);

AO21x2_ASAP7_75t_L g12050 ( 
.A1(n_11390),
.A2(n_1639),
.B(n_1640),
.Y(n_12050)
);

BUFx12f_ASAP7_75t_L g12051 ( 
.A(n_11560),
.Y(n_12051)
);

BUFx2_ASAP7_75t_L g12052 ( 
.A(n_11740),
.Y(n_12052)
);

AND2x2_ASAP7_75t_L g12053 ( 
.A(n_11884),
.B(n_1639),
.Y(n_12053)
);

OAI21xp5_ASAP7_75t_L g12054 ( 
.A1(n_11841),
.A2(n_1640),
.B(n_1641),
.Y(n_12054)
);

INVx2_ASAP7_75t_L g12055 ( 
.A(n_11836),
.Y(n_12055)
);

INVx8_ASAP7_75t_L g12056 ( 
.A(n_11367),
.Y(n_12056)
);

BUFx3_ASAP7_75t_L g12057 ( 
.A(n_11367),
.Y(n_12057)
);

OAI21x1_ASAP7_75t_L g12058 ( 
.A1(n_11409),
.A2(n_1641),
.B(n_1642),
.Y(n_12058)
);

OAI21x1_ASAP7_75t_L g12059 ( 
.A1(n_11412),
.A2(n_11879),
.B(n_11488),
.Y(n_12059)
);

INVxp67_ASAP7_75t_SL g12060 ( 
.A(n_11551),
.Y(n_12060)
);

BUFx3_ASAP7_75t_L g12061 ( 
.A(n_11582),
.Y(n_12061)
);

CKINVDCx20_ASAP7_75t_R g12062 ( 
.A(n_11791),
.Y(n_12062)
);

BUFx2_ASAP7_75t_L g12063 ( 
.A(n_11740),
.Y(n_12063)
);

INVx2_ASAP7_75t_SL g12064 ( 
.A(n_11723),
.Y(n_12064)
);

INVx2_ASAP7_75t_SL g12065 ( 
.A(n_11714),
.Y(n_12065)
);

OAI21x1_ASAP7_75t_L g12066 ( 
.A1(n_11484),
.A2(n_1643),
.B(n_1644),
.Y(n_12066)
);

INVx2_ASAP7_75t_L g12067 ( 
.A(n_11325),
.Y(n_12067)
);

AND2x2_ASAP7_75t_L g12068 ( 
.A(n_11712),
.B(n_1643),
.Y(n_12068)
);

OAI21xp5_ASAP7_75t_L g12069 ( 
.A1(n_11474),
.A2(n_1644),
.B(n_1645),
.Y(n_12069)
);

INVx1_ASAP7_75t_L g12070 ( 
.A(n_11747),
.Y(n_12070)
);

BUFx6f_ASAP7_75t_L g12071 ( 
.A(n_11701),
.Y(n_12071)
);

AND2x2_ASAP7_75t_L g12072 ( 
.A(n_11318),
.B(n_1645),
.Y(n_12072)
);

INVx1_ASAP7_75t_SL g12073 ( 
.A(n_11378),
.Y(n_12073)
);

INVx2_ASAP7_75t_SL g12074 ( 
.A(n_11746),
.Y(n_12074)
);

INVxp67_ASAP7_75t_SL g12075 ( 
.A(n_11590),
.Y(n_12075)
);

CKINVDCx8_ASAP7_75t_R g12076 ( 
.A(n_11740),
.Y(n_12076)
);

OAI21x1_ASAP7_75t_L g12077 ( 
.A1(n_11501),
.A2(n_1646),
.B(n_1647),
.Y(n_12077)
);

OAI21x1_ASAP7_75t_L g12078 ( 
.A1(n_11334),
.A2(n_1646),
.B(n_1648),
.Y(n_12078)
);

OR2x2_ASAP7_75t_L g12079 ( 
.A(n_11360),
.B(n_1648),
.Y(n_12079)
);

NAND2xp5_ASAP7_75t_SL g12080 ( 
.A(n_11746),
.B(n_1649),
.Y(n_12080)
);

AND2x4_ASAP7_75t_L g12081 ( 
.A(n_11372),
.B(n_1649),
.Y(n_12081)
);

INVx5_ASAP7_75t_SL g12082 ( 
.A(n_11612),
.Y(n_12082)
);

AND2x4_ASAP7_75t_L g12083 ( 
.A(n_11402),
.B(n_1650),
.Y(n_12083)
);

AO21x2_ASAP7_75t_L g12084 ( 
.A1(n_11356),
.A2(n_1650),
.B(n_1651),
.Y(n_12084)
);

INVx3_ASAP7_75t_L g12085 ( 
.A(n_11827),
.Y(n_12085)
);

OAI21x1_ASAP7_75t_L g12086 ( 
.A1(n_11413),
.A2(n_11446),
.B(n_11292),
.Y(n_12086)
);

BUFx3_ASAP7_75t_L g12087 ( 
.A(n_11599),
.Y(n_12087)
);

AO21x2_ASAP7_75t_L g12088 ( 
.A1(n_11406),
.A2(n_1651),
.B(n_1652),
.Y(n_12088)
);

BUFx2_ASAP7_75t_R g12089 ( 
.A(n_11475),
.Y(n_12089)
);

INVx1_ASAP7_75t_L g12090 ( 
.A(n_11331),
.Y(n_12090)
);

AND2x2_ASAP7_75t_L g12091 ( 
.A(n_11706),
.B(n_1652),
.Y(n_12091)
);

BUFx3_ASAP7_75t_L g12092 ( 
.A(n_11611),
.Y(n_12092)
);

AND2x2_ASAP7_75t_L g12093 ( 
.A(n_11812),
.B(n_1653),
.Y(n_12093)
);

NAND2xp5_ASAP7_75t_L g12094 ( 
.A(n_11421),
.B(n_1653),
.Y(n_12094)
);

AO21x2_ASAP7_75t_L g12095 ( 
.A1(n_11418),
.A2(n_11438),
.B(n_11429),
.Y(n_12095)
);

HB1xp67_ASAP7_75t_L g12096 ( 
.A(n_11455),
.Y(n_12096)
);

OAI21x1_ASAP7_75t_L g12097 ( 
.A1(n_11504),
.A2(n_11520),
.B(n_11514),
.Y(n_12097)
);

OAI21x1_ASAP7_75t_L g12098 ( 
.A1(n_11527),
.A2(n_1654),
.B(n_1655),
.Y(n_12098)
);

NAND2xp5_ASAP7_75t_L g12099 ( 
.A(n_11375),
.B(n_1654),
.Y(n_12099)
);

BUFx8_ASAP7_75t_L g12100 ( 
.A(n_11371),
.Y(n_12100)
);

INVx2_ASAP7_75t_L g12101 ( 
.A(n_11437),
.Y(n_12101)
);

INVx3_ASAP7_75t_L g12102 ( 
.A(n_11351),
.Y(n_12102)
);

OAI21x1_ASAP7_75t_L g12103 ( 
.A1(n_11530),
.A2(n_1655),
.B(n_1656),
.Y(n_12103)
);

BUFx2_ASAP7_75t_L g12104 ( 
.A(n_11333),
.Y(n_12104)
);

OAI21x1_ASAP7_75t_L g12105 ( 
.A1(n_11531),
.A2(n_1656),
.B(n_1657),
.Y(n_12105)
);

BUFx3_ASAP7_75t_L g12106 ( 
.A(n_11542),
.Y(n_12106)
);

INVx1_ASAP7_75t_SL g12107 ( 
.A(n_11648),
.Y(n_12107)
);

INVx3_ASAP7_75t_L g12108 ( 
.A(n_11837),
.Y(n_12108)
);

INVx4_ASAP7_75t_L g12109 ( 
.A(n_11663),
.Y(n_12109)
);

OAI21x1_ASAP7_75t_L g12110 ( 
.A1(n_11537),
.A2(n_1657),
.B(n_1658),
.Y(n_12110)
);

OAI21xp5_ASAP7_75t_L g12111 ( 
.A1(n_11631),
.A2(n_1658),
.B(n_1659),
.Y(n_12111)
);

INVx2_ASAP7_75t_SL g12112 ( 
.A(n_11485),
.Y(n_12112)
);

NAND2xp5_ASAP7_75t_L g12113 ( 
.A(n_11388),
.B(n_1659),
.Y(n_12113)
);

OAI21x1_ASAP7_75t_L g12114 ( 
.A1(n_11539),
.A2(n_1660),
.B(n_1661),
.Y(n_12114)
);

OAI21x1_ASAP7_75t_L g12115 ( 
.A1(n_11321),
.A2(n_1660),
.B(n_1662),
.Y(n_12115)
);

BUFx6f_ASAP7_75t_L g12116 ( 
.A(n_11699),
.Y(n_12116)
);

BUFx6f_ASAP7_75t_L g12117 ( 
.A(n_11789),
.Y(n_12117)
);

OAI21x1_ASAP7_75t_L g12118 ( 
.A1(n_11338),
.A2(n_1662),
.B(n_1663),
.Y(n_12118)
);

CKINVDCx16_ASAP7_75t_R g12119 ( 
.A(n_11614),
.Y(n_12119)
);

INVx2_ASAP7_75t_SL g12120 ( 
.A(n_11494),
.Y(n_12120)
);

INVx2_ASAP7_75t_L g12121 ( 
.A(n_11455),
.Y(n_12121)
);

BUFx10_ASAP7_75t_L g12122 ( 
.A(n_11546),
.Y(n_12122)
);

BUFx6f_ASAP7_75t_L g12123 ( 
.A(n_11813),
.Y(n_12123)
);

OAI21xp5_ASAP7_75t_L g12124 ( 
.A1(n_11880),
.A2(n_1664),
.B(n_1665),
.Y(n_12124)
);

HB1xp67_ASAP7_75t_L g12125 ( 
.A(n_11469),
.Y(n_12125)
);

OAI21x1_ASAP7_75t_L g12126 ( 
.A1(n_11293),
.A2(n_11457),
.B(n_11314),
.Y(n_12126)
);

INVx1_ASAP7_75t_L g12127 ( 
.A(n_11331),
.Y(n_12127)
);

BUFx2_ASAP7_75t_L g12128 ( 
.A(n_11585),
.Y(n_12128)
);

BUFx4f_ASAP7_75t_SL g12129 ( 
.A(n_11839),
.Y(n_12129)
);

INVx2_ASAP7_75t_L g12130 ( 
.A(n_11301),
.Y(n_12130)
);

AND2x2_ASAP7_75t_L g12131 ( 
.A(n_11346),
.B(n_11387),
.Y(n_12131)
);

INVx2_ASAP7_75t_L g12132 ( 
.A(n_11301),
.Y(n_12132)
);

INVx1_ASAP7_75t_L g12133 ( 
.A(n_11329),
.Y(n_12133)
);

INVx2_ASAP7_75t_SL g12134 ( 
.A(n_11645),
.Y(n_12134)
);

INVx1_ASAP7_75t_L g12135 ( 
.A(n_11329),
.Y(n_12135)
);

AO21x2_ASAP7_75t_L g12136 ( 
.A1(n_11440),
.A2(n_1664),
.B(n_1665),
.Y(n_12136)
);

OAI21x1_ASAP7_75t_L g12137 ( 
.A1(n_11751),
.A2(n_1666),
.B(n_1667),
.Y(n_12137)
);

INVx1_ASAP7_75t_L g12138 ( 
.A(n_11459),
.Y(n_12138)
);

INVx4_ASAP7_75t_L g12139 ( 
.A(n_11534),
.Y(n_12139)
);

INVx1_ASAP7_75t_L g12140 ( 
.A(n_11541),
.Y(n_12140)
);

BUFx12f_ASAP7_75t_L g12141 ( 
.A(n_11735),
.Y(n_12141)
);

OAI21x1_ASAP7_75t_L g12142 ( 
.A1(n_11374),
.A2(n_1666),
.B(n_1668),
.Y(n_12142)
);

CKINVDCx20_ASAP7_75t_R g12143 ( 
.A(n_11876),
.Y(n_12143)
);

OAI21x1_ASAP7_75t_L g12144 ( 
.A1(n_11878),
.A2(n_11875),
.B(n_11290),
.Y(n_12144)
);

AND2x2_ASAP7_75t_L g12145 ( 
.A(n_11428),
.B(n_1669),
.Y(n_12145)
);

NAND2x1p5_ASAP7_75t_L g12146 ( 
.A(n_11492),
.B(n_11493),
.Y(n_12146)
);

OAI21xp5_ASAP7_75t_L g12147 ( 
.A1(n_11589),
.A2(n_1670),
.B(n_1671),
.Y(n_12147)
);

INVx3_ASAP7_75t_L g12148 ( 
.A(n_11673),
.Y(n_12148)
);

BUFx12f_ASAP7_75t_L g12149 ( 
.A(n_11355),
.Y(n_12149)
);

INVx1_ASAP7_75t_SL g12150 ( 
.A(n_11829),
.Y(n_12150)
);

CKINVDCx16_ASAP7_75t_R g12151 ( 
.A(n_11877),
.Y(n_12151)
);

AO21x2_ASAP7_75t_L g12152 ( 
.A1(n_11441),
.A2(n_1671),
.B(n_1672),
.Y(n_12152)
);

INVx3_ASAP7_75t_L g12153 ( 
.A(n_11786),
.Y(n_12153)
);

INVx4_ASAP7_75t_L g12154 ( 
.A(n_11602),
.Y(n_12154)
);

BUFx2_ASAP7_75t_R g12155 ( 
.A(n_11597),
.Y(n_12155)
);

OAI21xp5_ASAP7_75t_L g12156 ( 
.A1(n_11310),
.A2(n_1672),
.B(n_1673),
.Y(n_12156)
);

INVx1_ASAP7_75t_L g12157 ( 
.A(n_11553),
.Y(n_12157)
);

AND2x4_ASAP7_75t_L g12158 ( 
.A(n_11618),
.B(n_1673),
.Y(n_12158)
);

BUFx2_ASAP7_75t_SL g12159 ( 
.A(n_11883),
.Y(n_12159)
);

INVx1_ASAP7_75t_L g12160 ( 
.A(n_11312),
.Y(n_12160)
);

BUFx12f_ASAP7_75t_L g12161 ( 
.A(n_11394),
.Y(n_12161)
);

NAND2x1_ASAP7_75t_L g12162 ( 
.A(n_11299),
.B(n_1674),
.Y(n_12162)
);

NAND2x1p5_ASAP7_75t_L g12163 ( 
.A(n_11711),
.B(n_11476),
.Y(n_12163)
);

INVx3_ASAP7_75t_SL g12164 ( 
.A(n_11866),
.Y(n_12164)
);

INVx1_ASAP7_75t_L g12165 ( 
.A(n_11679),
.Y(n_12165)
);

NOR2xp33_ASAP7_75t_L g12166 ( 
.A(n_11540),
.B(n_11882),
.Y(n_12166)
);

AND2x2_ASAP7_75t_L g12167 ( 
.A(n_11509),
.B(n_1674),
.Y(n_12167)
);

AO21x2_ASAP7_75t_L g12168 ( 
.A1(n_11449),
.A2(n_1676),
.B(n_1677),
.Y(n_12168)
);

CKINVDCx5p33_ASAP7_75t_R g12169 ( 
.A(n_11743),
.Y(n_12169)
);

BUFx3_ASAP7_75t_L g12170 ( 
.A(n_11416),
.Y(n_12170)
);

NAND2x1p5_ASAP7_75t_L g12171 ( 
.A(n_11779),
.B(n_1676),
.Y(n_12171)
);

AO21x2_ASAP7_75t_L g12172 ( 
.A1(n_11587),
.A2(n_1677),
.B(n_1678),
.Y(n_12172)
);

BUFx2_ASAP7_75t_L g12173 ( 
.A(n_11516),
.Y(n_12173)
);

CKINVDCx20_ASAP7_75t_R g12174 ( 
.A(n_11716),
.Y(n_12174)
);

INVxp67_ASAP7_75t_L g12175 ( 
.A(n_11577),
.Y(n_12175)
);

INVx1_ASAP7_75t_SL g12176 ( 
.A(n_11526),
.Y(n_12176)
);

NAND2xp5_ASAP7_75t_L g12177 ( 
.A(n_11359),
.B(n_1679),
.Y(n_12177)
);

INVx1_ASAP7_75t_SL g12178 ( 
.A(n_11575),
.Y(n_12178)
);

BUFx2_ASAP7_75t_L g12179 ( 
.A(n_11709),
.Y(n_12179)
);

INVx1_ASAP7_75t_L g12180 ( 
.A(n_11679),
.Y(n_12180)
);

INVx1_ASAP7_75t_L g12181 ( 
.A(n_11452),
.Y(n_12181)
);

NAND2xp5_ASAP7_75t_L g12182 ( 
.A(n_11359),
.B(n_1680),
.Y(n_12182)
);

AO21x2_ASAP7_75t_L g12183 ( 
.A1(n_11826),
.A2(n_1680),
.B(n_1681),
.Y(n_12183)
);

INVx3_ASAP7_75t_L g12184 ( 
.A(n_11621),
.Y(n_12184)
);

INVx8_ASAP7_75t_L g12185 ( 
.A(n_11678),
.Y(n_12185)
);

OAI21x1_ASAP7_75t_L g12186 ( 
.A1(n_11320),
.A2(n_1681),
.B(n_1682),
.Y(n_12186)
);

OAI21x1_ASAP7_75t_L g12187 ( 
.A1(n_11349),
.A2(n_1682),
.B(n_1683),
.Y(n_12187)
);

AO21x2_ASAP7_75t_L g12188 ( 
.A1(n_11633),
.A2(n_1684),
.B(n_1685),
.Y(n_12188)
);

AND2x4_ASAP7_75t_L g12189 ( 
.A(n_11522),
.B(n_1684),
.Y(n_12189)
);

INVx1_ASAP7_75t_L g12190 ( 
.A(n_11452),
.Y(n_12190)
);

NAND2xp5_ASAP7_75t_L g12191 ( 
.A(n_11454),
.B(n_1685),
.Y(n_12191)
);

BUFx3_ASAP7_75t_L g12192 ( 
.A(n_11636),
.Y(n_12192)
);

AND2x2_ASAP7_75t_L g12193 ( 
.A(n_11761),
.B(n_1686),
.Y(n_12193)
);

OR2x6_ASAP7_75t_L g12194 ( 
.A(n_11816),
.B(n_1687),
.Y(n_12194)
);

INVx2_ASAP7_75t_L g12195 ( 
.A(n_11308),
.Y(n_12195)
);

INVx2_ASAP7_75t_SL g12196 ( 
.A(n_11655),
.Y(n_12196)
);

INVx1_ASAP7_75t_L g12197 ( 
.A(n_11533),
.Y(n_12197)
);

NAND2x1p5_ASAP7_75t_L g12198 ( 
.A(n_11532),
.B(n_1687),
.Y(n_12198)
);

INVx2_ASAP7_75t_L g12199 ( 
.A(n_11414),
.Y(n_12199)
);

BUFx2_ASAP7_75t_L g12200 ( 
.A(n_11815),
.Y(n_12200)
);

NOR2xp67_ASAP7_75t_L g12201 ( 
.A(n_11639),
.B(n_1688),
.Y(n_12201)
);

INVx4_ASAP7_75t_L g12202 ( 
.A(n_11780),
.Y(n_12202)
);

AO21x2_ASAP7_75t_L g12203 ( 
.A1(n_11581),
.A2(n_1688),
.B(n_1689),
.Y(n_12203)
);

OAI21x1_ASAP7_75t_L g12204 ( 
.A1(n_11302),
.A2(n_1689),
.B(n_1690),
.Y(n_12204)
);

INVx3_ASAP7_75t_L g12205 ( 
.A(n_11643),
.Y(n_12205)
);

AOI22x1_ASAP7_75t_L g12206 ( 
.A1(n_11770),
.A2(n_1693),
.B1(n_1691),
.B2(n_1692),
.Y(n_12206)
);

NAND2xp5_ASAP7_75t_L g12207 ( 
.A(n_11596),
.B(n_1692),
.Y(n_12207)
);

INVx1_ASAP7_75t_L g12208 ( 
.A(n_11533),
.Y(n_12208)
);

BUFx12f_ASAP7_75t_L g12209 ( 
.A(n_11823),
.Y(n_12209)
);

INVx1_ASAP7_75t_SL g12210 ( 
.A(n_11831),
.Y(n_12210)
);

AOI21x1_ASAP7_75t_L g12211 ( 
.A1(n_11606),
.A2(n_1693),
.B(n_1694),
.Y(n_12211)
);

OAI21xp5_ASAP7_75t_L g12212 ( 
.A1(n_11309),
.A2(n_1694),
.B(n_1695),
.Y(n_12212)
);

OAI21xp5_ASAP7_75t_L g12213 ( 
.A1(n_11426),
.A2(n_11323),
.B(n_11680),
.Y(n_12213)
);

INVx8_ASAP7_75t_L g12214 ( 
.A(n_11622),
.Y(n_12214)
);

HB1xp67_ASAP7_75t_L g12215 ( 
.A(n_11468),
.Y(n_12215)
);

INVx1_ASAP7_75t_L g12216 ( 
.A(n_11536),
.Y(n_12216)
);

AOI22x1_ASAP7_75t_L g12217 ( 
.A1(n_11818),
.A2(n_1697),
.B1(n_1695),
.B2(n_1696),
.Y(n_12217)
);

HB1xp67_ASAP7_75t_L g12218 ( 
.A(n_11468),
.Y(n_12218)
);

OAI21x1_ASAP7_75t_L g12219 ( 
.A1(n_11296),
.A2(n_1696),
.B(n_1697),
.Y(n_12219)
);

INVx1_ASAP7_75t_L g12220 ( 
.A(n_11536),
.Y(n_12220)
);

INVxp67_ASAP7_75t_SL g12221 ( 
.A(n_11615),
.Y(n_12221)
);

NAND2xp5_ASAP7_75t_L g12222 ( 
.A(n_11671),
.B(n_1698),
.Y(n_12222)
);

AOI22x1_ASAP7_75t_L g12223 ( 
.A1(n_11460),
.A2(n_11295),
.B1(n_11600),
.B2(n_11591),
.Y(n_12223)
);

NOR2xp33_ASAP7_75t_L g12224 ( 
.A(n_11832),
.B(n_1698),
.Y(n_12224)
);

INVx1_ASAP7_75t_SL g12225 ( 
.A(n_11850),
.Y(n_12225)
);

HB1xp67_ASAP7_75t_L g12226 ( 
.A(n_11549),
.Y(n_12226)
);

NAND2xp5_ASAP7_75t_L g12227 ( 
.A(n_11683),
.B(n_1700),
.Y(n_12227)
);

AO21x2_ASAP7_75t_L g12228 ( 
.A1(n_11482),
.A2(n_1700),
.B(n_1701),
.Y(n_12228)
);

AOI22x1_ASAP7_75t_L g12229 ( 
.A1(n_11862),
.A2(n_11500),
.B1(n_11443),
.B2(n_11576),
.Y(n_12229)
);

AO21x2_ASAP7_75t_L g12230 ( 
.A1(n_11748),
.A2(n_1702),
.B(n_1703),
.Y(n_12230)
);

INVx2_ASAP7_75t_L g12231 ( 
.A(n_11549),
.Y(n_12231)
);

CKINVDCx5p33_ASAP7_75t_R g12232 ( 
.A(n_11696),
.Y(n_12232)
);

NOR2xp33_ASAP7_75t_L g12233 ( 
.A(n_11855),
.B(n_1702),
.Y(n_12233)
);

INVx2_ASAP7_75t_L g12234 ( 
.A(n_11825),
.Y(n_12234)
);

HB1xp67_ASAP7_75t_L g12235 ( 
.A(n_11458),
.Y(n_12235)
);

INVx4_ASAP7_75t_L g12236 ( 
.A(n_11363),
.Y(n_12236)
);

BUFx4_ASAP7_75t_SL g12237 ( 
.A(n_11739),
.Y(n_12237)
);

CKINVDCx5p33_ASAP7_75t_R g12238 ( 
.A(n_11828),
.Y(n_12238)
);

BUFx8_ASAP7_75t_L g12239 ( 
.A(n_11881),
.Y(n_12239)
);

BUFx3_ASAP7_75t_L g12240 ( 
.A(n_11684),
.Y(n_12240)
);

OAI21x1_ASAP7_75t_L g12241 ( 
.A1(n_11793),
.A2(n_1704),
.B(n_1705),
.Y(n_12241)
);

INVxp67_ASAP7_75t_L g12242 ( 
.A(n_11769),
.Y(n_12242)
);

INVx1_ASAP7_75t_L g12243 ( 
.A(n_11825),
.Y(n_12243)
);

INVx3_ASAP7_75t_L g12244 ( 
.A(n_11487),
.Y(n_12244)
);

INVxp67_ASAP7_75t_SL g12245 ( 
.A(n_11574),
.Y(n_12245)
);

AO21x2_ASAP7_75t_L g12246 ( 
.A1(n_11773),
.A2(n_1706),
.B(n_1707),
.Y(n_12246)
);

NAND2xp5_ASAP7_75t_L g12247 ( 
.A(n_11787),
.B(n_1706),
.Y(n_12247)
);

HB1xp67_ASAP7_75t_L g12248 ( 
.A(n_11458),
.Y(n_12248)
);

INVx5_ASAP7_75t_L g12249 ( 
.A(n_11353),
.Y(n_12249)
);

INVx3_ASAP7_75t_L g12250 ( 
.A(n_11467),
.Y(n_12250)
);

INVx3_ASAP7_75t_L g12251 ( 
.A(n_11538),
.Y(n_12251)
);

INVx2_ASAP7_75t_SL g12252 ( 
.A(n_11609),
.Y(n_12252)
);

INVx1_ASAP7_75t_L g12253 ( 
.A(n_11395),
.Y(n_12253)
);

CKINVDCx5p33_ASAP7_75t_R g12254 ( 
.A(n_11869),
.Y(n_12254)
);

INVx3_ASAP7_75t_L g12255 ( 
.A(n_11389),
.Y(n_12255)
);

AOI22x1_ASAP7_75t_L g12256 ( 
.A1(n_11852),
.A2(n_1710),
.B1(n_1707),
.B2(n_1708),
.Y(n_12256)
);

INVx2_ASAP7_75t_L g12257 ( 
.A(n_11400),
.Y(n_12257)
);

OAI21xp5_ASAP7_75t_L g12258 ( 
.A1(n_11771),
.A2(n_1708),
.B(n_1710),
.Y(n_12258)
);

INVx5_ASAP7_75t_L g12259 ( 
.A(n_11433),
.Y(n_12259)
);

NAND2x1p5_ASAP7_75t_L g12260 ( 
.A(n_11379),
.B(n_1711),
.Y(n_12260)
);

HB1xp67_ASAP7_75t_L g12261 ( 
.A(n_11797),
.Y(n_12261)
);

HB1xp67_ASAP7_75t_L g12262 ( 
.A(n_11797),
.Y(n_12262)
);

OAI21x1_ASAP7_75t_L g12263 ( 
.A1(n_11556),
.A2(n_1711),
.B(n_1712),
.Y(n_12263)
);

INVx1_ASAP7_75t_L g12264 ( 
.A(n_11700),
.Y(n_12264)
);

BUFx2_ASAP7_75t_L g12265 ( 
.A(n_11693),
.Y(n_12265)
);

INVx1_ASAP7_75t_L g12266 ( 
.A(n_11736),
.Y(n_12266)
);

BUFx8_ASAP7_75t_L g12267 ( 
.A(n_11881),
.Y(n_12267)
);

INVx1_ASAP7_75t_L g12268 ( 
.A(n_11744),
.Y(n_12268)
);

OAI21x1_ASAP7_75t_SL g12269 ( 
.A1(n_11352),
.A2(n_1712),
.B(n_1713),
.Y(n_12269)
);

BUFx3_ASAP7_75t_L g12270 ( 
.A(n_11762),
.Y(n_12270)
);

INVx3_ASAP7_75t_L g12271 ( 
.A(n_11358),
.Y(n_12271)
);

INVx3_ASAP7_75t_SL g12272 ( 
.A(n_11383),
.Y(n_12272)
);

BUFx2_ASAP7_75t_L g12273 ( 
.A(n_11693),
.Y(n_12273)
);

OAI21x1_ASAP7_75t_L g12274 ( 
.A1(n_11607),
.A2(n_1713),
.B(n_1714),
.Y(n_12274)
);

AO21x1_ASAP7_75t_L g12275 ( 
.A1(n_11324),
.A2(n_1714),
.B(n_1715),
.Y(n_12275)
);

NAND2x1p5_ASAP7_75t_L g12276 ( 
.A(n_11627),
.B(n_1715),
.Y(n_12276)
);

NAND2x1p5_ASAP7_75t_L g12277 ( 
.A(n_11686),
.B(n_11694),
.Y(n_12277)
);

NOR2xp33_ASAP7_75t_L g12278 ( 
.A(n_11798),
.B(n_1716),
.Y(n_12278)
);

AO21x2_ASAP7_75t_L g12279 ( 
.A1(n_11822),
.A2(n_1716),
.B(n_1717),
.Y(n_12279)
);

HB1xp67_ASAP7_75t_L g12280 ( 
.A(n_11744),
.Y(n_12280)
);

OA21x2_ASAP7_75t_L g12281 ( 
.A1(n_11340),
.A2(n_1717),
.B(n_1718),
.Y(n_12281)
);

OAI21x1_ASAP7_75t_L g12282 ( 
.A1(n_11778),
.A2(n_1718),
.B(n_1719),
.Y(n_12282)
);

OAI21xp33_ASAP7_75t_L g12283 ( 
.A1(n_11578),
.A2(n_1719),
.B(n_1720),
.Y(n_12283)
);

NAND2xp5_ASAP7_75t_L g12284 ( 
.A(n_11366),
.B(n_1720),
.Y(n_12284)
);

INVx1_ASAP7_75t_L g12285 ( 
.A(n_11745),
.Y(n_12285)
);

AND2x2_ASAP7_75t_L g12286 ( 
.A(n_11566),
.B(n_1721),
.Y(n_12286)
);

BUFx3_ASAP7_75t_L g12287 ( 
.A(n_11675),
.Y(n_12287)
);

OAI21x1_ASAP7_75t_L g12288 ( 
.A1(n_11342),
.A2(n_1722),
.B(n_1723),
.Y(n_12288)
);

AO21x1_ASAP7_75t_L g12289 ( 
.A1(n_11336),
.A2(n_1722),
.B(n_1723),
.Y(n_12289)
);

OAI21x1_ASAP7_75t_L g12290 ( 
.A1(n_11665),
.A2(n_1724),
.B(n_1725),
.Y(n_12290)
);

AND2x2_ASAP7_75t_L g12291 ( 
.A(n_11566),
.B(n_1724),
.Y(n_12291)
);

AOI22x1_ASAP7_75t_L g12292 ( 
.A1(n_11489),
.A2(n_1727),
.B1(n_1725),
.B2(n_1726),
.Y(n_12292)
);

INVx1_ASAP7_75t_L g12293 ( 
.A(n_11745),
.Y(n_12293)
);

BUFx3_ASAP7_75t_L g12294 ( 
.A(n_11732),
.Y(n_12294)
);

OA21x2_ASAP7_75t_L g12295 ( 
.A1(n_11362),
.A2(n_1726),
.B(n_1727),
.Y(n_12295)
);

BUFx6f_ASAP7_75t_L g12296 ( 
.A(n_11749),
.Y(n_12296)
);

OAI21x1_ASAP7_75t_SL g12297 ( 
.A1(n_11838),
.A2(n_1728),
.B(n_1730),
.Y(n_12297)
);

BUFx3_ASAP7_75t_L g12298 ( 
.A(n_11803),
.Y(n_12298)
);

INVx1_ASAP7_75t_L g12299 ( 
.A(n_11529),
.Y(n_12299)
);

INVx3_ASAP7_75t_L g12300 ( 
.A(n_11804),
.Y(n_12300)
);

INVx5_ASAP7_75t_L g12301 ( 
.A(n_11328),
.Y(n_12301)
);

INVx2_ASAP7_75t_L g12302 ( 
.A(n_11403),
.Y(n_12302)
);

NOR2xp67_ASAP7_75t_L g12303 ( 
.A(n_11417),
.B(n_1730),
.Y(n_12303)
);

NAND2x1p5_ASAP7_75t_L g12304 ( 
.A(n_11707),
.B(n_1731),
.Y(n_12304)
);

BUFx6f_ASAP7_75t_L g12305 ( 
.A(n_11820),
.Y(n_12305)
);

AND2x4_ASAP7_75t_L g12306 ( 
.A(n_11772),
.B(n_1731),
.Y(n_12306)
);

INVx1_ASAP7_75t_L g12307 ( 
.A(n_11864),
.Y(n_12307)
);

BUFx2_ASAP7_75t_SL g12308 ( 
.A(n_11405),
.Y(n_12308)
);

INVx2_ASAP7_75t_L g12309 ( 
.A(n_11424),
.Y(n_12309)
);

OAI21x1_ASAP7_75t_L g12310 ( 
.A1(n_11717),
.A2(n_1732),
.B(n_1733),
.Y(n_12310)
);

INVx1_ASAP7_75t_L g12311 ( 
.A(n_11864),
.Y(n_12311)
);

BUFx6f_ASAP7_75t_L g12312 ( 
.A(n_11874),
.Y(n_12312)
);

INVx1_ASAP7_75t_L g12313 ( 
.A(n_11592),
.Y(n_12313)
);

INVx1_ASAP7_75t_SL g12314 ( 
.A(n_11376),
.Y(n_12314)
);

BUFx3_ASAP7_75t_L g12315 ( 
.A(n_11860),
.Y(n_12315)
);

OAI21x1_ASAP7_75t_L g12316 ( 
.A1(n_12121),
.A2(n_11765),
.B(n_11734),
.Y(n_12316)
);

AOI22xp33_ASAP7_75t_L g12317 ( 
.A1(n_12239),
.A2(n_11848),
.B1(n_11764),
.B2(n_11733),
.Y(n_12317)
);

AOI22xp33_ASAP7_75t_L g12318 ( 
.A1(n_12267),
.A2(n_11781),
.B1(n_11439),
.B2(n_11456),
.Y(n_12318)
);

OAI22xp5_ASAP7_75t_L g12319 ( 
.A1(n_12265),
.A2(n_11595),
.B1(n_11594),
.B2(n_11763),
.Y(n_12319)
);

OAI22xp5_ASAP7_75t_SL g12320 ( 
.A1(n_12273),
.A2(n_11753),
.B1(n_11550),
.B2(n_11809),
.Y(n_12320)
);

AO32x2_ASAP7_75t_L g12321 ( 
.A1(n_12196),
.A2(n_11525),
.A3(n_11289),
.B1(n_11681),
.B2(n_11674),
.Y(n_12321)
);

AOI22xp33_ASAP7_75t_L g12322 ( 
.A1(n_12249),
.A2(n_11637),
.B1(n_11824),
.B2(n_11805),
.Y(n_12322)
);

INVx2_ASAP7_75t_SL g12323 ( 
.A(n_11899),
.Y(n_12323)
);

OAI22xp5_ASAP7_75t_L g12324 ( 
.A1(n_12249),
.A2(n_12301),
.B1(n_12000),
.B2(n_11974),
.Y(n_12324)
);

BUFx2_ASAP7_75t_L g12325 ( 
.A(n_11887),
.Y(n_12325)
);

NAND2x1p5_ASAP7_75t_L g12326 ( 
.A(n_11974),
.B(n_11608),
.Y(n_12326)
);

OA21x2_ASAP7_75t_L g12327 ( 
.A1(n_11905),
.A2(n_11796),
.B(n_11808),
.Y(n_12327)
);

HB1xp67_ASAP7_75t_L g12328 ( 
.A(n_12125),
.Y(n_12328)
);

O2A1O1Ixp33_ASAP7_75t_SL g12329 ( 
.A1(n_12064),
.A2(n_11844),
.B(n_11605),
.C(n_11784),
.Y(n_12329)
);

OAI21xp5_ASAP7_75t_L g12330 ( 
.A1(n_11902),
.A2(n_11491),
.B(n_11545),
.Y(n_12330)
);

NAND2xp5_ASAP7_75t_L g12331 ( 
.A(n_12006),
.B(n_11847),
.Y(n_12331)
);

INVx2_ASAP7_75t_L g12332 ( 
.A(n_12315),
.Y(n_12332)
);

OAI21x1_ASAP7_75t_L g12333 ( 
.A1(n_11894),
.A2(n_11782),
.B(n_11303),
.Y(n_12333)
);

AND2x2_ASAP7_75t_L g12334 ( 
.A(n_12052),
.B(n_11610),
.Y(n_12334)
);

OAI21x1_ASAP7_75t_L g12335 ( 
.A1(n_11888),
.A2(n_11506),
.B(n_11872),
.Y(n_12335)
);

INVx2_ASAP7_75t_L g12336 ( 
.A(n_12255),
.Y(n_12336)
);

OAI21x1_ASAP7_75t_L g12337 ( 
.A1(n_12086),
.A2(n_11512),
.B(n_11330),
.Y(n_12337)
);

INVx1_ASAP7_75t_L g12338 ( 
.A(n_12090),
.Y(n_12338)
);

AOI22xp33_ASAP7_75t_SL g12339 ( 
.A1(n_12075),
.A2(n_11856),
.B1(n_11767),
.B2(n_11572),
.Y(n_12339)
);

NOR2x1_ASAP7_75t_R g12340 ( 
.A(n_11895),
.B(n_11840),
.Y(n_12340)
);

AOI22xp33_ASAP7_75t_L g12341 ( 
.A1(n_12223),
.A2(n_11759),
.B1(n_11603),
.B2(n_11613),
.Y(n_12341)
);

NAND2xp5_ASAP7_75t_L g12342 ( 
.A(n_11928),
.B(n_11610),
.Y(n_12342)
);

NAND3xp33_ASAP7_75t_L g12343 ( 
.A(n_12229),
.B(n_12096),
.C(n_12025),
.Y(n_12343)
);

AND2x2_ASAP7_75t_L g12344 ( 
.A(n_12063),
.B(n_11427),
.Y(n_12344)
);

BUFx3_ASAP7_75t_L g12345 ( 
.A(n_11890),
.Y(n_12345)
);

NAND2xp5_ASAP7_75t_L g12346 ( 
.A(n_12221),
.B(n_11592),
.Y(n_12346)
);

INVx1_ASAP7_75t_L g12347 ( 
.A(n_12127),
.Y(n_12347)
);

INVx1_ASAP7_75t_SL g12348 ( 
.A(n_12155),
.Y(n_12348)
);

OAI21x1_ASAP7_75t_L g12349 ( 
.A1(n_12195),
.A2(n_11435),
.B(n_11431),
.Y(n_12349)
);

OAI21x1_ASAP7_75t_L g12350 ( 
.A1(n_12130),
.A2(n_11447),
.B(n_11436),
.Y(n_12350)
);

INVx8_ASAP7_75t_L g12351 ( 
.A(n_12023),
.Y(n_12351)
);

AO21x2_ASAP7_75t_L g12352 ( 
.A1(n_12177),
.A2(n_11658),
.B(n_11573),
.Y(n_12352)
);

INVx1_ASAP7_75t_SL g12353 ( 
.A(n_11947),
.Y(n_12353)
);

NAND2xp5_ASAP7_75t_L g12354 ( 
.A(n_12095),
.B(n_11845),
.Y(n_12354)
);

OA21x2_ASAP7_75t_L g12355 ( 
.A1(n_12200),
.A2(n_11535),
.B(n_11835),
.Y(n_12355)
);

INVx1_ASAP7_75t_L g12356 ( 
.A(n_11934),
.Y(n_12356)
);

OAI21x1_ASAP7_75t_L g12357 ( 
.A1(n_12132),
.A2(n_11451),
.B(n_11471),
.Y(n_12357)
);

AO21x2_ASAP7_75t_L g12358 ( 
.A1(n_12182),
.A2(n_11423),
.B(n_11345),
.Y(n_12358)
);

OAI21x1_ASAP7_75t_L g12359 ( 
.A1(n_12244),
.A2(n_11472),
.B(n_11294),
.Y(n_12359)
);

OA21x2_ASAP7_75t_L g12360 ( 
.A1(n_11904),
.A2(n_11365),
.B(n_11332),
.Y(n_12360)
);

INVx2_ASAP7_75t_L g12361 ( 
.A(n_12205),
.Y(n_12361)
);

OAI21x1_ASAP7_75t_L g12362 ( 
.A1(n_12181),
.A2(n_11370),
.B(n_11368),
.Y(n_12362)
);

AOI21x1_ASAP7_75t_L g12363 ( 
.A1(n_11892),
.A2(n_11644),
.B(n_11624),
.Y(n_12363)
);

AO31x2_ASAP7_75t_L g12364 ( 
.A1(n_12236),
.A2(n_11430),
.A3(n_11861),
.B(n_11664),
.Y(n_12364)
);

INVx1_ASAP7_75t_L g12365 ( 
.A(n_11937),
.Y(n_12365)
);

INVx2_ASAP7_75t_L g12366 ( 
.A(n_12298),
.Y(n_12366)
);

OAI21x1_ASAP7_75t_L g12367 ( 
.A1(n_12190),
.A2(n_11398),
.B(n_11396),
.Y(n_12367)
);

OAI21x1_ASAP7_75t_L g12368 ( 
.A1(n_12313),
.A2(n_11350),
.B(n_11384),
.Y(n_12368)
);

AOI21xp5_ASAP7_75t_L g12369 ( 
.A1(n_12213),
.A2(n_11586),
.B(n_11719),
.Y(n_12369)
);

INVx1_ASAP7_75t_L g12370 ( 
.A(n_11939),
.Y(n_12370)
);

CKINVDCx5p33_ASAP7_75t_R g12371 ( 
.A(n_11941),
.Y(n_12371)
);

OAI211xp5_ASAP7_75t_SL g12372 ( 
.A1(n_11893),
.A2(n_11783),
.B(n_11386),
.C(n_11794),
.Y(n_12372)
);

AO31x2_ASAP7_75t_L g12373 ( 
.A1(n_12199),
.A2(n_11790),
.A3(n_11721),
.B(n_11776),
.Y(n_12373)
);

INVxp67_ASAP7_75t_SL g12374 ( 
.A(n_11942),
.Y(n_12374)
);

NOR2xp33_ASAP7_75t_L g12375 ( 
.A(n_11896),
.B(n_11677),
.Y(n_12375)
);

INVx2_ASAP7_75t_L g12376 ( 
.A(n_12251),
.Y(n_12376)
);

OAI21x1_ASAP7_75t_L g12377 ( 
.A1(n_11977),
.A2(n_11415),
.B(n_11547),
.Y(n_12377)
);

OAI21x1_ASAP7_75t_L g12378 ( 
.A1(n_12307),
.A2(n_11559),
.B(n_11554),
.Y(n_12378)
);

NOR2xp67_ASAP7_75t_L g12379 ( 
.A(n_12000),
.B(n_11698),
.Y(n_12379)
);

BUFx3_ASAP7_75t_L g12380 ( 
.A(n_11968),
.Y(n_12380)
);

AO31x2_ASAP7_75t_L g12381 ( 
.A1(n_12311),
.A2(n_11601),
.A3(n_11619),
.B(n_11552),
.Y(n_12381)
);

OAI21x1_ASAP7_75t_L g12382 ( 
.A1(n_12231),
.A2(n_11583),
.B(n_11561),
.Y(n_12382)
);

OAI21x1_ASAP7_75t_L g12383 ( 
.A1(n_12133),
.A2(n_11629),
.B(n_11598),
.Y(n_12383)
);

INVx2_ASAP7_75t_L g12384 ( 
.A(n_12250),
.Y(n_12384)
);

BUFx3_ASAP7_75t_L g12385 ( 
.A(n_11970),
.Y(n_12385)
);

INVx1_ASAP7_75t_L g12386 ( 
.A(n_12261),
.Y(n_12386)
);

OAI21x1_ASAP7_75t_L g12387 ( 
.A1(n_12135),
.A2(n_11649),
.B(n_11646),
.Y(n_12387)
);

INVx3_ASAP7_75t_L g12388 ( 
.A(n_11903),
.Y(n_12388)
);

AND2x2_ASAP7_75t_L g12389 ( 
.A(n_12019),
.B(n_11845),
.Y(n_12389)
);

AOI21xp5_ASAP7_75t_L g12390 ( 
.A1(n_12111),
.A2(n_11635),
.B(n_11548),
.Y(n_12390)
);

AOI21xp33_ASAP7_75t_SL g12391 ( 
.A1(n_11950),
.A2(n_11670),
.B(n_11579),
.Y(n_12391)
);

OAI21x1_ASAP7_75t_L g12392 ( 
.A1(n_12234),
.A2(n_11657),
.B(n_11656),
.Y(n_12392)
);

INVx1_ASAP7_75t_L g12393 ( 
.A(n_12262),
.Y(n_12393)
);

NAND2xp5_ASAP7_75t_L g12394 ( 
.A(n_12041),
.B(n_11486),
.Y(n_12394)
);

INVxp67_ASAP7_75t_L g12395 ( 
.A(n_11930),
.Y(n_12395)
);

AO21x2_ASAP7_75t_L g12396 ( 
.A1(n_11897),
.A2(n_11867),
.B(n_11788),
.Y(n_12396)
);

NAND2xp5_ASAP7_75t_L g12397 ( 
.A(n_12015),
.B(n_11486),
.Y(n_12397)
);

OA21x2_ASAP7_75t_L g12398 ( 
.A1(n_11901),
.A2(n_11638),
.B(n_11623),
.Y(n_12398)
);

OAI22xp5_ASAP7_75t_L g12399 ( 
.A1(n_12301),
.A2(n_11304),
.B1(n_11800),
.B2(n_11502),
.Y(n_12399)
);

AND2x4_ASAP7_75t_L g12400 ( 
.A(n_11951),
.B(n_11507),
.Y(n_12400)
);

AND2x2_ASAP7_75t_L g12401 ( 
.A(n_11993),
.B(n_11616),
.Y(n_12401)
);

HB1xp67_ASAP7_75t_L g12402 ( 
.A(n_11949),
.Y(n_12402)
);

AOI221xp5_ASAP7_75t_L g12403 ( 
.A1(n_12286),
.A2(n_11343),
.B1(n_11863),
.B2(n_11737),
.C(n_11738),
.Y(n_12403)
);

AO21x2_ASAP7_75t_L g12404 ( 
.A1(n_12291),
.A2(n_11569),
.B(n_11543),
.Y(n_12404)
);

INVx1_ASAP7_75t_SL g12405 ( 
.A(n_11926),
.Y(n_12405)
);

OAI21xp5_ASAP7_75t_L g12406 ( 
.A1(n_11915),
.A2(n_11393),
.B(n_11834),
.Y(n_12406)
);

AOI21xp5_ASAP7_75t_L g12407 ( 
.A1(n_12284),
.A2(n_11651),
.B(n_11641),
.Y(n_12407)
);

INVx1_ASAP7_75t_SL g12408 ( 
.A(n_11911),
.Y(n_12408)
);

NOR2xp33_ASAP7_75t_L g12409 ( 
.A(n_12073),
.B(n_11361),
.Y(n_12409)
);

NAND2xp5_ASAP7_75t_L g12410 ( 
.A(n_11920),
.B(n_11507),
.Y(n_12410)
);

INVx1_ASAP7_75t_L g12411 ( 
.A(n_12280),
.Y(n_12411)
);

AOI21xp33_ASAP7_75t_L g12412 ( 
.A1(n_12215),
.A2(n_11369),
.B(n_11807),
.Y(n_12412)
);

OAI21x1_ASAP7_75t_L g12413 ( 
.A1(n_11918),
.A2(n_11667),
.B(n_11659),
.Y(n_12413)
);

OAI21x1_ASAP7_75t_L g12414 ( 
.A1(n_12165),
.A2(n_12180),
.B(n_12268),
.Y(n_12414)
);

INVx1_ASAP7_75t_L g12415 ( 
.A(n_11961),
.Y(n_12415)
);

OAI21x1_ASAP7_75t_L g12416 ( 
.A1(n_12285),
.A2(n_11685),
.B(n_11672),
.Y(n_12416)
);

AOI221xp5_ASAP7_75t_L g12417 ( 
.A1(n_12253),
.A2(n_11729),
.B1(n_11710),
.B2(n_11669),
.C(n_11682),
.Y(n_12417)
);

INVx2_ASAP7_75t_L g12418 ( 
.A(n_12302),
.Y(n_12418)
);

OAI21xp33_ASAP7_75t_L g12419 ( 
.A1(n_12054),
.A2(n_11854),
.B(n_11660),
.Y(n_12419)
);

AO21x2_ASAP7_75t_L g12420 ( 
.A1(n_12293),
.A2(n_11702),
.B(n_11515),
.Y(n_12420)
);

AND2x4_ASAP7_75t_L g12421 ( 
.A(n_11996),
.B(n_11859),
.Y(n_12421)
);

O2A1O1Ixp33_ASAP7_75t_SL g12422 ( 
.A1(n_12112),
.A2(n_12120),
.B(n_11997),
.C(n_12080),
.Y(n_12422)
);

INVx4_ASAP7_75t_L g12423 ( 
.A(n_11889),
.Y(n_12423)
);

OAI21x1_ASAP7_75t_L g12424 ( 
.A1(n_11936),
.A2(n_11691),
.B(n_11690),
.Y(n_12424)
);

HB1xp67_ASAP7_75t_SL g12425 ( 
.A(n_12089),
.Y(n_12425)
);

BUFx2_ASAP7_75t_L g12426 ( 
.A(n_12003),
.Y(n_12426)
);

AND2x2_ASAP7_75t_L g12427 ( 
.A(n_11908),
.B(n_11616),
.Y(n_12427)
);

INVx2_ASAP7_75t_L g12428 ( 
.A(n_12309),
.Y(n_12428)
);

AOI22xp33_ASAP7_75t_L g12429 ( 
.A1(n_12308),
.A2(n_11511),
.B1(n_11728),
.B2(n_11715),
.Y(n_12429)
);

CKINVDCx5p33_ASAP7_75t_R g12430 ( 
.A(n_11921),
.Y(n_12430)
);

OR2x2_ASAP7_75t_L g12431 ( 
.A(n_11886),
.B(n_11766),
.Y(n_12431)
);

OAI21xp5_ASAP7_75t_L g12432 ( 
.A1(n_12126),
.A2(n_11410),
.B(n_11377),
.Y(n_12432)
);

INVx4_ASAP7_75t_L g12433 ( 
.A(n_11933),
.Y(n_12433)
);

AOI21xp33_ASAP7_75t_L g12434 ( 
.A1(n_12218),
.A2(n_11885),
.B(n_11849),
.Y(n_12434)
);

AND2x4_ASAP7_75t_L g12435 ( 
.A(n_11982),
.B(n_11870),
.Y(n_12435)
);

NAND2xp5_ASAP7_75t_L g12436 ( 
.A(n_12138),
.B(n_11676),
.Y(n_12436)
);

OAI21x1_ASAP7_75t_L g12437 ( 
.A1(n_12197),
.A2(n_11713),
.B(n_11703),
.Y(n_12437)
);

NAND2xp5_ASAP7_75t_L g12438 ( 
.A(n_12140),
.B(n_11676),
.Y(n_12438)
);

AND2x2_ASAP7_75t_L g12439 ( 
.A(n_11919),
.B(n_11766),
.Y(n_12439)
);

AND2x2_ASAP7_75t_L g12440 ( 
.A(n_11940),
.B(n_11871),
.Y(n_12440)
);

NOR2xp33_ASAP7_75t_L g12441 ( 
.A(n_12109),
.B(n_11364),
.Y(n_12441)
);

HB1xp67_ASAP7_75t_L g12442 ( 
.A(n_12038),
.Y(n_12442)
);

NAND2x1p5_ASAP7_75t_L g12443 ( 
.A(n_11973),
.B(n_11722),
.Y(n_12443)
);

OAI22xp33_ASAP7_75t_L g12444 ( 
.A1(n_12259),
.A2(n_11401),
.B1(n_11785),
.B2(n_11802),
.Y(n_12444)
);

AND2x2_ASAP7_75t_L g12445 ( 
.A(n_12153),
.B(n_11909),
.Y(n_12445)
);

INVx1_ASAP7_75t_L g12446 ( 
.A(n_11962),
.Y(n_12446)
);

OAI22xp5_ASAP7_75t_L g12447 ( 
.A1(n_12272),
.A2(n_11811),
.B1(n_11795),
.B2(n_11724),
.Y(n_12447)
);

INVx1_ASAP7_75t_L g12448 ( 
.A(n_11967),
.Y(n_12448)
);

INVx2_ASAP7_75t_L g12449 ( 
.A(n_12257),
.Y(n_12449)
);

NOR2xp33_ASAP7_75t_L g12450 ( 
.A(n_12018),
.B(n_11720),
.Y(n_12450)
);

AOI21xp5_ASAP7_75t_L g12451 ( 
.A1(n_11931),
.A2(n_11725),
.B(n_11705),
.Y(n_12451)
);

OAI21x1_ASAP7_75t_L g12452 ( 
.A1(n_12208),
.A2(n_11853),
.B(n_11833),
.Y(n_12452)
);

NAND2x1p5_ASAP7_75t_L g12453 ( 
.A(n_11979),
.B(n_11774),
.Y(n_12453)
);

OAI21x1_ASAP7_75t_L g12454 ( 
.A1(n_12216),
.A2(n_11858),
.B(n_11777),
.Y(n_12454)
);

AND2x2_ASAP7_75t_L g12455 ( 
.A(n_11944),
.B(n_11775),
.Y(n_12455)
);

OAI21xp5_ASAP7_75t_L g12456 ( 
.A1(n_12201),
.A2(n_11792),
.B(n_1732),
.Y(n_12456)
);

NOR2xp33_ASAP7_75t_L g12457 ( 
.A(n_12021),
.B(n_1733),
.Y(n_12457)
);

INVx3_ASAP7_75t_L g12458 ( 
.A(n_11983),
.Y(n_12458)
);

OAI21x1_ASAP7_75t_L g12459 ( 
.A1(n_12220),
.A2(n_1734),
.B(n_1735),
.Y(n_12459)
);

OAI21x1_ASAP7_75t_L g12460 ( 
.A1(n_12243),
.A2(n_1734),
.B(n_1735),
.Y(n_12460)
);

INVx1_ASAP7_75t_L g12461 ( 
.A(n_11972),
.Y(n_12461)
);

AOI21xp5_ASAP7_75t_L g12462 ( 
.A1(n_11914),
.A2(n_1736),
.B(n_1737),
.Y(n_12462)
);

BUFx2_ASAP7_75t_L g12463 ( 
.A(n_12062),
.Y(n_12463)
);

NAND2xp5_ASAP7_75t_L g12464 ( 
.A(n_12157),
.B(n_1737),
.Y(n_12464)
);

OAI21x1_ASAP7_75t_SL g12465 ( 
.A1(n_11953),
.A2(n_1738),
.B(n_1739),
.Y(n_12465)
);

HB1xp67_ASAP7_75t_L g12466 ( 
.A(n_11975),
.Y(n_12466)
);

OA21x2_ASAP7_75t_L g12467 ( 
.A1(n_12264),
.A2(n_1739),
.B(n_1741),
.Y(n_12467)
);

OAI21x1_ASAP7_75t_L g12468 ( 
.A1(n_11929),
.A2(n_1742),
.B(n_1743),
.Y(n_12468)
);

AND2x4_ASAP7_75t_L g12469 ( 
.A(n_11932),
.B(n_1742),
.Y(n_12469)
);

INVx2_ASAP7_75t_SL g12470 ( 
.A(n_12214),
.Y(n_12470)
);

AOI22xp33_ASAP7_75t_L g12471 ( 
.A1(n_12266),
.A2(n_1745),
.B1(n_1743),
.B2(n_1744),
.Y(n_12471)
);

OA21x2_ASAP7_75t_L g12472 ( 
.A1(n_11976),
.A2(n_1744),
.B(n_1745),
.Y(n_12472)
);

OAI22xp33_ASAP7_75t_L g12473 ( 
.A1(n_12259),
.A2(n_1748),
.B1(n_1746),
.B2(n_1747),
.Y(n_12473)
);

NAND2xp5_ASAP7_75t_L g12474 ( 
.A(n_12175),
.B(n_1746),
.Y(n_12474)
);

NOR2xp33_ASAP7_75t_L g12475 ( 
.A(n_12119),
.B(n_1747),
.Y(n_12475)
);

CKINVDCx5p33_ASAP7_75t_R g12476 ( 
.A(n_11963),
.Y(n_12476)
);

INVx1_ASAP7_75t_L g12477 ( 
.A(n_11984),
.Y(n_12477)
);

OAI21x1_ASAP7_75t_L g12478 ( 
.A1(n_11990),
.A2(n_1748),
.B(n_1749),
.Y(n_12478)
);

HB1xp67_ASAP7_75t_L g12479 ( 
.A(n_11987),
.Y(n_12479)
);

AND2x2_ASAP7_75t_L g12480 ( 
.A(n_12032),
.B(n_1750),
.Y(n_12480)
);

AOI21x1_ASAP7_75t_L g12481 ( 
.A1(n_12235),
.A2(n_1750),
.B(n_1751),
.Y(n_12481)
);

OAI21x1_ASAP7_75t_L g12482 ( 
.A1(n_11966),
.A2(n_1751),
.B(n_1753),
.Y(n_12482)
);

OAI21x1_ASAP7_75t_L g12483 ( 
.A1(n_12248),
.A2(n_1754),
.B(n_1755),
.Y(n_12483)
);

BUFx2_ASAP7_75t_L g12484 ( 
.A(n_12100),
.Y(n_12484)
);

AOI221x1_ASAP7_75t_L g12485 ( 
.A1(n_12001),
.A2(n_1756),
.B1(n_1754),
.B2(n_1755),
.C(n_1757),
.Y(n_12485)
);

INVx2_ASAP7_75t_L g12486 ( 
.A(n_12271),
.Y(n_12486)
);

INVx1_ASAP7_75t_L g12487 ( 
.A(n_11989),
.Y(n_12487)
);

OR2x6_ASAP7_75t_L g12488 ( 
.A(n_11978),
.B(n_1756),
.Y(n_12488)
);

AOI21x1_ASAP7_75t_L g12489 ( 
.A1(n_12104),
.A2(n_1758),
.B(n_1759),
.Y(n_12489)
);

AND2x2_ASAP7_75t_L g12490 ( 
.A(n_12049),
.B(n_1758),
.Y(n_12490)
);

OAI22xp5_ASAP7_75t_SL g12491 ( 
.A1(n_12151),
.A2(n_12129),
.B1(n_12016),
.B2(n_12143),
.Y(n_12491)
);

INVx2_ASAP7_75t_L g12492 ( 
.A(n_11910),
.Y(n_12492)
);

INVx1_ASAP7_75t_L g12493 ( 
.A(n_11991),
.Y(n_12493)
);

AND2x2_ASAP7_75t_L g12494 ( 
.A(n_12004),
.B(n_1759),
.Y(n_12494)
);

INVx1_ASAP7_75t_L g12495 ( 
.A(n_11994),
.Y(n_12495)
);

INVx1_ASAP7_75t_L g12496 ( 
.A(n_11995),
.Y(n_12496)
);

AO31x2_ASAP7_75t_L g12497 ( 
.A1(n_12179),
.A2(n_1762),
.A3(n_1760),
.B(n_1761),
.Y(n_12497)
);

HB1xp67_ASAP7_75t_L g12498 ( 
.A(n_11998),
.Y(n_12498)
);

INVx4_ASAP7_75t_L g12499 ( 
.A(n_11933),
.Y(n_12499)
);

OAI21x1_ASAP7_75t_L g12500 ( 
.A1(n_12226),
.A2(n_1761),
.B(n_1763),
.Y(n_12500)
);

OAI22xp5_ASAP7_75t_L g12501 ( 
.A1(n_11917),
.A2(n_1765),
.B1(n_1763),
.B2(n_1764),
.Y(n_12501)
);

BUFx3_ASAP7_75t_L g12502 ( 
.A(n_11969),
.Y(n_12502)
);

OAI21x1_ASAP7_75t_L g12503 ( 
.A1(n_11898),
.A2(n_1764),
.B(n_1765),
.Y(n_12503)
);

AO21x2_ASAP7_75t_L g12504 ( 
.A1(n_12011),
.A2(n_1766),
.B(n_1767),
.Y(n_12504)
);

OA21x2_ASAP7_75t_L g12505 ( 
.A1(n_11999),
.A2(n_11952),
.B(n_11945),
.Y(n_12505)
);

O2A1O1Ixp33_ASAP7_75t_L g12506 ( 
.A1(n_12124),
.A2(n_1768),
.B(n_1766),
.C(n_1767),
.Y(n_12506)
);

OAI21x1_ASAP7_75t_L g12507 ( 
.A1(n_12067),
.A2(n_1768),
.B(n_1769),
.Y(n_12507)
);

OAI21x1_ASAP7_75t_L g12508 ( 
.A1(n_11935),
.A2(n_1769),
.B(n_1770),
.Y(n_12508)
);

OAI21x1_ASAP7_75t_L g12509 ( 
.A1(n_11925),
.A2(n_1770),
.B(n_1771),
.Y(n_12509)
);

INVx8_ASAP7_75t_L g12510 ( 
.A(n_12056),
.Y(n_12510)
);

OA21x2_ASAP7_75t_L g12511 ( 
.A1(n_11954),
.A2(n_1771),
.B(n_1772),
.Y(n_12511)
);

HB1xp67_ASAP7_75t_L g12512 ( 
.A(n_11900),
.Y(n_12512)
);

OAI21x1_ASAP7_75t_L g12513 ( 
.A1(n_12184),
.A2(n_1772),
.B(n_1773),
.Y(n_12513)
);

OAI22xp33_ASAP7_75t_L g12514 ( 
.A1(n_12076),
.A2(n_12107),
.B1(n_12245),
.B2(n_11964),
.Y(n_12514)
);

AND2x4_ASAP7_75t_L g12515 ( 
.A(n_11988),
.B(n_1773),
.Y(n_12515)
);

BUFx12f_ASAP7_75t_L g12516 ( 
.A(n_12051),
.Y(n_12516)
);

OAI21x1_ASAP7_75t_L g12517 ( 
.A1(n_11891),
.A2(n_1774),
.B(n_1775),
.Y(n_12517)
);

AO21x2_ASAP7_75t_L g12518 ( 
.A1(n_12160),
.A2(n_1776),
.B(n_1777),
.Y(n_12518)
);

A2O1A1Ixp33_ASAP7_75t_L g12519 ( 
.A1(n_12283),
.A2(n_1780),
.B(n_1778),
.C(n_1779),
.Y(n_12519)
);

CKINVDCx5p33_ASAP7_75t_R g12520 ( 
.A(n_11980),
.Y(n_12520)
);

INVx2_ASAP7_75t_L g12521 ( 
.A(n_11912),
.Y(n_12521)
);

AND2x4_ASAP7_75t_L g12522 ( 
.A(n_12106),
.B(n_1778),
.Y(n_12522)
);

BUFx2_ASAP7_75t_SL g12523 ( 
.A(n_12037),
.Y(n_12523)
);

AO31x2_ASAP7_75t_L g12524 ( 
.A1(n_12173),
.A2(n_1782),
.A3(n_1780),
.B(n_1781),
.Y(n_12524)
);

AND2x4_ASAP7_75t_L g12525 ( 
.A(n_11985),
.B(n_1781),
.Y(n_12525)
);

OAI221xp5_ASAP7_75t_L g12526 ( 
.A1(n_12069),
.A2(n_1785),
.B1(n_1783),
.B2(n_1784),
.C(n_1786),
.Y(n_12526)
);

HB1xp67_ASAP7_75t_L g12527 ( 
.A(n_12242),
.Y(n_12527)
);

INVx2_ASAP7_75t_L g12528 ( 
.A(n_11913),
.Y(n_12528)
);

NOR2xp33_ASAP7_75t_L g12529 ( 
.A(n_12164),
.B(n_1783),
.Y(n_12529)
);

CKINVDCx5p33_ASAP7_75t_R g12530 ( 
.A(n_11960),
.Y(n_12530)
);

AOI222xp33_ASAP7_75t_L g12531 ( 
.A1(n_12147),
.A2(n_12156),
.B1(n_12082),
.B2(n_12303),
.C1(n_12191),
.C2(n_12306),
.Y(n_12531)
);

AO21x2_ASAP7_75t_L g12532 ( 
.A1(n_12094),
.A2(n_1785),
.B(n_1786),
.Y(n_12532)
);

CKINVDCx16_ASAP7_75t_R g12533 ( 
.A(n_11943),
.Y(n_12533)
);

BUFx2_ASAP7_75t_SL g12534 ( 
.A(n_12061),
.Y(n_12534)
);

OR2x2_ASAP7_75t_L g12535 ( 
.A(n_12150),
.B(n_1787),
.Y(n_12535)
);

INVx2_ASAP7_75t_L g12536 ( 
.A(n_11958),
.Y(n_12536)
);

NAND2xp5_ASAP7_75t_L g12537 ( 
.A(n_12210),
.B(n_1787),
.Y(n_12537)
);

AOI22xp33_ASAP7_75t_L g12538 ( 
.A1(n_12289),
.A2(n_1790),
.B1(n_1788),
.B2(n_1789),
.Y(n_12538)
);

AO21x2_ASAP7_75t_L g12539 ( 
.A1(n_12099),
.A2(n_1788),
.B(n_1789),
.Y(n_12539)
);

OA21x2_ASAP7_75t_L g12540 ( 
.A1(n_12028),
.A2(n_1791),
.B(n_1792),
.Y(n_12540)
);

OAI21xp5_ASAP7_75t_L g12541 ( 
.A1(n_12029),
.A2(n_1791),
.B(n_1792),
.Y(n_12541)
);

INVx3_ASAP7_75t_L g12542 ( 
.A(n_11981),
.Y(n_12542)
);

NAND2xp5_ASAP7_75t_L g12543 ( 
.A(n_12225),
.B(n_1793),
.Y(n_12543)
);

INVx6_ASAP7_75t_L g12544 ( 
.A(n_12117),
.Y(n_12544)
);

INVx1_ASAP7_75t_L g12545 ( 
.A(n_12030),
.Y(n_12545)
);

OAI21x1_ASAP7_75t_SL g12546 ( 
.A1(n_12134),
.A2(n_1794),
.B(n_1795),
.Y(n_12546)
);

INVx1_ASAP7_75t_L g12547 ( 
.A(n_12034),
.Y(n_12547)
);

OAI21x1_ASAP7_75t_L g12548 ( 
.A1(n_12300),
.A2(n_1794),
.B(n_1796),
.Y(n_12548)
);

A2O1A1Ixp33_ASAP7_75t_L g12549 ( 
.A1(n_12224),
.A2(n_1798),
.B(n_1796),
.C(n_1797),
.Y(n_12549)
);

A2O1A1Ixp33_ASAP7_75t_L g12550 ( 
.A1(n_12233),
.A2(n_1799),
.B(n_1797),
.C(n_1798),
.Y(n_12550)
);

AND2x4_ASAP7_75t_L g12551 ( 
.A(n_12148),
.B(n_1799),
.Y(n_12551)
);

NAND2x1p5_ASAP7_75t_L g12552 ( 
.A(n_11916),
.B(n_12010),
.Y(n_12552)
);

INVx1_ASAP7_75t_SL g12553 ( 
.A(n_12036),
.Y(n_12553)
);

AOI21x1_ASAP7_75t_L g12554 ( 
.A1(n_12162),
.A2(n_12128),
.B(n_12299),
.Y(n_12554)
);

HB1xp67_ASAP7_75t_L g12555 ( 
.A(n_12050),
.Y(n_12555)
);

OR2x2_ASAP7_75t_L g12556 ( 
.A(n_12044),
.B(n_1800),
.Y(n_12556)
);

O2A1O1Ixp33_ASAP7_75t_SL g12557 ( 
.A1(n_12026),
.A2(n_1802),
.B(n_1800),
.C(n_1801),
.Y(n_12557)
);

CKINVDCx6p67_ASAP7_75t_R g12558 ( 
.A(n_12141),
.Y(n_12558)
);

INVx3_ASAP7_75t_L g12559 ( 
.A(n_12117),
.Y(n_12559)
);

AOI21x1_ASAP7_75t_L g12560 ( 
.A1(n_12211),
.A2(n_1801),
.B(n_1803),
.Y(n_12560)
);

OAI21x1_ASAP7_75t_L g12561 ( 
.A1(n_12108),
.A2(n_12039),
.B(n_12070),
.Y(n_12561)
);

INVx2_ASAP7_75t_L g12562 ( 
.A(n_11986),
.Y(n_12562)
);

NAND2xp5_ASAP7_75t_L g12563 ( 
.A(n_12176),
.B(n_1803),
.Y(n_12563)
);

OR2x6_ASAP7_75t_L g12564 ( 
.A(n_12159),
.B(n_1804),
.Y(n_12564)
);

INVx2_ASAP7_75t_L g12565 ( 
.A(n_12024),
.Y(n_12565)
);

OAI22xp33_ASAP7_75t_L g12566 ( 
.A1(n_12087),
.A2(n_1806),
.B1(n_1804),
.B2(n_1805),
.Y(n_12566)
);

CKINVDCx16_ASAP7_75t_R g12567 ( 
.A(n_12149),
.Y(n_12567)
);

AOI22xp33_ASAP7_75t_L g12568 ( 
.A1(n_12217),
.A2(n_1808),
.B1(n_1806),
.B2(n_1807),
.Y(n_12568)
);

INVx1_ASAP7_75t_L g12569 ( 
.A(n_12007),
.Y(n_12569)
);

OAI21x1_ASAP7_75t_L g12570 ( 
.A1(n_11946),
.A2(n_1807),
.B(n_1809),
.Y(n_12570)
);

AOI22xp33_ASAP7_75t_L g12571 ( 
.A1(n_12228),
.A2(n_1811),
.B1(n_1809),
.B2(n_1810),
.Y(n_12571)
);

OAI21xp5_ASAP7_75t_L g12572 ( 
.A1(n_11948),
.A2(n_1810),
.B(n_1811),
.Y(n_12572)
);

HB1xp67_ASAP7_75t_L g12573 ( 
.A(n_12084),
.Y(n_12573)
);

AND2x2_ASAP7_75t_L g12574 ( 
.A(n_12065),
.B(n_1812),
.Y(n_12574)
);

BUFx3_ASAP7_75t_L g12575 ( 
.A(n_12092),
.Y(n_12575)
);

CKINVDCx5p33_ASAP7_75t_R g12576 ( 
.A(n_12047),
.Y(n_12576)
);

BUFx6f_ASAP7_75t_L g12577 ( 
.A(n_12209),
.Y(n_12577)
);

A2O1A1Ixp33_ASAP7_75t_L g12578 ( 
.A1(n_12278),
.A2(n_1814),
.B(n_1812),
.C(n_1813),
.Y(n_12578)
);

NAND3xp33_ASAP7_75t_L g12579 ( 
.A(n_11965),
.B(n_1813),
.C(n_1814),
.Y(n_12579)
);

INVx2_ASAP7_75t_L g12580 ( 
.A(n_12046),
.Y(n_12580)
);

OAI21x1_ASAP7_75t_L g12581 ( 
.A1(n_11955),
.A2(n_1815),
.B(n_1816),
.Y(n_12581)
);

OA21x2_ASAP7_75t_L g12582 ( 
.A1(n_12040),
.A2(n_12060),
.B(n_12055),
.Y(n_12582)
);

NOR2xp67_ASAP7_75t_SL g12583 ( 
.A(n_12161),
.B(n_1815),
.Y(n_12583)
);

NAND2xp5_ASAP7_75t_L g12584 ( 
.A(n_12166),
.B(n_1816),
.Y(n_12584)
);

AO31x2_ASAP7_75t_L g12585 ( 
.A1(n_12275),
.A2(n_1819),
.A3(n_1817),
.B(n_1818),
.Y(n_12585)
);

AND2x4_ASAP7_75t_L g12586 ( 
.A(n_12009),
.B(n_1817),
.Y(n_12586)
);

OAI22xp5_ASAP7_75t_L g12587 ( 
.A1(n_11938),
.A2(n_1820),
.B1(n_1818),
.B2(n_1819),
.Y(n_12587)
);

INVx1_ASAP7_75t_L g12588 ( 
.A(n_12013),
.Y(n_12588)
);

OAI21x1_ASAP7_75t_L g12589 ( 
.A1(n_12085),
.A2(n_1820),
.B(n_1821),
.Y(n_12589)
);

AOI22xp33_ASAP7_75t_L g12590 ( 
.A1(n_12305),
.A2(n_1823),
.B1(n_1821),
.B2(n_1822),
.Y(n_12590)
);

AND2x2_ASAP7_75t_L g12591 ( 
.A(n_12102),
.B(n_1823),
.Y(n_12591)
);

OAI21x1_ASAP7_75t_L g12592 ( 
.A1(n_12097),
.A2(n_1824),
.B(n_1825),
.Y(n_12592)
);

INVxp67_ASAP7_75t_L g12593 ( 
.A(n_12008),
.Y(n_12593)
);

OAI21x1_ASAP7_75t_SL g12594 ( 
.A1(n_12139),
.A2(n_1824),
.B(n_1825),
.Y(n_12594)
);

INVx6_ASAP7_75t_L g12595 ( 
.A(n_12123),
.Y(n_12595)
);

NAND2x1p5_ASAP7_75t_L g12596 ( 
.A(n_12116),
.B(n_1826),
.Y(n_12596)
);

AND2x2_ASAP7_75t_L g12597 ( 
.A(n_12074),
.B(n_1826),
.Y(n_12597)
);

AOI22xp33_ASAP7_75t_L g12598 ( 
.A1(n_12305),
.A2(n_1829),
.B1(n_1827),
.B2(n_1828),
.Y(n_12598)
);

OR2x6_ASAP7_75t_L g12599 ( 
.A(n_12185),
.B(n_12005),
.Y(n_12599)
);

AOI21xp33_ASAP7_75t_L g12600 ( 
.A1(n_12297),
.A2(n_1827),
.B(n_1830),
.Y(n_12600)
);

INVx2_ASAP7_75t_L g12601 ( 
.A(n_12312),
.Y(n_12601)
);

OAI22xp5_ASAP7_75t_L g12602 ( 
.A1(n_12277),
.A2(n_1833),
.B1(n_1831),
.B2(n_1832),
.Y(n_12602)
);

INVx2_ASAP7_75t_L g12603 ( 
.A(n_12312),
.Y(n_12603)
);

CKINVDCx20_ASAP7_75t_R g12604 ( 
.A(n_12174),
.Y(n_12604)
);

OAI21x1_ASAP7_75t_L g12605 ( 
.A1(n_11956),
.A2(n_1831),
.B(n_1832),
.Y(n_12605)
);

HB1xp67_ASAP7_75t_L g12606 ( 
.A(n_12230),
.Y(n_12606)
);

AO21x2_ASAP7_75t_L g12607 ( 
.A1(n_12113),
.A2(n_1834),
.B(n_1835),
.Y(n_12607)
);

OAI21x1_ASAP7_75t_L g12608 ( 
.A1(n_12059),
.A2(n_1835),
.B(n_1836),
.Y(n_12608)
);

NAND2x1p5_ASAP7_75t_L g12609 ( 
.A(n_12116),
.B(n_1836),
.Y(n_12609)
);

AO21x2_ASAP7_75t_L g12610 ( 
.A1(n_12207),
.A2(n_1837),
.B(n_1838),
.Y(n_12610)
);

OAI22xp5_ASAP7_75t_L g12611 ( 
.A1(n_12163),
.A2(n_1840),
.B1(n_1837),
.B2(n_1839),
.Y(n_12611)
);

OAI21x1_ASAP7_75t_L g12612 ( 
.A1(n_12146),
.A2(n_1841),
.B(n_1842),
.Y(n_12612)
);

NOR2xp67_ASAP7_75t_L g12613 ( 
.A(n_12154),
.B(n_1841),
.Y(n_12613)
);

OR2x2_ASAP7_75t_L g12614 ( 
.A(n_12178),
.B(n_12192),
.Y(n_12614)
);

OR2x2_ASAP7_75t_L g12615 ( 
.A(n_12131),
.B(n_12270),
.Y(n_12615)
);

BUFx3_ASAP7_75t_L g12616 ( 
.A(n_12123),
.Y(n_12616)
);

OAI21x1_ASAP7_75t_L g12617 ( 
.A1(n_12101),
.A2(n_1842),
.B(n_1843),
.Y(n_12617)
);

OAI21x1_ASAP7_75t_L g12618 ( 
.A1(n_12144),
.A2(n_1844),
.B(n_1845),
.Y(n_12618)
);

CKINVDCx20_ASAP7_75t_R g12619 ( 
.A(n_12048),
.Y(n_12619)
);

NAND2xp5_ASAP7_75t_L g12620 ( 
.A(n_12252),
.B(n_1844),
.Y(n_12620)
);

OAI21x1_ASAP7_75t_L g12621 ( 
.A1(n_11906),
.A2(n_1846),
.B(n_1847),
.Y(n_12621)
);

AOI22xp33_ASAP7_75t_L g12622 ( 
.A1(n_12020),
.A2(n_1849),
.B1(n_1846),
.B2(n_1848),
.Y(n_12622)
);

AO21x2_ASAP7_75t_L g12623 ( 
.A1(n_12222),
.A2(n_1848),
.B(n_1849),
.Y(n_12623)
);

AOI22xp33_ASAP7_75t_L g12624 ( 
.A1(n_12269),
.A2(n_1853),
.B1(n_1850),
.B2(n_1852),
.Y(n_12624)
);

AND2x4_ASAP7_75t_L g12625 ( 
.A(n_12240),
.B(n_1852),
.Y(n_12625)
);

OAI21x1_ASAP7_75t_L g12626 ( 
.A1(n_11924),
.A2(n_1853),
.B(n_1854),
.Y(n_12626)
);

AND2x2_ASAP7_75t_L g12627 ( 
.A(n_12057),
.B(n_12017),
.Y(n_12627)
);

OR2x2_ASAP7_75t_L g12628 ( 
.A(n_12079),
.B(n_1855),
.Y(n_12628)
);

AND2x4_ASAP7_75t_L g12629 ( 
.A(n_12287),
.B(n_1855),
.Y(n_12629)
);

OAI211xp5_ASAP7_75t_L g12630 ( 
.A1(n_12256),
.A2(n_1858),
.B(n_1856),
.C(n_1857),
.Y(n_12630)
);

BUFx12f_ASAP7_75t_L g12631 ( 
.A(n_12122),
.Y(n_12631)
);

INVx1_ASAP7_75t_SL g12632 ( 
.A(n_12232),
.Y(n_12632)
);

HB1xp67_ASAP7_75t_L g12633 ( 
.A(n_12172),
.Y(n_12633)
);

OA21x2_ASAP7_75t_L g12634 ( 
.A1(n_12169),
.A2(n_1856),
.B(n_1857),
.Y(n_12634)
);

HB1xp67_ASAP7_75t_L g12635 ( 
.A(n_12045),
.Y(n_12635)
);

OAI21x1_ASAP7_75t_L g12636 ( 
.A1(n_11907),
.A2(n_1858),
.B(n_1859),
.Y(n_12636)
);

BUFx2_ASAP7_75t_L g12637 ( 
.A(n_11957),
.Y(n_12637)
);

CKINVDCx5p33_ASAP7_75t_R g12638 ( 
.A(n_12238),
.Y(n_12638)
);

OR2x2_ASAP7_75t_L g12639 ( 
.A(n_12203),
.B(n_1859),
.Y(n_12639)
);

INVx1_ASAP7_75t_L g12640 ( 
.A(n_12088),
.Y(n_12640)
);

A2O1A1Ixp33_ASAP7_75t_L g12641 ( 
.A1(n_12258),
.A2(n_1862),
.B(n_1860),
.C(n_1861),
.Y(n_12641)
);

INVx2_ASAP7_75t_L g12642 ( 
.A(n_12136),
.Y(n_12642)
);

NOR2xp33_ASAP7_75t_L g12643 ( 
.A(n_12254),
.B(n_1861),
.Y(n_12643)
);

OR2x6_ASAP7_75t_L g12644 ( 
.A(n_12012),
.B(n_1862),
.Y(n_12644)
);

OA21x2_ASAP7_75t_L g12645 ( 
.A1(n_12227),
.A2(n_1864),
.B(n_1865),
.Y(n_12645)
);

INVx2_ASAP7_75t_SL g12646 ( 
.A(n_12296),
.Y(n_12646)
);

A2O1A1Ixp33_ASAP7_75t_L g12647 ( 
.A1(n_12212),
.A2(n_1866),
.B(n_1864),
.C(n_1865),
.Y(n_12647)
);

BUFx2_ASAP7_75t_L g12648 ( 
.A(n_11957),
.Y(n_12648)
);

OAI21x1_ASAP7_75t_L g12649 ( 
.A1(n_11922),
.A2(n_1866),
.B(n_1867),
.Y(n_12649)
);

INVx1_ASAP7_75t_L g12650 ( 
.A(n_12152),
.Y(n_12650)
);

CKINVDCx20_ASAP7_75t_R g12651 ( 
.A(n_12170),
.Y(n_12651)
);

OAI21x1_ASAP7_75t_L g12652 ( 
.A1(n_11959),
.A2(n_1867),
.B(n_1868),
.Y(n_12652)
);

BUFx6f_ASAP7_75t_L g12653 ( 
.A(n_11971),
.Y(n_12653)
);

OA21x2_ASAP7_75t_L g12654 ( 
.A1(n_12241),
.A2(n_1868),
.B(n_1869),
.Y(n_12654)
);

INVx1_ASAP7_75t_L g12655 ( 
.A(n_12168),
.Y(n_12655)
);

INVx1_ASAP7_75t_L g12656 ( 
.A(n_12246),
.Y(n_12656)
);

AO21x2_ASAP7_75t_L g12657 ( 
.A1(n_12247),
.A2(n_1870),
.B(n_1871),
.Y(n_12657)
);

INVx3_ASAP7_75t_L g12658 ( 
.A(n_12296),
.Y(n_12658)
);

OAI21xp5_ASAP7_75t_L g12659 ( 
.A1(n_11927),
.A2(n_1870),
.B(n_1871),
.Y(n_12659)
);

NOR2xp33_ASAP7_75t_L g12660 ( 
.A(n_12202),
.B(n_1872),
.Y(n_12660)
);

INVx1_ASAP7_75t_L g12661 ( 
.A(n_12279),
.Y(n_12661)
);

BUFx3_ASAP7_75t_L g12662 ( 
.A(n_12294),
.Y(n_12662)
);

AND2x4_ASAP7_75t_SL g12663 ( 
.A(n_11971),
.B(n_1872),
.Y(n_12663)
);

OAI21x1_ASAP7_75t_L g12664 ( 
.A1(n_12002),
.A2(n_1873),
.B(n_1874),
.Y(n_12664)
);

NOR2xp33_ASAP7_75t_R g12665 ( 
.A(n_12027),
.B(n_1873),
.Y(n_12665)
);

INVx1_ASAP7_75t_L g12666 ( 
.A(n_12188),
.Y(n_12666)
);

AOI22xp33_ASAP7_75t_SL g12667 ( 
.A1(n_12206),
.A2(n_1878),
.B1(n_1875),
.B2(n_1876),
.Y(n_12667)
);

AOI221xp5_ASAP7_75t_L g12668 ( 
.A1(n_12314),
.A2(n_1879),
.B1(n_1875),
.B2(n_1878),
.C(n_1880),
.Y(n_12668)
);

OAI21x1_ASAP7_75t_L g12669 ( 
.A1(n_12042),
.A2(n_1879),
.B(n_1880),
.Y(n_12669)
);

OAI21x1_ASAP7_75t_L g12670 ( 
.A1(n_12022),
.A2(n_1881),
.B(n_1882),
.Y(n_12670)
);

HB1xp67_ASAP7_75t_L g12671 ( 
.A(n_12053),
.Y(n_12671)
);

BUFx3_ASAP7_75t_L g12672 ( 
.A(n_12145),
.Y(n_12672)
);

OAI21x1_ASAP7_75t_L g12673 ( 
.A1(n_12263),
.A2(n_1883),
.B(n_1884),
.Y(n_12673)
);

BUFx12f_ASAP7_75t_L g12674 ( 
.A(n_12193),
.Y(n_12674)
);

INVx1_ASAP7_75t_L g12675 ( 
.A(n_12281),
.Y(n_12675)
);

OAI22xp33_ASAP7_75t_L g12676 ( 
.A1(n_12198),
.A2(n_1885),
.B1(n_1883),
.B2(n_1884),
.Y(n_12676)
);

INVx2_ASAP7_75t_L g12677 ( 
.A(n_12033),
.Y(n_12677)
);

AND2x4_ASAP7_75t_L g12678 ( 
.A(n_12027),
.B(n_1885),
.Y(n_12678)
);

INVx2_ASAP7_75t_L g12679 ( 
.A(n_12081),
.Y(n_12679)
);

INVx4_ASAP7_75t_L g12680 ( 
.A(n_12043),
.Y(n_12680)
);

AO31x2_ASAP7_75t_L g12681 ( 
.A1(n_12237),
.A2(n_1888),
.A3(n_1886),
.B(n_1887),
.Y(n_12681)
);

OA21x2_ASAP7_75t_L g12682 ( 
.A1(n_12068),
.A2(n_1886),
.B(n_1887),
.Y(n_12682)
);

OAI21x1_ASAP7_75t_L g12683 ( 
.A1(n_12274),
.A2(n_12282),
.B(n_12114),
.Y(n_12683)
);

INVx2_ASAP7_75t_SL g12684 ( 
.A(n_12043),
.Y(n_12684)
);

AOI21xp5_ASAP7_75t_L g12685 ( 
.A1(n_12183),
.A2(n_12189),
.B(n_12194),
.Y(n_12685)
);

OA21x2_ASAP7_75t_L g12686 ( 
.A1(n_12167),
.A2(n_1888),
.B(n_1889),
.Y(n_12686)
);

OAI211xp5_ASAP7_75t_L g12687 ( 
.A1(n_12292),
.A2(n_1892),
.B(n_1889),
.C(n_1891),
.Y(n_12687)
);

OA21x2_ASAP7_75t_L g12688 ( 
.A1(n_11923),
.A2(n_1892),
.B(n_1893),
.Y(n_12688)
);

OAI21x1_ASAP7_75t_SL g12689 ( 
.A1(n_12324),
.A2(n_12295),
.B(n_12171),
.Y(n_12689)
);

OAI21x1_ASAP7_75t_L g12690 ( 
.A1(n_12414),
.A2(n_12035),
.B(n_12072),
.Y(n_12690)
);

HB1xp67_ASAP7_75t_L g12691 ( 
.A(n_12402),
.Y(n_12691)
);

AOI21xp5_ASAP7_75t_L g12692 ( 
.A1(n_12462),
.A2(n_12260),
.B(n_12276),
.Y(n_12692)
);

INVx2_ASAP7_75t_L g12693 ( 
.A(n_12615),
.Y(n_12693)
);

OR2x2_ASAP7_75t_L g12694 ( 
.A(n_12442),
.B(n_12527),
.Y(n_12694)
);

CKINVDCx6p67_ASAP7_75t_R g12695 ( 
.A(n_12502),
.Y(n_12695)
);

INVx1_ASAP7_75t_L g12696 ( 
.A(n_12466),
.Y(n_12696)
);

INVx1_ASAP7_75t_L g12697 ( 
.A(n_12479),
.Y(n_12697)
);

AOI21xp5_ASAP7_75t_L g12698 ( 
.A1(n_12369),
.A2(n_12304),
.B(n_12158),
.Y(n_12698)
);

AND2x4_ASAP7_75t_L g12699 ( 
.A(n_12575),
.B(n_12083),
.Y(n_12699)
);

INVx1_ASAP7_75t_L g12700 ( 
.A(n_12498),
.Y(n_12700)
);

CKINVDCx5p33_ASAP7_75t_R g12701 ( 
.A(n_12430),
.Y(n_12701)
);

INVx2_ASAP7_75t_L g12702 ( 
.A(n_12453),
.Y(n_12702)
);

BUFx2_ASAP7_75t_R g12703 ( 
.A(n_12523),
.Y(n_12703)
);

INVx2_ASAP7_75t_L g12704 ( 
.A(n_12505),
.Y(n_12704)
);

INVx1_ASAP7_75t_L g12705 ( 
.A(n_12512),
.Y(n_12705)
);

INVx1_ASAP7_75t_L g12706 ( 
.A(n_12338),
.Y(n_12706)
);

OAI21x1_ASAP7_75t_L g12707 ( 
.A1(n_12561),
.A2(n_12014),
.B(n_11992),
.Y(n_12707)
);

INVx1_ASAP7_75t_L g12708 ( 
.A(n_12347),
.Y(n_12708)
);

OAI21xp5_ASAP7_75t_L g12709 ( 
.A1(n_12343),
.A2(n_12310),
.B(n_12290),
.Y(n_12709)
);

HB1xp67_ASAP7_75t_L g12710 ( 
.A(n_12675),
.Y(n_12710)
);

AOI21xp5_ASAP7_75t_L g12711 ( 
.A1(n_12319),
.A2(n_12091),
.B(n_12093),
.Y(n_12711)
);

CKINVDCx5p33_ASAP7_75t_R g12712 ( 
.A(n_12371),
.Y(n_12712)
);

INVx2_ASAP7_75t_L g12713 ( 
.A(n_12377),
.Y(n_12713)
);

INVx1_ASAP7_75t_L g12714 ( 
.A(n_12356),
.Y(n_12714)
);

AND2x2_ASAP7_75t_L g12715 ( 
.A(n_12344),
.B(n_12071),
.Y(n_12715)
);

OAI21x1_ASAP7_75t_L g12716 ( 
.A1(n_12342),
.A2(n_12077),
.B(n_12066),
.Y(n_12716)
);

OR2x2_ASAP7_75t_L g12717 ( 
.A(n_12588),
.B(n_12331),
.Y(n_12717)
);

AO21x2_ASAP7_75t_L g12718 ( 
.A1(n_12374),
.A2(n_12078),
.B(n_12058),
.Y(n_12718)
);

INVx1_ASAP7_75t_L g12719 ( 
.A(n_12365),
.Y(n_12719)
);

A2O1A1Ixp33_ASAP7_75t_L g12720 ( 
.A1(n_12330),
.A2(n_12098),
.B(n_12105),
.C(n_12103),
.Y(n_12720)
);

BUFx6f_ASAP7_75t_SL g12721 ( 
.A(n_12345),
.Y(n_12721)
);

NAND2xp5_ASAP7_75t_L g12722 ( 
.A(n_12396),
.B(n_12110),
.Y(n_12722)
);

AOI21xp33_ASAP7_75t_L g12723 ( 
.A1(n_12410),
.A2(n_12137),
.B(n_12031),
.Y(n_12723)
);

NAND2xp5_ASAP7_75t_L g12724 ( 
.A(n_12346),
.B(n_12071),
.Y(n_12724)
);

OAI21x1_ASAP7_75t_L g12725 ( 
.A1(n_12361),
.A2(n_12115),
.B(n_12118),
.Y(n_12725)
);

AOI21xp5_ASAP7_75t_L g12726 ( 
.A1(n_12320),
.A2(n_12219),
.B(n_12204),
.Y(n_12726)
);

AOI21xp33_ASAP7_75t_L g12727 ( 
.A1(n_12514),
.A2(n_12395),
.B(n_12354),
.Y(n_12727)
);

AND2x2_ASAP7_75t_L g12728 ( 
.A(n_12534),
.B(n_12325),
.Y(n_12728)
);

OA21x2_ASAP7_75t_L g12729 ( 
.A1(n_12593),
.A2(n_12186),
.B(n_12187),
.Y(n_12729)
);

AO31x2_ASAP7_75t_L g12730 ( 
.A1(n_12642),
.A2(n_12288),
.A3(n_12142),
.B(n_1895),
.Y(n_12730)
);

OR2x2_ASAP7_75t_L g12731 ( 
.A(n_12397),
.B(n_1893),
.Y(n_12731)
);

AND2x2_ASAP7_75t_L g12732 ( 
.A(n_12440),
.B(n_1894),
.Y(n_12732)
);

AOI21xp5_ASAP7_75t_L g12733 ( 
.A1(n_12322),
.A2(n_1894),
.B(n_1896),
.Y(n_12733)
);

BUFx4f_ASAP7_75t_SL g12734 ( 
.A(n_12516),
.Y(n_12734)
);

NAND2xp5_ASAP7_75t_L g12735 ( 
.A(n_12436),
.B(n_1896),
.Y(n_12735)
);

NOR2xp33_ASAP7_75t_L g12736 ( 
.A(n_12533),
.B(n_12425),
.Y(n_12736)
);

AND2x2_ASAP7_75t_L g12737 ( 
.A(n_12388),
.B(n_1897),
.Y(n_12737)
);

NAND2xp5_ASAP7_75t_L g12738 ( 
.A(n_12438),
.B(n_1897),
.Y(n_12738)
);

HB1xp67_ASAP7_75t_L g12739 ( 
.A(n_12328),
.Y(n_12739)
);

OA21x2_ASAP7_75t_L g12740 ( 
.A1(n_12366),
.A2(n_1898),
.B(n_1899),
.Y(n_12740)
);

INVx2_ASAP7_75t_L g12741 ( 
.A(n_12554),
.Y(n_12741)
);

NAND2xp5_ASAP7_75t_L g12742 ( 
.A(n_12555),
.B(n_1898),
.Y(n_12742)
);

AOI21xp5_ASAP7_75t_L g12743 ( 
.A1(n_12422),
.A2(n_1900),
.B(n_1901),
.Y(n_12743)
);

OAI21x1_ASAP7_75t_L g12744 ( 
.A1(n_12486),
.A2(n_1901),
.B(n_1902),
.Y(n_12744)
);

INVx1_ASAP7_75t_L g12745 ( 
.A(n_12370),
.Y(n_12745)
);

AND2x2_ASAP7_75t_L g12746 ( 
.A(n_12426),
.B(n_1902),
.Y(n_12746)
);

BUFx10_ASAP7_75t_L g12747 ( 
.A(n_12660),
.Y(n_12747)
);

INVx1_ASAP7_75t_SL g12748 ( 
.A(n_12604),
.Y(n_12748)
);

INVx2_ASAP7_75t_L g12749 ( 
.A(n_12424),
.Y(n_12749)
);

NAND2xp5_ASAP7_75t_L g12750 ( 
.A(n_12573),
.B(n_1903),
.Y(n_12750)
);

NAND2xp5_ASAP7_75t_L g12751 ( 
.A(n_12635),
.B(n_1903),
.Y(n_12751)
);

AOI21xp5_ASAP7_75t_SL g12752 ( 
.A1(n_12472),
.A2(n_1904),
.B(n_1905),
.Y(n_12752)
);

NAND2xp5_ASAP7_75t_L g12753 ( 
.A(n_12633),
.B(n_1904),
.Y(n_12753)
);

INVx2_ASAP7_75t_SL g12754 ( 
.A(n_12458),
.Y(n_12754)
);

NOR2xp33_ASAP7_75t_L g12755 ( 
.A(n_12405),
.B(n_12423),
.Y(n_12755)
);

OAI21xp33_ASAP7_75t_SL g12756 ( 
.A1(n_12334),
.A2(n_12401),
.B(n_12564),
.Y(n_12756)
);

INVx2_ASAP7_75t_L g12757 ( 
.A(n_12327),
.Y(n_12757)
);

OAI21x1_ASAP7_75t_L g12758 ( 
.A1(n_12376),
.A2(n_1905),
.B(n_1906),
.Y(n_12758)
);

OAI21x1_ASAP7_75t_L g12759 ( 
.A1(n_12384),
.A2(n_1906),
.B(n_1907),
.Y(n_12759)
);

INVx1_ASAP7_75t_L g12760 ( 
.A(n_12415),
.Y(n_12760)
);

OAI21x1_ASAP7_75t_L g12761 ( 
.A1(n_12336),
.A2(n_1908),
.B(n_1909),
.Y(n_12761)
);

INVx1_ASAP7_75t_L g12762 ( 
.A(n_12446),
.Y(n_12762)
);

A2O1A1Ixp33_ASAP7_75t_L g12763 ( 
.A1(n_12475),
.A2(n_1910),
.B(n_1908),
.C(n_1909),
.Y(n_12763)
);

OR2x2_ASAP7_75t_L g12764 ( 
.A(n_12431),
.B(n_1910),
.Y(n_12764)
);

NAND2xp5_ASAP7_75t_L g12765 ( 
.A(n_12606),
.B(n_1911),
.Y(n_12765)
);

AO31x2_ASAP7_75t_L g12766 ( 
.A1(n_12656),
.A2(n_1915),
.A3(n_1912),
.B(n_1913),
.Y(n_12766)
);

INVx2_ASAP7_75t_L g12767 ( 
.A(n_12478),
.Y(n_12767)
);

OAI21x1_ASAP7_75t_SL g12768 ( 
.A1(n_12465),
.A2(n_12685),
.B(n_12546),
.Y(n_12768)
);

NOR2xp33_ASAP7_75t_L g12769 ( 
.A(n_12408),
.B(n_12567),
.Y(n_12769)
);

NAND2xp5_ASAP7_75t_L g12770 ( 
.A(n_12569),
.B(n_1912),
.Y(n_12770)
);

AO21x2_ASAP7_75t_L g12771 ( 
.A1(n_12386),
.A2(n_1913),
.B(n_1916),
.Y(n_12771)
);

OAI21x1_ASAP7_75t_L g12772 ( 
.A1(n_12332),
.A2(n_1917),
.B(n_1918),
.Y(n_12772)
);

AND2x4_ASAP7_75t_L g12773 ( 
.A(n_12662),
.B(n_1917),
.Y(n_12773)
);

INVx1_ASAP7_75t_L g12774 ( 
.A(n_12448),
.Y(n_12774)
);

AND2x2_ASAP7_75t_L g12775 ( 
.A(n_12455),
.B(n_1919),
.Y(n_12775)
);

NOR2xp33_ASAP7_75t_L g12776 ( 
.A(n_12348),
.B(n_12433),
.Y(n_12776)
);

AND2x2_ASAP7_75t_L g12777 ( 
.A(n_12427),
.B(n_1919),
.Y(n_12777)
);

INVx2_ASAP7_75t_L g12778 ( 
.A(n_12614),
.Y(n_12778)
);

INVx1_ASAP7_75t_L g12779 ( 
.A(n_12461),
.Y(n_12779)
);

OAI21x1_ASAP7_75t_L g12780 ( 
.A1(n_12418),
.A2(n_1920),
.B(n_1921),
.Y(n_12780)
);

NAND2x1p5_ASAP7_75t_L g12781 ( 
.A(n_12551),
.B(n_1920),
.Y(n_12781)
);

AND2x2_ASAP7_75t_L g12782 ( 
.A(n_12439),
.B(n_1921),
.Y(n_12782)
);

AO31x2_ASAP7_75t_L g12783 ( 
.A1(n_12661),
.A2(n_12666),
.A3(n_12393),
.B(n_12411),
.Y(n_12783)
);

AOI21xp33_ASAP7_75t_SL g12784 ( 
.A1(n_12491),
.A2(n_1922),
.B(n_1923),
.Y(n_12784)
);

AOI21xp5_ASAP7_75t_L g12785 ( 
.A1(n_12390),
.A2(n_1923),
.B(n_1924),
.Y(n_12785)
);

HB1xp67_ASAP7_75t_L g12786 ( 
.A(n_12389),
.Y(n_12786)
);

AO21x1_ASAP7_75t_L g12787 ( 
.A1(n_12450),
.A2(n_1924),
.B(n_1925),
.Y(n_12787)
);

AO21x2_ASAP7_75t_L g12788 ( 
.A1(n_12640),
.A2(n_1925),
.B(n_1926),
.Y(n_12788)
);

INVx2_ASAP7_75t_L g12789 ( 
.A(n_12509),
.Y(n_12789)
);

NAND2xp5_ASAP7_75t_L g12790 ( 
.A(n_12650),
.B(n_1926),
.Y(n_12790)
);

INVx1_ASAP7_75t_L g12791 ( 
.A(n_12477),
.Y(n_12791)
);

BUFx6f_ASAP7_75t_L g12792 ( 
.A(n_12577),
.Y(n_12792)
);

OA21x2_ASAP7_75t_L g12793 ( 
.A1(n_12394),
.A2(n_1927),
.B(n_1928),
.Y(n_12793)
);

BUFx3_ASAP7_75t_L g12794 ( 
.A(n_12380),
.Y(n_12794)
);

AND2x2_ASAP7_75t_L g12795 ( 
.A(n_12445),
.B(n_1927),
.Y(n_12795)
);

AOI22xp33_ASAP7_75t_L g12796 ( 
.A1(n_12404),
.A2(n_1930),
.B1(n_1928),
.B2(n_1929),
.Y(n_12796)
);

INVx1_ASAP7_75t_L g12797 ( 
.A(n_12487),
.Y(n_12797)
);

AO31x2_ASAP7_75t_L g12798 ( 
.A1(n_12655),
.A2(n_1932),
.A3(n_1929),
.B(n_1931),
.Y(n_12798)
);

NAND2xp5_ASAP7_75t_L g12799 ( 
.A(n_12358),
.B(n_1931),
.Y(n_12799)
);

OAI21x1_ASAP7_75t_L g12800 ( 
.A1(n_12449),
.A2(n_12428),
.B(n_12601),
.Y(n_12800)
);

INVx2_ASAP7_75t_L g12801 ( 
.A(n_12337),
.Y(n_12801)
);

INVx2_ASAP7_75t_L g12802 ( 
.A(n_12482),
.Y(n_12802)
);

INVx2_ASAP7_75t_L g12803 ( 
.A(n_12582),
.Y(n_12803)
);

NAND2xp5_ASAP7_75t_L g12804 ( 
.A(n_12511),
.B(n_12540),
.Y(n_12804)
);

NOR2xp33_ASAP7_75t_SL g12805 ( 
.A(n_12499),
.B(n_12484),
.Y(n_12805)
);

INVx2_ASAP7_75t_L g12806 ( 
.A(n_12443),
.Y(n_12806)
);

AO21x2_ASAP7_75t_L g12807 ( 
.A1(n_12464),
.A2(n_1932),
.B(n_1933),
.Y(n_12807)
);

INVx1_ASAP7_75t_L g12808 ( 
.A(n_12493),
.Y(n_12808)
);

NAND2xp5_ASAP7_75t_L g12809 ( 
.A(n_12495),
.B(n_1934),
.Y(n_12809)
);

AO21x2_ASAP7_75t_L g12810 ( 
.A1(n_12563),
.A2(n_1935),
.B(n_1936),
.Y(n_12810)
);

NAND2xp5_ASAP7_75t_L g12811 ( 
.A(n_12496),
.B(n_12645),
.Y(n_12811)
);

BUFx2_ASAP7_75t_SL g12812 ( 
.A(n_12651),
.Y(n_12812)
);

AND2x2_ASAP7_75t_L g12813 ( 
.A(n_12637),
.B(n_1936),
.Y(n_12813)
);

INVx2_ASAP7_75t_L g12814 ( 
.A(n_12368),
.Y(n_12814)
);

OAI21xp5_ASAP7_75t_L g12815 ( 
.A1(n_12339),
.A2(n_1937),
.B(n_1939),
.Y(n_12815)
);

AO31x2_ASAP7_75t_L g12816 ( 
.A1(n_12603),
.A2(n_1941),
.A3(n_1939),
.B(n_1940),
.Y(n_12816)
);

INVx3_ASAP7_75t_L g12817 ( 
.A(n_12385),
.Y(n_12817)
);

BUFx2_ASAP7_75t_L g12818 ( 
.A(n_12631),
.Y(n_12818)
);

INVx1_ASAP7_75t_L g12819 ( 
.A(n_12545),
.Y(n_12819)
);

NAND2xp5_ASAP7_75t_L g12820 ( 
.A(n_12547),
.B(n_1941),
.Y(n_12820)
);

NAND2xp5_ASAP7_75t_L g12821 ( 
.A(n_12504),
.B(n_1943),
.Y(n_12821)
);

OR2x2_ASAP7_75t_L g12822 ( 
.A(n_12671),
.B(n_1943),
.Y(n_12822)
);

OAI21x1_ASAP7_75t_L g12823 ( 
.A1(n_12552),
.A2(n_1944),
.B(n_1945),
.Y(n_12823)
);

INVx2_ASAP7_75t_L g12824 ( 
.A(n_12608),
.Y(n_12824)
);

NAND2xp5_ASAP7_75t_L g12825 ( 
.A(n_12352),
.B(n_1944),
.Y(n_12825)
);

INVx2_ASAP7_75t_L g12826 ( 
.A(n_12683),
.Y(n_12826)
);

OA21x2_ASAP7_75t_L g12827 ( 
.A1(n_12316),
.A2(n_1945),
.B(n_1946),
.Y(n_12827)
);

OAI21x1_ASAP7_75t_L g12828 ( 
.A1(n_12492),
.A2(n_1947),
.B(n_1948),
.Y(n_12828)
);

INVx2_ASAP7_75t_SL g12829 ( 
.A(n_12510),
.Y(n_12829)
);

AOI22xp5_ASAP7_75t_L g12830 ( 
.A1(n_12318),
.A2(n_1950),
.B1(n_1948),
.B2(n_1949),
.Y(n_12830)
);

OAI21x1_ASAP7_75t_L g12831 ( 
.A1(n_12521),
.A2(n_1949),
.B(n_1950),
.Y(n_12831)
);

INVx2_ASAP7_75t_L g12832 ( 
.A(n_12349),
.Y(n_12832)
);

INVx1_ASAP7_75t_L g12833 ( 
.A(n_12378),
.Y(n_12833)
);

INVx1_ASAP7_75t_L g12834 ( 
.A(n_12383),
.Y(n_12834)
);

BUFx3_ASAP7_75t_L g12835 ( 
.A(n_12463),
.Y(n_12835)
);

NAND2xp5_ASAP7_75t_L g12836 ( 
.A(n_12360),
.B(n_1951),
.Y(n_12836)
);

OAI21x1_ASAP7_75t_L g12837 ( 
.A1(n_12528),
.A2(n_1951),
.B(n_1952),
.Y(n_12837)
);

AND3x4_ASAP7_75t_L g12838 ( 
.A(n_12672),
.B(n_1952),
.C(n_1954),
.Y(n_12838)
);

INVx2_ASAP7_75t_L g12839 ( 
.A(n_12621),
.Y(n_12839)
);

AND2x2_ASAP7_75t_L g12840 ( 
.A(n_12648),
.B(n_1954),
.Y(n_12840)
);

AOI21xp5_ASAP7_75t_L g12841 ( 
.A1(n_12379),
.A2(n_1955),
.B(n_1956),
.Y(n_12841)
);

INVx1_ASAP7_75t_L g12842 ( 
.A(n_12387),
.Y(n_12842)
);

NOR2xp33_ASAP7_75t_L g12843 ( 
.A(n_12558),
.B(n_1955),
.Y(n_12843)
);

AO21x2_ASAP7_75t_L g12844 ( 
.A1(n_12537),
.A2(n_1956),
.B(n_1957),
.Y(n_12844)
);

INVx1_ASAP7_75t_L g12845 ( 
.A(n_12416),
.Y(n_12845)
);

BUFx2_ASAP7_75t_L g12846 ( 
.A(n_12674),
.Y(n_12846)
);

NOR2xp33_ASAP7_75t_L g12847 ( 
.A(n_12476),
.B(n_1957),
.Y(n_12847)
);

NAND2xp5_ASAP7_75t_L g12848 ( 
.A(n_12400),
.B(n_1958),
.Y(n_12848)
);

AOI22xp33_ASAP7_75t_L g12849 ( 
.A1(n_12355),
.A2(n_1961),
.B1(n_1959),
.B2(n_1960),
.Y(n_12849)
);

OR2x6_ASAP7_75t_L g12850 ( 
.A(n_12351),
.B(n_1959),
.Y(n_12850)
);

INVx1_ASAP7_75t_L g12851 ( 
.A(n_12437),
.Y(n_12851)
);

OAI21xp5_ASAP7_75t_L g12852 ( 
.A1(n_12406),
.A2(n_1960),
.B(n_1961),
.Y(n_12852)
);

OA21x2_ASAP7_75t_L g12853 ( 
.A1(n_12553),
.A2(n_1962),
.B(n_1963),
.Y(n_12853)
);

BUFx2_ASAP7_75t_L g12854 ( 
.A(n_12619),
.Y(n_12854)
);

NAND3xp33_ASAP7_75t_L g12855 ( 
.A(n_12317),
.B(n_1962),
.C(n_1963),
.Y(n_12855)
);

INVx2_ASAP7_75t_L g12856 ( 
.A(n_12413),
.Y(n_12856)
);

AOI21xp5_ASAP7_75t_L g12857 ( 
.A1(n_12407),
.A2(n_1964),
.B(n_1965),
.Y(n_12857)
);

INVx1_ASAP7_75t_L g12858 ( 
.A(n_12452),
.Y(n_12858)
);

AOI21xp5_ASAP7_75t_L g12859 ( 
.A1(n_12399),
.A2(n_1964),
.B(n_1966),
.Y(n_12859)
);

OR2x2_ASAP7_75t_L g12860 ( 
.A(n_12556),
.B(n_1966),
.Y(n_12860)
);

O2A1O1Ixp33_ASAP7_75t_L g12861 ( 
.A1(n_12372),
.A2(n_1969),
.B(n_1967),
.C(n_1968),
.Y(n_12861)
);

OR2x2_ASAP7_75t_L g12862 ( 
.A(n_12535),
.B(n_12362),
.Y(n_12862)
);

NOR2x1_ASAP7_75t_SL g12863 ( 
.A(n_12564),
.B(n_1967),
.Y(n_12863)
);

INVx1_ASAP7_75t_L g12864 ( 
.A(n_12454),
.Y(n_12864)
);

NAND2x1p5_ASAP7_75t_L g12865 ( 
.A(n_12613),
.B(n_1968),
.Y(n_12865)
);

INVx1_ASAP7_75t_L g12866 ( 
.A(n_12481),
.Y(n_12866)
);

BUFx6f_ASAP7_75t_L g12867 ( 
.A(n_12577),
.Y(n_12867)
);

AOI22xp33_ASAP7_75t_L g12868 ( 
.A1(n_12420),
.A2(n_1972),
.B1(n_1970),
.B2(n_1971),
.Y(n_12868)
);

AO31x2_ASAP7_75t_L g12869 ( 
.A1(n_12529),
.A2(n_12409),
.A3(n_12643),
.B(n_12447),
.Y(n_12869)
);

AOI21xp5_ASAP7_75t_L g12870 ( 
.A1(n_12432),
.A2(n_12444),
.B(n_12451),
.Y(n_12870)
);

INVx1_ASAP7_75t_L g12871 ( 
.A(n_12367),
.Y(n_12871)
);

INVx2_ASAP7_75t_L g12872 ( 
.A(n_12468),
.Y(n_12872)
);

INVx1_ASAP7_75t_L g12873 ( 
.A(n_12382),
.Y(n_12873)
);

OAI21x1_ASAP7_75t_L g12874 ( 
.A1(n_12536),
.A2(n_1970),
.B(n_1971),
.Y(n_12874)
);

AO21x2_ASAP7_75t_L g12875 ( 
.A1(n_12543),
.A2(n_12474),
.B(n_12584),
.Y(n_12875)
);

INVx2_ASAP7_75t_L g12876 ( 
.A(n_12618),
.Y(n_12876)
);

INVx2_ASAP7_75t_L g12877 ( 
.A(n_12350),
.Y(n_12877)
);

AND2x2_ASAP7_75t_L g12878 ( 
.A(n_12627),
.B(n_12421),
.Y(n_12878)
);

OA21x2_ASAP7_75t_L g12879 ( 
.A1(n_12335),
.A2(n_1972),
.B(n_1973),
.Y(n_12879)
);

INVx1_ASAP7_75t_L g12880 ( 
.A(n_12392),
.Y(n_12880)
);

NAND2xp5_ASAP7_75t_L g12881 ( 
.A(n_12623),
.B(n_1973),
.Y(n_12881)
);

AO31x2_ASAP7_75t_L g12882 ( 
.A1(n_12485),
.A2(n_1976),
.A3(n_1974),
.B(n_1975),
.Y(n_12882)
);

INVx6_ASAP7_75t_L g12883 ( 
.A(n_12351),
.Y(n_12883)
);

OAI21xp5_ASAP7_75t_L g12884 ( 
.A1(n_12579),
.A2(n_1974),
.B(n_1975),
.Y(n_12884)
);

OAI21x1_ASAP7_75t_L g12885 ( 
.A1(n_12562),
.A2(n_1976),
.B(n_1977),
.Y(n_12885)
);

OR2x2_ASAP7_75t_L g12886 ( 
.A(n_12357),
.B(n_1977),
.Y(n_12886)
);

OR2x6_ASAP7_75t_L g12887 ( 
.A(n_12488),
.B(n_1978),
.Y(n_12887)
);

AOI21xp5_ASAP7_75t_L g12888 ( 
.A1(n_12412),
.A2(n_1979),
.B(n_1980),
.Y(n_12888)
);

INVx2_ASAP7_75t_L g12889 ( 
.A(n_12435),
.Y(n_12889)
);

HB1xp67_ASAP7_75t_L g12890 ( 
.A(n_12688),
.Y(n_12890)
);

INVx2_ASAP7_75t_L g12891 ( 
.A(n_12664),
.Y(n_12891)
);

OAI21x1_ASAP7_75t_L g12892 ( 
.A1(n_12565),
.A2(n_1979),
.B(n_1981),
.Y(n_12892)
);

AOI21xp5_ASAP7_75t_L g12893 ( 
.A1(n_12541),
.A2(n_1981),
.B(n_1982),
.Y(n_12893)
);

OR2x2_ASAP7_75t_L g12894 ( 
.A(n_12381),
.B(n_1982),
.Y(n_12894)
);

NAND2x1p5_ASAP7_75t_L g12895 ( 
.A(n_12522),
.B(n_1983),
.Y(n_12895)
);

AND2x4_ASAP7_75t_L g12896 ( 
.A(n_12323),
.B(n_1983),
.Y(n_12896)
);

OAI21xp5_ASAP7_75t_L g12897 ( 
.A1(n_12572),
.A2(n_1984),
.B(n_1985),
.Y(n_12897)
);

OAI21x1_ASAP7_75t_L g12898 ( 
.A1(n_12580),
.A2(n_1984),
.B(n_1986),
.Y(n_12898)
);

HB1xp67_ASAP7_75t_L g12899 ( 
.A(n_12518),
.Y(n_12899)
);

AOI21xp5_ASAP7_75t_L g12900 ( 
.A1(n_12329),
.A2(n_1986),
.B(n_1987),
.Y(n_12900)
);

INVx6_ASAP7_75t_L g12901 ( 
.A(n_12510),
.Y(n_12901)
);

INVx2_ASAP7_75t_L g12902 ( 
.A(n_12548),
.Y(n_12902)
);

AND2x2_ASAP7_75t_L g12903 ( 
.A(n_12559),
.B(n_1987),
.Y(n_12903)
);

INVx1_ASAP7_75t_L g12904 ( 
.A(n_12497),
.Y(n_12904)
);

BUFx10_ASAP7_75t_L g12905 ( 
.A(n_12488),
.Y(n_12905)
);

AO21x2_ASAP7_75t_L g12906 ( 
.A1(n_12620),
.A2(n_1988),
.B(n_1989),
.Y(n_12906)
);

NOR2xp33_ASAP7_75t_L g12907 ( 
.A(n_12520),
.B(n_1989),
.Y(n_12907)
);

AOI22xp33_ASAP7_75t_L g12908 ( 
.A1(n_12403),
.A2(n_1992),
.B1(n_1990),
.B2(n_1991),
.Y(n_12908)
);

AND2x4_ASAP7_75t_SL g12909 ( 
.A(n_12599),
.B(n_1990),
.Y(n_12909)
);

OAI21xp33_ASAP7_75t_L g12910 ( 
.A1(n_12419),
.A2(n_1992),
.B(n_1993),
.Y(n_12910)
);

NAND2xp5_ASAP7_75t_L g12911 ( 
.A(n_12657),
.B(n_1993),
.Y(n_12911)
);

AND2x4_ASAP7_75t_L g12912 ( 
.A(n_12616),
.B(n_1994),
.Y(n_12912)
);

HB1xp67_ASAP7_75t_L g12913 ( 
.A(n_12359),
.Y(n_12913)
);

OAI21xp5_ASAP7_75t_L g12914 ( 
.A1(n_12531),
.A2(n_1994),
.B(n_1995),
.Y(n_12914)
);

OR2x6_ASAP7_75t_L g12915 ( 
.A(n_12599),
.B(n_1995),
.Y(n_12915)
);

NAND2xp5_ASAP7_75t_L g12916 ( 
.A(n_12532),
.B(n_1997),
.Y(n_12916)
);

INVx1_ASAP7_75t_L g12917 ( 
.A(n_12497),
.Y(n_12917)
);

INVx2_ASAP7_75t_SL g12918 ( 
.A(n_12544),
.Y(n_12918)
);

INVx1_ASAP7_75t_L g12919 ( 
.A(n_12524),
.Y(n_12919)
);

OAI21xp5_ASAP7_75t_L g12920 ( 
.A1(n_12391),
.A2(n_1998),
.B(n_2000),
.Y(n_12920)
);

INVx3_ASAP7_75t_L g12921 ( 
.A(n_12542),
.Y(n_12921)
);

INVx2_ASAP7_75t_L g12922 ( 
.A(n_12483),
.Y(n_12922)
);

OAI21x1_ASAP7_75t_L g12923 ( 
.A1(n_12658),
.A2(n_12326),
.B(n_12333),
.Y(n_12923)
);

INVx2_ASAP7_75t_SL g12924 ( 
.A(n_12595),
.Y(n_12924)
);

BUFx8_ASAP7_75t_L g12925 ( 
.A(n_12597),
.Y(n_12925)
);

INVx2_ASAP7_75t_L g12926 ( 
.A(n_12500),
.Y(n_12926)
);

INVx1_ASAP7_75t_L g12927 ( 
.A(n_12524),
.Y(n_12927)
);

AO31x2_ASAP7_75t_L g12928 ( 
.A1(n_12441),
.A2(n_2001),
.A3(n_1998),
.B(n_2000),
.Y(n_12928)
);

BUFx12f_ASAP7_75t_L g12929 ( 
.A(n_12530),
.Y(n_12929)
);

OAI21x1_ASAP7_75t_L g12930 ( 
.A1(n_12677),
.A2(n_2001),
.B(n_2002),
.Y(n_12930)
);

OA21x2_ASAP7_75t_L g12931 ( 
.A1(n_12576),
.A2(n_12679),
.B(n_12646),
.Y(n_12931)
);

OA21x2_ASAP7_75t_L g12932 ( 
.A1(n_12638),
.A2(n_2003),
.B(n_2004),
.Y(n_12932)
);

AOI21xp5_ASAP7_75t_L g12933 ( 
.A1(n_12434),
.A2(n_2003),
.B(n_2004),
.Y(n_12933)
);

AOI21xp5_ASAP7_75t_L g12934 ( 
.A1(n_12659),
.A2(n_2005),
.B(n_2006),
.Y(n_12934)
);

INVx1_ASAP7_75t_L g12935 ( 
.A(n_12467),
.Y(n_12935)
);

INVx1_ASAP7_75t_L g12936 ( 
.A(n_12639),
.Y(n_12936)
);

AND2x2_ASAP7_75t_L g12937 ( 
.A(n_12684),
.B(n_2005),
.Y(n_12937)
);

AO21x2_ASAP7_75t_L g12938 ( 
.A1(n_12665),
.A2(n_2006),
.B(n_2007),
.Y(n_12938)
);

NAND2xp5_ASAP7_75t_L g12939 ( 
.A(n_12539),
.B(n_12607),
.Y(n_12939)
);

INVx1_ASAP7_75t_L g12940 ( 
.A(n_12459),
.Y(n_12940)
);

OA21x2_ASAP7_75t_L g12941 ( 
.A1(n_12605),
.A2(n_2007),
.B(n_2008),
.Y(n_12941)
);

INVx2_ASAP7_75t_L g12942 ( 
.A(n_12592),
.Y(n_12942)
);

AOI21xp5_ASAP7_75t_L g12943 ( 
.A1(n_12473),
.A2(n_2008),
.B(n_2009),
.Y(n_12943)
);

BUFx10_ASAP7_75t_L g12944 ( 
.A(n_12457),
.Y(n_12944)
);

NAND3xp33_ASAP7_75t_L g12945 ( 
.A(n_12417),
.B(n_2009),
.C(n_2010),
.Y(n_12945)
);

OA21x2_ASAP7_75t_L g12946 ( 
.A1(n_12574),
.A2(n_2010),
.B(n_2011),
.Y(n_12946)
);

OR2x2_ASAP7_75t_L g12947 ( 
.A(n_12381),
.B(n_2011),
.Y(n_12947)
);

AOI21xp5_ASAP7_75t_L g12948 ( 
.A1(n_12634),
.A2(n_2012),
.B(n_2013),
.Y(n_12948)
);

AOI21xp5_ASAP7_75t_L g12949 ( 
.A1(n_12506),
.A2(n_2013),
.B(n_2014),
.Y(n_12949)
);

INVx1_ASAP7_75t_SL g12950 ( 
.A(n_12632),
.Y(n_12950)
);

AOI222xp33_ASAP7_75t_SL g12951 ( 
.A1(n_12353),
.A2(n_12501),
.B1(n_12321),
.B2(n_12587),
.C1(n_12602),
.C2(n_12611),
.Y(n_12951)
);

OA21x2_ASAP7_75t_L g12952 ( 
.A1(n_12649),
.A2(n_2014),
.B(n_2015),
.Y(n_12952)
);

NAND2xp5_ASAP7_75t_L g12953 ( 
.A(n_12610),
.B(n_2015),
.Y(n_12953)
);

NAND2xp5_ASAP7_75t_L g12954 ( 
.A(n_12686),
.B(n_2016),
.Y(n_12954)
);

INVx1_ASAP7_75t_L g12955 ( 
.A(n_12460),
.Y(n_12955)
);

NAND2xp5_ASAP7_75t_L g12956 ( 
.A(n_12682),
.B(n_2016),
.Y(n_12956)
);

AOI21xp5_ASAP7_75t_L g12957 ( 
.A1(n_12549),
.A2(n_2017),
.B(n_2018),
.Y(n_12957)
);

INVx1_ASAP7_75t_L g12958 ( 
.A(n_12517),
.Y(n_12958)
);

AOI22xp33_ASAP7_75t_L g12959 ( 
.A1(n_12398),
.A2(n_2020),
.B1(n_2018),
.B2(n_2019),
.Y(n_12959)
);

INVx2_ASAP7_75t_L g12960 ( 
.A(n_12652),
.Y(n_12960)
);

INVx2_ASAP7_75t_L g12961 ( 
.A(n_12489),
.Y(n_12961)
);

INVx1_ASAP7_75t_L g12962 ( 
.A(n_12628),
.Y(n_12962)
);

BUFx2_ASAP7_75t_L g12963 ( 
.A(n_12321),
.Y(n_12963)
);

INVx2_ASAP7_75t_L g12964 ( 
.A(n_12503),
.Y(n_12964)
);

AO21x2_ASAP7_75t_L g12965 ( 
.A1(n_12494),
.A2(n_2019),
.B(n_2020),
.Y(n_12965)
);

OA21x2_ASAP7_75t_L g12966 ( 
.A1(n_12591),
.A2(n_2021),
.B(n_2022),
.Y(n_12966)
);

INVx3_ASAP7_75t_L g12967 ( 
.A(n_12680),
.Y(n_12967)
);

AO31x2_ASAP7_75t_L g12968 ( 
.A1(n_12375),
.A2(n_2024),
.A3(n_2022),
.B(n_2023),
.Y(n_12968)
);

OAI21xp33_ASAP7_75t_L g12969 ( 
.A1(n_12341),
.A2(n_2024),
.B(n_2025),
.Y(n_12969)
);

OR2x2_ASAP7_75t_L g12970 ( 
.A(n_12373),
.B(n_12681),
.Y(n_12970)
);

OA21x2_ASAP7_75t_L g12971 ( 
.A1(n_12470),
.A2(n_2025),
.B(n_2026),
.Y(n_12971)
);

NAND2xp5_ASAP7_75t_L g12972 ( 
.A(n_12480),
.B(n_2026),
.Y(n_12972)
);

NAND2xp5_ASAP7_75t_L g12973 ( 
.A(n_12490),
.B(n_2027),
.Y(n_12973)
);

OAI21x1_ASAP7_75t_L g12974 ( 
.A1(n_12560),
.A2(n_2027),
.B(n_2028),
.Y(n_12974)
);

OA21x2_ASAP7_75t_L g12975 ( 
.A1(n_12625),
.A2(n_2028),
.B(n_2029),
.Y(n_12975)
);

INVx1_ASAP7_75t_L g12976 ( 
.A(n_12507),
.Y(n_12976)
);

NAND2xp5_ASAP7_75t_L g12977 ( 
.A(n_12681),
.B(n_2029),
.Y(n_12977)
);

CKINVDCx20_ASAP7_75t_R g12978 ( 
.A(n_12663),
.Y(n_12978)
);

INVx1_ASAP7_75t_L g12979 ( 
.A(n_12513),
.Y(n_12979)
);

AND2x4_ASAP7_75t_L g12980 ( 
.A(n_12525),
.B(n_12653),
.Y(n_12980)
);

INVx1_ASAP7_75t_SL g12981 ( 
.A(n_12629),
.Y(n_12981)
);

OAI21x1_ASAP7_75t_L g12982 ( 
.A1(n_12363),
.A2(n_2030),
.B(n_2031),
.Y(n_12982)
);

A2O1A1Ixp33_ASAP7_75t_L g12983 ( 
.A1(n_12456),
.A2(n_2032),
.B(n_2030),
.C(n_2031),
.Y(n_12983)
);

OR2x2_ASAP7_75t_L g12984 ( 
.A(n_12373),
.B(n_2032),
.Y(n_12984)
);

NAND2xp5_ASAP7_75t_L g12985 ( 
.A(n_12586),
.B(n_2033),
.Y(n_12985)
);

INVx1_ASAP7_75t_L g12986 ( 
.A(n_12654),
.Y(n_12986)
);

INVx1_ASAP7_75t_L g12987 ( 
.A(n_12617),
.Y(n_12987)
);

INVx1_ASAP7_75t_L g12988 ( 
.A(n_12581),
.Y(n_12988)
);

A2O1A1Ixp33_ASAP7_75t_L g12989 ( 
.A1(n_12550),
.A2(n_2036),
.B(n_2034),
.C(n_2035),
.Y(n_12989)
);

INVx3_ASAP7_75t_L g12990 ( 
.A(n_12469),
.Y(n_12990)
);

BUFx3_ASAP7_75t_L g12991 ( 
.A(n_12515),
.Y(n_12991)
);

AOI21xp33_ASAP7_75t_SL g12992 ( 
.A1(n_12594),
.A2(n_2034),
.B(n_2036),
.Y(n_12992)
);

AOI21xp5_ASAP7_75t_L g12993 ( 
.A1(n_12578),
.A2(n_2037),
.B(n_2038),
.Y(n_12993)
);

NAND2xp5_ASAP7_75t_L g12994 ( 
.A(n_12585),
.B(n_2037),
.Y(n_12994)
);

AND2x2_ASAP7_75t_L g12995 ( 
.A(n_12653),
.B(n_2038),
.Y(n_12995)
);

BUFx12f_ASAP7_75t_L g12996 ( 
.A(n_12644),
.Y(n_12996)
);

AOI21x1_ASAP7_75t_L g12997 ( 
.A1(n_12583),
.A2(n_2039),
.B(n_2040),
.Y(n_12997)
);

NAND2x1p5_ASAP7_75t_L g12998 ( 
.A(n_12678),
.B(n_2039),
.Y(n_12998)
);

AOI21xp5_ASAP7_75t_L g12999 ( 
.A1(n_12429),
.A2(n_12519),
.B(n_12641),
.Y(n_12999)
);

OAI21x1_ASAP7_75t_L g13000 ( 
.A1(n_12596),
.A2(n_2040),
.B(n_2041),
.Y(n_13000)
);

AOI21xp5_ASAP7_75t_L g13001 ( 
.A1(n_12647),
.A2(n_2041),
.B(n_2042),
.Y(n_13001)
);

AND2x2_ASAP7_75t_L g13002 ( 
.A(n_12644),
.B(n_2042),
.Y(n_13002)
);

OA21x2_ASAP7_75t_L g13003 ( 
.A1(n_12626),
.A2(n_2043),
.B(n_2044),
.Y(n_13003)
);

OR2x2_ASAP7_75t_L g13004 ( 
.A(n_12364),
.B(n_2043),
.Y(n_13004)
);

OAI21x1_ASAP7_75t_L g13005 ( 
.A1(n_12609),
.A2(n_2045),
.B(n_2046),
.Y(n_13005)
);

AOI21x1_ASAP7_75t_L g13006 ( 
.A1(n_12636),
.A2(n_2045),
.B(n_2046),
.Y(n_13006)
);

INVx1_ASAP7_75t_L g13007 ( 
.A(n_12669),
.Y(n_13007)
);

NAND2xp5_ASAP7_75t_L g13008 ( 
.A(n_12585),
.B(n_2047),
.Y(n_13008)
);

NAND2xp5_ASAP7_75t_L g13009 ( 
.A(n_12364),
.B(n_2047),
.Y(n_13009)
);

OAI21x1_ASAP7_75t_L g13010 ( 
.A1(n_12612),
.A2(n_12670),
.B(n_12589),
.Y(n_13010)
);

AO21x2_ASAP7_75t_L g13011 ( 
.A1(n_12566),
.A2(n_2048),
.B(n_2049),
.Y(n_13011)
);

OAI21x1_ASAP7_75t_SL g13012 ( 
.A1(n_12600),
.A2(n_2048),
.B(n_2049),
.Y(n_13012)
);

AND2x2_ASAP7_75t_L g13013 ( 
.A(n_12508),
.B(n_2050),
.Y(n_13013)
);

BUFx6f_ASAP7_75t_L g13014 ( 
.A(n_12570),
.Y(n_13014)
);

NAND2xp5_ASAP7_75t_L g13015 ( 
.A(n_12571),
.B(n_2050),
.Y(n_13015)
);

NAND2x1p5_ASAP7_75t_L g13016 ( 
.A(n_12673),
.B(n_12340),
.Y(n_13016)
);

OR2x2_ASAP7_75t_L g13017 ( 
.A(n_12471),
.B(n_2051),
.Y(n_13017)
);

AO21x1_ASAP7_75t_L g13018 ( 
.A1(n_12676),
.A2(n_2052),
.B(n_2053),
.Y(n_13018)
);

AOI21xp5_ASAP7_75t_L g13019 ( 
.A1(n_12557),
.A2(n_2052),
.B(n_2054),
.Y(n_13019)
);

INVx2_ASAP7_75t_SL g13020 ( 
.A(n_12590),
.Y(n_13020)
);

INVx2_ASAP7_75t_L g13021 ( 
.A(n_12526),
.Y(n_13021)
);

INVx1_ASAP7_75t_L g13022 ( 
.A(n_12538),
.Y(n_13022)
);

HB1xp67_ASAP7_75t_L g13023 ( 
.A(n_12668),
.Y(n_13023)
);

INVx3_ASAP7_75t_L g13024 ( 
.A(n_12598),
.Y(n_13024)
);

AOI21xp5_ASAP7_75t_L g13025 ( 
.A1(n_12630),
.A2(n_2054),
.B(n_2055),
.Y(n_13025)
);

NOR2xp33_ASAP7_75t_L g13026 ( 
.A(n_12687),
.B(n_2055),
.Y(n_13026)
);

OA21x2_ASAP7_75t_L g13027 ( 
.A1(n_12624),
.A2(n_2056),
.B(n_2057),
.Y(n_13027)
);

INVx1_ASAP7_75t_L g13028 ( 
.A(n_12667),
.Y(n_13028)
);

AO21x2_ASAP7_75t_L g13029 ( 
.A1(n_12568),
.A2(n_2056),
.B(n_2057),
.Y(n_13029)
);

INVxp33_ASAP7_75t_L g13030 ( 
.A(n_12622),
.Y(n_13030)
);

INVx2_ASAP7_75t_SL g13031 ( 
.A(n_12458),
.Y(n_13031)
);

NAND2xp5_ASAP7_75t_L g13032 ( 
.A(n_12527),
.B(n_2058),
.Y(n_13032)
);

CKINVDCx8_ASAP7_75t_R g13033 ( 
.A(n_12523),
.Y(n_13033)
);

OAI21x1_ASAP7_75t_SL g13034 ( 
.A1(n_12324),
.A2(n_2058),
.B(n_2059),
.Y(n_13034)
);

AND2x2_ASAP7_75t_L g13035 ( 
.A(n_12344),
.B(n_2060),
.Y(n_13035)
);

AOI21xp33_ASAP7_75t_SL g13036 ( 
.A1(n_12533),
.A2(n_2060),
.B(n_2061),
.Y(n_13036)
);

XNOR2xp5_ASAP7_75t_L g13037 ( 
.A(n_12425),
.B(n_2061),
.Y(n_13037)
);

AND2x2_ASAP7_75t_L g13038 ( 
.A(n_12344),
.B(n_2062),
.Y(n_13038)
);

INVx2_ASAP7_75t_SL g13039 ( 
.A(n_12458),
.Y(n_13039)
);

INVx6_ASAP7_75t_L g13040 ( 
.A(n_12516),
.Y(n_13040)
);

INVx2_ASAP7_75t_SL g13041 ( 
.A(n_13040),
.Y(n_13041)
);

HB1xp67_ASAP7_75t_L g13042 ( 
.A(n_12879),
.Y(n_13042)
);

INVx2_ASAP7_75t_L g13043 ( 
.A(n_12835),
.Y(n_13043)
);

OAI21xp33_ASAP7_75t_SL g13044 ( 
.A1(n_12704),
.A2(n_2062),
.B(n_2063),
.Y(n_13044)
);

BUFx2_ASAP7_75t_L g13045 ( 
.A(n_12818),
.Y(n_13045)
);

INVx2_ASAP7_75t_L g13046 ( 
.A(n_12854),
.Y(n_13046)
);

INVx1_ASAP7_75t_L g13047 ( 
.A(n_12766),
.Y(n_13047)
);

INVx3_ASAP7_75t_L g13048 ( 
.A(n_13033),
.Y(n_13048)
);

INVx3_ASAP7_75t_L g13049 ( 
.A(n_12929),
.Y(n_13049)
);

AND2x2_ASAP7_75t_L g13050 ( 
.A(n_12878),
.B(n_2063),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_12766),
.Y(n_13051)
);

INVx1_ASAP7_75t_L g13052 ( 
.A(n_12798),
.Y(n_13052)
);

INVx2_ASAP7_75t_L g13053 ( 
.A(n_12794),
.Y(n_13053)
);

INVx1_ASAP7_75t_L g13054 ( 
.A(n_12798),
.Y(n_13054)
);

INVx1_ASAP7_75t_L g13055 ( 
.A(n_12710),
.Y(n_13055)
);

INVx1_ASAP7_75t_L g13056 ( 
.A(n_12706),
.Y(n_13056)
);

OAI21x1_ASAP7_75t_L g13057 ( 
.A1(n_12800),
.A2(n_2064),
.B(n_2065),
.Y(n_13057)
);

INVx1_ASAP7_75t_L g13058 ( 
.A(n_12708),
.Y(n_13058)
);

AND2x2_ASAP7_75t_L g13059 ( 
.A(n_12728),
.B(n_2064),
.Y(n_13059)
);

INVx2_ASAP7_75t_L g13060 ( 
.A(n_12730),
.Y(n_13060)
);

INVx1_ASAP7_75t_L g13061 ( 
.A(n_12714),
.Y(n_13061)
);

OAI21x1_ASAP7_75t_L g13062 ( 
.A1(n_12741),
.A2(n_2065),
.B(n_2066),
.Y(n_13062)
);

AND2x4_ASAP7_75t_L g13063 ( 
.A(n_12754),
.B(n_2066),
.Y(n_13063)
);

INVx2_ASAP7_75t_L g13064 ( 
.A(n_12730),
.Y(n_13064)
);

AO21x2_ASAP7_75t_L g13065 ( 
.A1(n_12727),
.A2(n_12799),
.B(n_12825),
.Y(n_13065)
);

INVx2_ASAP7_75t_L g13066 ( 
.A(n_13010),
.Y(n_13066)
);

INVx2_ASAP7_75t_L g13067 ( 
.A(n_12707),
.Y(n_13067)
);

OAI21x1_ASAP7_75t_L g13068 ( 
.A1(n_12803),
.A2(n_2067),
.B(n_2068),
.Y(n_13068)
);

HB1xp67_ASAP7_75t_L g13069 ( 
.A(n_12866),
.Y(n_13069)
);

BUFx2_ASAP7_75t_L g13070 ( 
.A(n_12846),
.Y(n_13070)
);

INVx1_ASAP7_75t_SL g13071 ( 
.A(n_12812),
.Y(n_13071)
);

BUFx2_ASAP7_75t_L g13072 ( 
.A(n_13031),
.Y(n_13072)
);

INVx2_ASAP7_75t_L g13073 ( 
.A(n_12982),
.Y(n_13073)
);

AND2x2_ASAP7_75t_L g13074 ( 
.A(n_12715),
.B(n_2067),
.Y(n_13074)
);

INVx1_ASAP7_75t_L g13075 ( 
.A(n_12719),
.Y(n_13075)
);

AOI22xp33_ASAP7_75t_L g13076 ( 
.A1(n_12963),
.A2(n_2070),
.B1(n_2068),
.B2(n_2069),
.Y(n_13076)
);

INVx1_ASAP7_75t_L g13077 ( 
.A(n_12745),
.Y(n_13077)
);

OAI22xp5_ASAP7_75t_L g13078 ( 
.A1(n_12849),
.A2(n_2072),
.B1(n_2069),
.B2(n_2071),
.Y(n_13078)
);

INVx1_ASAP7_75t_L g13079 ( 
.A(n_12760),
.Y(n_13079)
);

INVx1_ASAP7_75t_L g13080 ( 
.A(n_12762),
.Y(n_13080)
);

INVx1_ASAP7_75t_L g13081 ( 
.A(n_12774),
.Y(n_13081)
);

AOI21x1_ASAP7_75t_L g13082 ( 
.A1(n_12890),
.A2(n_2072),
.B(n_2073),
.Y(n_13082)
);

INVx1_ASAP7_75t_L g13083 ( 
.A(n_12779),
.Y(n_13083)
);

INVx1_ASAP7_75t_L g13084 ( 
.A(n_12791),
.Y(n_13084)
);

INVx2_ASAP7_75t_L g13085 ( 
.A(n_12817),
.Y(n_13085)
);

CKINVDCx11_ASAP7_75t_R g13086 ( 
.A(n_12695),
.Y(n_13086)
);

INVx1_ASAP7_75t_L g13087 ( 
.A(n_12797),
.Y(n_13087)
);

INVx3_ASAP7_75t_L g13088 ( 
.A(n_12883),
.Y(n_13088)
);

INVx2_ASAP7_75t_L g13089 ( 
.A(n_12905),
.Y(n_13089)
);

INVx1_ASAP7_75t_L g13090 ( 
.A(n_12808),
.Y(n_13090)
);

INVx2_ASAP7_75t_L g13091 ( 
.A(n_12740),
.Y(n_13091)
);

INVx1_ASAP7_75t_L g13092 ( 
.A(n_12819),
.Y(n_13092)
);

INVx2_ASAP7_75t_L g13093 ( 
.A(n_13014),
.Y(n_13093)
);

HB1xp67_ASAP7_75t_L g13094 ( 
.A(n_12729),
.Y(n_13094)
);

AND2x2_ASAP7_75t_L g13095 ( 
.A(n_12921),
.B(n_2074),
.Y(n_13095)
);

INVx3_ASAP7_75t_L g13096 ( 
.A(n_12792),
.Y(n_13096)
);

HB1xp67_ASAP7_75t_L g13097 ( 
.A(n_12691),
.Y(n_13097)
);

INVx4_ASAP7_75t_L g13098 ( 
.A(n_12734),
.Y(n_13098)
);

OA21x2_ASAP7_75t_L g13099 ( 
.A1(n_12870),
.A2(n_2074),
.B(n_2076),
.Y(n_13099)
);

AND2x2_ASAP7_75t_L g13100 ( 
.A(n_12736),
.B(n_2076),
.Y(n_13100)
);

INVx1_ASAP7_75t_SL g13101 ( 
.A(n_12703),
.Y(n_13101)
);

INVx2_ASAP7_75t_L g13102 ( 
.A(n_13014),
.Y(n_13102)
);

INVx2_ASAP7_75t_SL g13103 ( 
.A(n_12901),
.Y(n_13103)
);

INVx1_ASAP7_75t_L g13104 ( 
.A(n_12904),
.Y(n_13104)
);

AND2x2_ASAP7_75t_L g13105 ( 
.A(n_12889),
.B(n_2077),
.Y(n_13105)
);

INVx2_ASAP7_75t_L g13106 ( 
.A(n_12886),
.Y(n_13106)
);

BUFx3_ASAP7_75t_L g13107 ( 
.A(n_12978),
.Y(n_13107)
);

INVx1_ASAP7_75t_L g13108 ( 
.A(n_12917),
.Y(n_13108)
);

INVx3_ASAP7_75t_L g13109 ( 
.A(n_12792),
.Y(n_13109)
);

INVx4_ASAP7_75t_L g13110 ( 
.A(n_12867),
.Y(n_13110)
);

INVx3_ASAP7_75t_L g13111 ( 
.A(n_12867),
.Y(n_13111)
);

INVx1_ASAP7_75t_L g13112 ( 
.A(n_12919),
.Y(n_13112)
);

INVx2_ASAP7_75t_L g13113 ( 
.A(n_12718),
.Y(n_13113)
);

INVx1_ASAP7_75t_L g13114 ( 
.A(n_12927),
.Y(n_13114)
);

AND2x2_ASAP7_75t_L g13115 ( 
.A(n_12967),
.B(n_2078),
.Y(n_13115)
);

AO21x2_ASAP7_75t_L g13116 ( 
.A1(n_12742),
.A2(n_2078),
.B(n_2079),
.Y(n_13116)
);

CKINVDCx6p67_ASAP7_75t_R g13117 ( 
.A(n_12721),
.Y(n_13117)
);

AO21x2_ASAP7_75t_L g13118 ( 
.A1(n_12750),
.A2(n_2079),
.B(n_2080),
.Y(n_13118)
);

INVx1_ASAP7_75t_L g13119 ( 
.A(n_12788),
.Y(n_13119)
);

AO21x2_ASAP7_75t_L g13120 ( 
.A1(n_12751),
.A2(n_2080),
.B(n_2081),
.Y(n_13120)
);

INVx1_ASAP7_75t_L g13121 ( 
.A(n_12962),
.Y(n_13121)
);

BUFx2_ASAP7_75t_SL g13122 ( 
.A(n_12748),
.Y(n_13122)
);

NAND2xp5_ASAP7_75t_L g13123 ( 
.A(n_12894),
.B(n_2081),
.Y(n_13123)
);

INVx1_ASAP7_75t_L g13124 ( 
.A(n_12986),
.Y(n_13124)
);

INVx1_ASAP7_75t_L g13125 ( 
.A(n_12936),
.Y(n_13125)
);

OAI21x1_ASAP7_75t_L g13126 ( 
.A1(n_12811),
.A2(n_2082),
.B(n_2083),
.Y(n_13126)
);

BUFx2_ASAP7_75t_L g13127 ( 
.A(n_13039),
.Y(n_13127)
);

OAI21xp5_ASAP7_75t_L g13128 ( 
.A1(n_12900),
.A2(n_2082),
.B(n_2083),
.Y(n_13128)
);

CKINVDCx20_ASAP7_75t_R g13129 ( 
.A(n_12925),
.Y(n_13129)
);

BUFx10_ASAP7_75t_L g13130 ( 
.A(n_12843),
.Y(n_13130)
);

INVx1_ASAP7_75t_L g13131 ( 
.A(n_12696),
.Y(n_13131)
);

OAI21x1_ASAP7_75t_L g13132 ( 
.A1(n_12757),
.A2(n_2084),
.B(n_2086),
.Y(n_13132)
);

AO21x2_ASAP7_75t_L g13133 ( 
.A1(n_12753),
.A2(n_2084),
.B(n_2086),
.Y(n_13133)
);

OAI21x1_ASAP7_75t_L g13134 ( 
.A1(n_12694),
.A2(n_2087),
.B(n_2088),
.Y(n_13134)
);

INVx1_ASAP7_75t_L g13135 ( 
.A(n_12697),
.Y(n_13135)
);

AND2x4_ASAP7_75t_L g13136 ( 
.A(n_12991),
.B(n_2088),
.Y(n_13136)
);

INVx2_ASAP7_75t_L g13137 ( 
.A(n_12827),
.Y(n_13137)
);

AND2x2_ASAP7_75t_L g13138 ( 
.A(n_12990),
.B(n_2089),
.Y(n_13138)
);

OAI21x1_ASAP7_75t_L g13139 ( 
.A1(n_12814),
.A2(n_2089),
.B(n_2090),
.Y(n_13139)
);

CKINVDCx5p33_ASAP7_75t_R g13140 ( 
.A(n_12701),
.Y(n_13140)
);

INVx1_ASAP7_75t_L g13141 ( 
.A(n_12700),
.Y(n_13141)
);

BUFx2_ASAP7_75t_L g13142 ( 
.A(n_12756),
.Y(n_13142)
);

AND2x2_ASAP7_75t_L g13143 ( 
.A(n_12693),
.B(n_12769),
.Y(n_13143)
);

INVx1_ASAP7_75t_L g13144 ( 
.A(n_12705),
.Y(n_13144)
);

INVx2_ASAP7_75t_L g13145 ( 
.A(n_12966),
.Y(n_13145)
);

INVx1_ASAP7_75t_L g13146 ( 
.A(n_12783),
.Y(n_13146)
);

INVx3_ASAP7_75t_L g13147 ( 
.A(n_12996),
.Y(n_13147)
);

INVx2_ASAP7_75t_SL g13148 ( 
.A(n_12915),
.Y(n_13148)
);

INVx1_ASAP7_75t_L g13149 ( 
.A(n_12783),
.Y(n_13149)
);

INVx1_ASAP7_75t_L g13150 ( 
.A(n_12947),
.Y(n_13150)
);

INVx3_ASAP7_75t_L g13151 ( 
.A(n_12915),
.Y(n_13151)
);

OA21x2_ASAP7_75t_L g13152 ( 
.A1(n_12935),
.A2(n_2090),
.B(n_2091),
.Y(n_13152)
);

INVx2_ASAP7_75t_L g13153 ( 
.A(n_12690),
.Y(n_13153)
);

BUFx3_ASAP7_75t_L g13154 ( 
.A(n_12850),
.Y(n_13154)
);

AO21x2_ASAP7_75t_L g13155 ( 
.A1(n_12765),
.A2(n_2092),
.B(n_2093),
.Y(n_13155)
);

INVx2_ASAP7_75t_L g13156 ( 
.A(n_12971),
.Y(n_13156)
);

INVx1_ASAP7_75t_L g13157 ( 
.A(n_12899),
.Y(n_13157)
);

INVx2_ASAP7_75t_L g13158 ( 
.A(n_13004),
.Y(n_13158)
);

AOI21x1_ASAP7_75t_L g13159 ( 
.A1(n_12848),
.A2(n_12836),
.B(n_12775),
.Y(n_13159)
);

INVx1_ASAP7_75t_L g13160 ( 
.A(n_12994),
.Y(n_13160)
);

BUFx3_ASAP7_75t_L g13161 ( 
.A(n_12850),
.Y(n_13161)
);

HB1xp67_ASAP7_75t_L g13162 ( 
.A(n_12739),
.Y(n_13162)
);

INVx3_ASAP7_75t_L g13163 ( 
.A(n_12699),
.Y(n_13163)
);

BUFx2_ASAP7_75t_L g13164 ( 
.A(n_12931),
.Y(n_13164)
);

INVx1_ASAP7_75t_L g13165 ( 
.A(n_13008),
.Y(n_13165)
);

BUFx3_ASAP7_75t_L g13166 ( 
.A(n_12909),
.Y(n_13166)
);

INVx2_ASAP7_75t_L g13167 ( 
.A(n_12946),
.Y(n_13167)
);

INVxp67_ASAP7_75t_SL g13168 ( 
.A(n_12787),
.Y(n_13168)
);

INVx2_ASAP7_75t_L g13169 ( 
.A(n_12802),
.Y(n_13169)
);

INVxp67_ASAP7_75t_L g13170 ( 
.A(n_12755),
.Y(n_13170)
);

INVx1_ASAP7_75t_L g13171 ( 
.A(n_13007),
.Y(n_13171)
);

INVx1_ASAP7_75t_L g13172 ( 
.A(n_12717),
.Y(n_13172)
);

INVx2_ASAP7_75t_L g13173 ( 
.A(n_12767),
.Y(n_13173)
);

INVx1_ASAP7_75t_L g13174 ( 
.A(n_12790),
.Y(n_13174)
);

AO21x2_ASAP7_75t_L g13175 ( 
.A1(n_13009),
.A2(n_2092),
.B(n_2093),
.Y(n_13175)
);

INVx1_ASAP7_75t_L g13176 ( 
.A(n_12958),
.Y(n_13176)
);

INVxp33_ASAP7_75t_L g13177 ( 
.A(n_13037),
.Y(n_13177)
);

NAND2xp5_ASAP7_75t_L g13178 ( 
.A(n_12793),
.B(n_2094),
.Y(n_13178)
);

AOI21x1_ASAP7_75t_L g13179 ( 
.A1(n_12939),
.A2(n_2095),
.B(n_2096),
.Y(n_13179)
);

HB1xp67_ASAP7_75t_L g13180 ( 
.A(n_12942),
.Y(n_13180)
);

INVx1_ASAP7_75t_L g13181 ( 
.A(n_12940),
.Y(n_13181)
);

HB1xp67_ASAP7_75t_L g13182 ( 
.A(n_12872),
.Y(n_13182)
);

INVx1_ASAP7_75t_L g13183 ( 
.A(n_12955),
.Y(n_13183)
);

NOR2xp33_ASAP7_75t_L g13184 ( 
.A(n_12805),
.B(n_2095),
.Y(n_13184)
);

AND2x2_ASAP7_75t_L g13185 ( 
.A(n_12732),
.B(n_2097),
.Y(n_13185)
);

INVx1_ASAP7_75t_L g13186 ( 
.A(n_12976),
.Y(n_13186)
);

INVx2_ASAP7_75t_L g13187 ( 
.A(n_12950),
.Y(n_13187)
);

INVx1_ASAP7_75t_L g13188 ( 
.A(n_12954),
.Y(n_13188)
);

BUFx2_ASAP7_75t_L g13189 ( 
.A(n_12932),
.Y(n_13189)
);

INVx2_ASAP7_75t_L g13190 ( 
.A(n_12922),
.Y(n_13190)
);

NAND2xp5_ASAP7_75t_L g13191 ( 
.A(n_12777),
.B(n_2097),
.Y(n_13191)
);

HB1xp67_ASAP7_75t_L g13192 ( 
.A(n_12876),
.Y(n_13192)
);

OAI21x1_ASAP7_75t_L g13193 ( 
.A1(n_12801),
.A2(n_2098),
.B(n_2099),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_12956),
.Y(n_13194)
);

INVx1_ASAP7_75t_L g13195 ( 
.A(n_12770),
.Y(n_13195)
);

INVx1_ASAP7_75t_L g13196 ( 
.A(n_12804),
.Y(n_13196)
);

AOI22xp33_ASAP7_75t_L g13197 ( 
.A1(n_13023),
.A2(n_2101),
.B1(n_2099),
.B2(n_2100),
.Y(n_13197)
);

INVx2_ASAP7_75t_L g13198 ( 
.A(n_12926),
.Y(n_13198)
);

AO21x2_ASAP7_75t_L g13199 ( 
.A1(n_12722),
.A2(n_2100),
.B(n_2102),
.Y(n_13199)
);

INVx1_ASAP7_75t_L g13200 ( 
.A(n_12771),
.Y(n_13200)
);

INVx1_ASAP7_75t_L g13201 ( 
.A(n_12822),
.Y(n_13201)
);

OAI21x1_ASAP7_75t_L g13202 ( 
.A1(n_12713),
.A2(n_2102),
.B(n_2103),
.Y(n_13202)
);

INVx1_ASAP7_75t_L g13203 ( 
.A(n_12735),
.Y(n_13203)
);

INVx2_ASAP7_75t_L g13204 ( 
.A(n_12902),
.Y(n_13204)
);

INVx1_ASAP7_75t_L g13205 ( 
.A(n_12738),
.Y(n_13205)
);

AOI22xp33_ASAP7_75t_L g13206 ( 
.A1(n_12914),
.A2(n_2106),
.B1(n_2104),
.B2(n_2105),
.Y(n_13206)
);

INVx1_ASAP7_75t_L g13207 ( 
.A(n_12809),
.Y(n_13207)
);

INVx1_ASAP7_75t_L g13208 ( 
.A(n_12820),
.Y(n_13208)
);

INVx2_ASAP7_75t_L g13209 ( 
.A(n_12853),
.Y(n_13209)
);

INVx1_ASAP7_75t_L g13210 ( 
.A(n_12987),
.Y(n_13210)
);

INVx2_ASAP7_75t_L g13211 ( 
.A(n_12960),
.Y(n_13211)
);

HB1xp67_ASAP7_75t_SL g13212 ( 
.A(n_12829),
.Y(n_13212)
);

AND2x4_ASAP7_75t_L g13213 ( 
.A(n_12918),
.B(n_2104),
.Y(n_13213)
);

AOI21xp5_ASAP7_75t_L g13214 ( 
.A1(n_12743),
.A2(n_2106),
.B(n_2107),
.Y(n_13214)
);

INVx2_ASAP7_75t_L g13215 ( 
.A(n_12816),
.Y(n_13215)
);

INVx1_ASAP7_75t_L g13216 ( 
.A(n_12988),
.Y(n_13216)
);

INVx2_ASAP7_75t_L g13217 ( 
.A(n_12816),
.Y(n_13217)
);

AND2x2_ASAP7_75t_L g13218 ( 
.A(n_12924),
.B(n_2108),
.Y(n_13218)
);

AND2x2_ASAP7_75t_L g13219 ( 
.A(n_12980),
.B(n_2108),
.Y(n_13219)
);

AOI221xp5_ASAP7_75t_L g13220 ( 
.A1(n_12959),
.A2(n_12999),
.B1(n_12815),
.B2(n_12871),
.C(n_12726),
.Y(n_13220)
);

INVx1_ASAP7_75t_L g13221 ( 
.A(n_13032),
.Y(n_13221)
);

INVx1_ASAP7_75t_L g13222 ( 
.A(n_12984),
.Y(n_13222)
);

BUFx2_ASAP7_75t_L g13223 ( 
.A(n_13016),
.Y(n_13223)
);

OAI21x1_ASAP7_75t_L g13224 ( 
.A1(n_12778),
.A2(n_2109),
.B(n_2110),
.Y(n_13224)
);

OR2x6_ASAP7_75t_L g13225 ( 
.A(n_12887),
.B(n_12859),
.Y(n_13225)
);

INVx1_ASAP7_75t_L g13226 ( 
.A(n_12979),
.Y(n_13226)
);

OAI21xp5_ASAP7_75t_L g13227 ( 
.A1(n_12945),
.A2(n_2110),
.B(n_2111),
.Y(n_13227)
);

INVx1_ASAP7_75t_L g13228 ( 
.A(n_12789),
.Y(n_13228)
);

AND2x4_ASAP7_75t_L g13229 ( 
.A(n_12981),
.B(n_2111),
.Y(n_13229)
);

AND2x2_ASAP7_75t_L g13230 ( 
.A(n_12776),
.B(n_12786),
.Y(n_13230)
);

AND2x2_ASAP7_75t_L g13231 ( 
.A(n_12806),
.B(n_12702),
.Y(n_13231)
);

OAI21x1_ASAP7_75t_L g13232 ( 
.A1(n_12724),
.A2(n_2112),
.B(n_2113),
.Y(n_13232)
);

INVx1_ASAP7_75t_L g13233 ( 
.A(n_12891),
.Y(n_13233)
);

AND2x4_ASAP7_75t_L g13234 ( 
.A(n_12813),
.B(n_2112),
.Y(n_13234)
);

INVx1_ASAP7_75t_L g13235 ( 
.A(n_12824),
.Y(n_13235)
);

INVx1_ASAP7_75t_L g13236 ( 
.A(n_12839),
.Y(n_13236)
);

INVx1_ASAP7_75t_L g13237 ( 
.A(n_12881),
.Y(n_13237)
);

INVx2_ASAP7_75t_L g13238 ( 
.A(n_12964),
.Y(n_13238)
);

NAND2xp33_ASAP7_75t_R g13239 ( 
.A(n_12975),
.B(n_2113),
.Y(n_13239)
);

INVx1_ASAP7_75t_L g13240 ( 
.A(n_12911),
.Y(n_13240)
);

INVx1_ASAP7_75t_L g13241 ( 
.A(n_12916),
.Y(n_13241)
);

BUFx6f_ASAP7_75t_L g13242 ( 
.A(n_12773),
.Y(n_13242)
);

BUFx2_ASAP7_75t_R g13243 ( 
.A(n_12938),
.Y(n_13243)
);

INVx1_ASAP7_75t_L g13244 ( 
.A(n_12953),
.Y(n_13244)
);

OAI21x1_ASAP7_75t_L g13245 ( 
.A1(n_12856),
.A2(n_2114),
.B(n_2115),
.Y(n_13245)
);

INVx3_ASAP7_75t_L g13246 ( 
.A(n_12912),
.Y(n_13246)
);

INVxp67_ASAP7_75t_SL g13247 ( 
.A(n_12863),
.Y(n_13247)
);

INVx3_ASAP7_75t_L g13248 ( 
.A(n_12944),
.Y(n_13248)
);

INVx1_ASAP7_75t_SL g13249 ( 
.A(n_12712),
.Y(n_13249)
);

HB1xp67_ASAP7_75t_L g13250 ( 
.A(n_12961),
.Y(n_13250)
);

AOI22xp5_ASAP7_75t_L g13251 ( 
.A1(n_12951),
.A2(n_2117),
.B1(n_2115),
.B2(n_2116),
.Y(n_13251)
);

AND2x2_ASAP7_75t_L g13252 ( 
.A(n_12746),
.B(n_2116),
.Y(n_13252)
);

INVx3_ASAP7_75t_L g13253 ( 
.A(n_12887),
.Y(n_13253)
);

NAND2xp5_ASAP7_75t_L g13254 ( 
.A(n_12782),
.B(n_2118),
.Y(n_13254)
);

NAND2xp5_ASAP7_75t_L g13255 ( 
.A(n_12875),
.B(n_2119),
.Y(n_13255)
);

CKINVDCx20_ASAP7_75t_R g13256 ( 
.A(n_12830),
.Y(n_13256)
);

INVx1_ASAP7_75t_L g13257 ( 
.A(n_12821),
.Y(n_13257)
);

NAND2xp5_ASAP7_75t_L g13258 ( 
.A(n_12807),
.B(n_2119),
.Y(n_13258)
);

NOR2x1_ASAP7_75t_SL g13259 ( 
.A(n_12965),
.B(n_2120),
.Y(n_13259)
);

INVx2_ASAP7_75t_L g13260 ( 
.A(n_12716),
.Y(n_13260)
);

INVx1_ASAP7_75t_L g13261 ( 
.A(n_12977),
.Y(n_13261)
);

INVx1_ASAP7_75t_L g13262 ( 
.A(n_12928),
.Y(n_13262)
);

NOR2x1_ASAP7_75t_L g13263 ( 
.A(n_12920),
.B(n_12731),
.Y(n_13263)
);

INVx3_ASAP7_75t_L g13264 ( 
.A(n_12747),
.Y(n_13264)
);

INVx1_ASAP7_75t_L g13265 ( 
.A(n_12928),
.Y(n_13265)
);

AND2x4_ASAP7_75t_L g13266 ( 
.A(n_12840),
.B(n_2120),
.Y(n_13266)
);

OR2x2_ASAP7_75t_L g13267 ( 
.A(n_12862),
.B(n_2121),
.Y(n_13267)
);

AND2x4_ASAP7_75t_L g13268 ( 
.A(n_12795),
.B(n_2121),
.Y(n_13268)
);

INVx1_ASAP7_75t_L g13269 ( 
.A(n_12764),
.Y(n_13269)
);

OAI21x1_ASAP7_75t_L g13270 ( 
.A1(n_12749),
.A2(n_2122),
.B(n_2123),
.Y(n_13270)
);

OAI21xp5_ASAP7_75t_L g13271 ( 
.A1(n_12857),
.A2(n_2122),
.B(n_2123),
.Y(n_13271)
);

INVxp67_ASAP7_75t_L g13272 ( 
.A(n_12970),
.Y(n_13272)
);

INVx1_ASAP7_75t_L g13273 ( 
.A(n_13022),
.Y(n_13273)
);

INVx1_ASAP7_75t_L g13274 ( 
.A(n_12780),
.Y(n_13274)
);

INVx2_ASAP7_75t_L g13275 ( 
.A(n_12689),
.Y(n_13275)
);

AND2x2_ASAP7_75t_L g13276 ( 
.A(n_13035),
.B(n_2124),
.Y(n_13276)
);

HB1xp67_ASAP7_75t_L g13277 ( 
.A(n_12709),
.Y(n_13277)
);

INVx3_ASAP7_75t_L g13278 ( 
.A(n_12896),
.Y(n_13278)
);

AOI22xp33_ASAP7_75t_L g13279 ( 
.A1(n_13021),
.A2(n_2126),
.B1(n_2124),
.B2(n_2125),
.Y(n_13279)
);

OAI22xp5_ASAP7_75t_L g13280 ( 
.A1(n_12711),
.A2(n_2127),
.B1(n_2125),
.B2(n_2126),
.Y(n_13280)
);

BUFx3_ASAP7_75t_L g13281 ( 
.A(n_12838),
.Y(n_13281)
);

AND2x4_ASAP7_75t_L g13282 ( 
.A(n_12737),
.B(n_2127),
.Y(n_13282)
);

INVx1_ASAP7_75t_L g13283 ( 
.A(n_13038),
.Y(n_13283)
);

BUFx3_ASAP7_75t_L g13284 ( 
.A(n_12895),
.Y(n_13284)
);

AND2x2_ASAP7_75t_L g13285 ( 
.A(n_12923),
.B(n_2128),
.Y(n_13285)
);

NAND2xp5_ASAP7_75t_L g13286 ( 
.A(n_12906),
.B(n_2128),
.Y(n_13286)
);

BUFx4f_ASAP7_75t_L g13287 ( 
.A(n_13002),
.Y(n_13287)
);

INVx2_ASAP7_75t_L g13288 ( 
.A(n_12952),
.Y(n_13288)
);

OAI21xp5_ASAP7_75t_L g13289 ( 
.A1(n_12752),
.A2(n_2129),
.B(n_2130),
.Y(n_13289)
);

INVx1_ASAP7_75t_L g13290 ( 
.A(n_12810),
.Y(n_13290)
);

AND2x2_ASAP7_75t_L g13291 ( 
.A(n_12869),
.B(n_2129),
.Y(n_13291)
);

INVx1_ASAP7_75t_L g13292 ( 
.A(n_12844),
.Y(n_13292)
);

INVx2_ASAP7_75t_L g13293 ( 
.A(n_12725),
.Y(n_13293)
);

INVx3_ASAP7_75t_L g13294 ( 
.A(n_12781),
.Y(n_13294)
);

INVx1_ASAP7_75t_L g13295 ( 
.A(n_12974),
.Y(n_13295)
);

NAND2xp5_ASAP7_75t_L g13296 ( 
.A(n_12948),
.B(n_2130),
.Y(n_13296)
);

BUFx3_ASAP7_75t_L g13297 ( 
.A(n_12998),
.Y(n_13297)
);

INVx1_ASAP7_75t_L g13298 ( 
.A(n_12826),
.Y(n_13298)
);

INVx1_ASAP7_75t_L g13299 ( 
.A(n_12828),
.Y(n_13299)
);

INVx1_ASAP7_75t_L g13300 ( 
.A(n_12831),
.Y(n_13300)
);

INVx1_ASAP7_75t_L g13301 ( 
.A(n_12837),
.Y(n_13301)
);

INVx2_ASAP7_75t_L g13302 ( 
.A(n_12941),
.Y(n_13302)
);

INVx3_ASAP7_75t_L g13303 ( 
.A(n_12903),
.Y(n_13303)
);

INVx1_ASAP7_75t_L g13304 ( 
.A(n_12874),
.Y(n_13304)
);

INVx2_ASAP7_75t_L g13305 ( 
.A(n_13003),
.Y(n_13305)
);

OA21x2_ASAP7_75t_L g13306 ( 
.A1(n_12833),
.A2(n_2131),
.B(n_2132),
.Y(n_13306)
);

OR2x2_ASAP7_75t_L g13307 ( 
.A(n_12869),
.B(n_2131),
.Y(n_13307)
);

INVx1_ASAP7_75t_L g13308 ( 
.A(n_12885),
.Y(n_13308)
);

INVx1_ASAP7_75t_L g13309 ( 
.A(n_12892),
.Y(n_13309)
);

BUFx3_ASAP7_75t_L g13310 ( 
.A(n_12865),
.Y(n_13310)
);

AND2x2_ASAP7_75t_L g13311 ( 
.A(n_12913),
.B(n_2132),
.Y(n_13311)
);

INVx2_ASAP7_75t_L g13312 ( 
.A(n_12968),
.Y(n_13312)
);

OAI21x1_ASAP7_75t_L g13313 ( 
.A1(n_12877),
.A2(n_2133),
.B(n_2134),
.Y(n_13313)
);

INVx1_ASAP7_75t_L g13314 ( 
.A(n_12898),
.Y(n_13314)
);

HB1xp67_ASAP7_75t_L g13315 ( 
.A(n_12834),
.Y(n_13315)
);

INVx1_ASAP7_75t_L g13316 ( 
.A(n_12968),
.Y(n_13316)
);

INVx2_ASAP7_75t_L g13317 ( 
.A(n_12744),
.Y(n_13317)
);

OR2x6_ASAP7_75t_L g13318 ( 
.A(n_12893),
.B(n_2133),
.Y(n_13318)
);

BUFx8_ASAP7_75t_L g13319 ( 
.A(n_12995),
.Y(n_13319)
);

INVx1_ASAP7_75t_SL g13320 ( 
.A(n_12860),
.Y(n_13320)
);

INVx1_ASAP7_75t_L g13321 ( 
.A(n_12758),
.Y(n_13321)
);

INVx2_ASAP7_75t_L g13322 ( 
.A(n_12759),
.Y(n_13322)
);

HB1xp67_ASAP7_75t_L g13323 ( 
.A(n_12842),
.Y(n_13323)
);

INVx2_ASAP7_75t_SL g13324 ( 
.A(n_12937),
.Y(n_13324)
);

NAND2xp5_ASAP7_75t_L g13325 ( 
.A(n_12868),
.B(n_2135),
.Y(n_13325)
);

INVx1_ASAP7_75t_L g13326 ( 
.A(n_12761),
.Y(n_13326)
);

INVx2_ASAP7_75t_SL g13327 ( 
.A(n_12972),
.Y(n_13327)
);

INVxp67_ASAP7_75t_L g13328 ( 
.A(n_12768),
.Y(n_13328)
);

INVx1_ASAP7_75t_L g13329 ( 
.A(n_12772),
.Y(n_13329)
);

OAI21x1_ASAP7_75t_L g13330 ( 
.A1(n_12832),
.A2(n_2135),
.B(n_2136),
.Y(n_13330)
);

INVx2_ASAP7_75t_L g13331 ( 
.A(n_12845),
.Y(n_13331)
);

INVx2_ASAP7_75t_L g13332 ( 
.A(n_12851),
.Y(n_13332)
);

INVxp67_ASAP7_75t_L g13333 ( 
.A(n_13028),
.Y(n_13333)
);

INVx3_ASAP7_75t_L g13334 ( 
.A(n_12823),
.Y(n_13334)
);

INVx1_ASAP7_75t_L g13335 ( 
.A(n_12858),
.Y(n_13335)
);

NAND2xp5_ASAP7_75t_L g13336 ( 
.A(n_12720),
.B(n_12933),
.Y(n_13336)
);

HB1xp67_ASAP7_75t_L g13337 ( 
.A(n_12864),
.Y(n_13337)
);

OA21x2_ASAP7_75t_L g13338 ( 
.A1(n_12873),
.A2(n_2136),
.B(n_2137),
.Y(n_13338)
);

INVx1_ASAP7_75t_L g13339 ( 
.A(n_12880),
.Y(n_13339)
);

OR2x2_ASAP7_75t_L g13340 ( 
.A(n_12723),
.B(n_2137),
.Y(n_13340)
);

INVx1_ASAP7_75t_L g13341 ( 
.A(n_13020),
.Y(n_13341)
);

INVx2_ASAP7_75t_L g13342 ( 
.A(n_12930),
.Y(n_13342)
);

INVx1_ASAP7_75t_L g13343 ( 
.A(n_13024),
.Y(n_13343)
);

HB1xp67_ASAP7_75t_L g13344 ( 
.A(n_12973),
.Y(n_13344)
);

INVx8_ASAP7_75t_L g13345 ( 
.A(n_13013),
.Y(n_13345)
);

HB1xp67_ASAP7_75t_L g13346 ( 
.A(n_13006),
.Y(n_13346)
);

INVx1_ASAP7_75t_L g13347 ( 
.A(n_12985),
.Y(n_13347)
);

AND2x2_ASAP7_75t_L g13348 ( 
.A(n_12784),
.B(n_2138),
.Y(n_13348)
);

INVx1_ASAP7_75t_L g13349 ( 
.A(n_13011),
.Y(n_13349)
);

NAND3x1_ASAP7_75t_L g13350 ( 
.A(n_12698),
.B(n_2138),
.C(n_2139),
.Y(n_13350)
);

INVx2_ASAP7_75t_L g13351 ( 
.A(n_13012),
.Y(n_13351)
);

INVx2_ASAP7_75t_L g13352 ( 
.A(n_13000),
.Y(n_13352)
);

INVx3_ASAP7_75t_L g13353 ( 
.A(n_12997),
.Y(n_13353)
);

INVx2_ASAP7_75t_L g13354 ( 
.A(n_13005),
.Y(n_13354)
);

AOI21x1_ASAP7_75t_L g13355 ( 
.A1(n_12841),
.A2(n_2139),
.B(n_2140),
.Y(n_13355)
);

BUFx4f_ASAP7_75t_SL g13356 ( 
.A(n_12847),
.Y(n_13356)
);

AOI221xp5_ASAP7_75t_L g13357 ( 
.A1(n_12861),
.A2(n_2142),
.B1(n_2140),
.B2(n_2141),
.C(n_2143),
.Y(n_13357)
);

INVx1_ASAP7_75t_L g13358 ( 
.A(n_13027),
.Y(n_13358)
);

INVx3_ASAP7_75t_L g13359 ( 
.A(n_12882),
.Y(n_13359)
);

INVx1_ASAP7_75t_L g13360 ( 
.A(n_13015),
.Y(n_13360)
);

OAI21x1_ASAP7_75t_L g13361 ( 
.A1(n_12692),
.A2(n_2141),
.B(n_2142),
.Y(n_13361)
);

OAI21x1_ASAP7_75t_L g13362 ( 
.A1(n_12888),
.A2(n_2143),
.B(n_2144),
.Y(n_13362)
);

HB1xp67_ASAP7_75t_L g13363 ( 
.A(n_12855),
.Y(n_13363)
);

INVx1_ASAP7_75t_L g13364 ( 
.A(n_12796),
.Y(n_13364)
);

INVx1_ASAP7_75t_L g13365 ( 
.A(n_13018),
.Y(n_13365)
);

BUFx2_ASAP7_75t_L g13366 ( 
.A(n_12852),
.Y(n_13366)
);

BUFx6f_ASAP7_75t_L g13367 ( 
.A(n_12907),
.Y(n_13367)
);

INVx2_ASAP7_75t_L g13368 ( 
.A(n_13034),
.Y(n_13368)
);

INVx1_ASAP7_75t_L g13369 ( 
.A(n_13030),
.Y(n_13369)
);

INVx2_ASAP7_75t_L g13370 ( 
.A(n_13029),
.Y(n_13370)
);

BUFx2_ASAP7_75t_L g13371 ( 
.A(n_12884),
.Y(n_13371)
);

OAI21x1_ASAP7_75t_L g13372 ( 
.A1(n_12733),
.A2(n_2145),
.B(n_2146),
.Y(n_13372)
);

INVx1_ASAP7_75t_L g13373 ( 
.A(n_12882),
.Y(n_13373)
);

NAND2x1p5_ASAP7_75t_L g13374 ( 
.A(n_13019),
.B(n_2145),
.Y(n_13374)
);

NAND2xp5_ASAP7_75t_L g13375 ( 
.A(n_12785),
.B(n_2147),
.Y(n_13375)
);

AND2x2_ASAP7_75t_L g13376 ( 
.A(n_12897),
.B(n_12910),
.Y(n_13376)
);

INVx2_ASAP7_75t_L g13377 ( 
.A(n_13017),
.Y(n_13377)
);

INVx1_ASAP7_75t_L g13378 ( 
.A(n_12969),
.Y(n_13378)
);

INVx1_ASAP7_75t_L g13379 ( 
.A(n_12983),
.Y(n_13379)
);

OR2x6_ASAP7_75t_L g13380 ( 
.A(n_12957),
.B(n_2147),
.Y(n_13380)
);

OA21x2_ASAP7_75t_L g13381 ( 
.A1(n_12763),
.A2(n_2148),
.B(n_2149),
.Y(n_13381)
);

AOI21x1_ASAP7_75t_L g13382 ( 
.A1(n_12934),
.A2(n_2149),
.B(n_2150),
.Y(n_13382)
);

INVx2_ASAP7_75t_L g13383 ( 
.A(n_13026),
.Y(n_13383)
);

INVx1_ASAP7_75t_L g13384 ( 
.A(n_12949),
.Y(n_13384)
);

INVx1_ASAP7_75t_L g13385 ( 
.A(n_12992),
.Y(n_13385)
);

INVx2_ASAP7_75t_L g13386 ( 
.A(n_13036),
.Y(n_13386)
);

INVx1_ASAP7_75t_L g13387 ( 
.A(n_12943),
.Y(n_13387)
);

INVx1_ASAP7_75t_L g13388 ( 
.A(n_12989),
.Y(n_13388)
);

AOI22xp33_ASAP7_75t_L g13389 ( 
.A1(n_13383),
.A2(n_13001),
.B1(n_13025),
.B2(n_12993),
.Y(n_13389)
);

AOI22xp33_ASAP7_75t_L g13390 ( 
.A1(n_13168),
.A2(n_12908),
.B1(n_2152),
.B2(n_2150),
.Y(n_13390)
);

OAI221xp5_ASAP7_75t_L g13391 ( 
.A1(n_13251),
.A2(n_2153),
.B1(n_2151),
.B2(n_2152),
.C(n_2154),
.Y(n_13391)
);

AOI221xp5_ASAP7_75t_L g13392 ( 
.A1(n_13277),
.A2(n_2155),
.B1(n_2153),
.B2(n_2154),
.C(n_2156),
.Y(n_13392)
);

INVx3_ASAP7_75t_L g13393 ( 
.A(n_13107),
.Y(n_13393)
);

AOI221xp5_ASAP7_75t_L g13394 ( 
.A1(n_13336),
.A2(n_2158),
.B1(n_2156),
.B2(n_2157),
.C(n_2159),
.Y(n_13394)
);

AOI221xp5_ASAP7_75t_L g13395 ( 
.A1(n_13196),
.A2(n_2160),
.B1(n_2157),
.B2(n_2159),
.C(n_2161),
.Y(n_13395)
);

BUFx4f_ASAP7_75t_SL g13396 ( 
.A(n_13129),
.Y(n_13396)
);

AOI22xp33_ASAP7_75t_L g13397 ( 
.A1(n_13220),
.A2(n_2164),
.B1(n_2162),
.B2(n_2163),
.Y(n_13397)
);

AOI22xp33_ASAP7_75t_L g13398 ( 
.A1(n_13377),
.A2(n_2164),
.B1(n_2162),
.B2(n_2163),
.Y(n_13398)
);

INVx2_ASAP7_75t_L g13399 ( 
.A(n_13154),
.Y(n_13399)
);

AOI22xp33_ASAP7_75t_L g13400 ( 
.A1(n_13150),
.A2(n_2167),
.B1(n_2165),
.B2(n_2166),
.Y(n_13400)
);

OAI21x1_ASAP7_75t_L g13401 ( 
.A1(n_13113),
.A2(n_2165),
.B(n_2168),
.Y(n_13401)
);

AND2x4_ASAP7_75t_L g13402 ( 
.A(n_13147),
.B(n_2169),
.Y(n_13402)
);

BUFx12f_ASAP7_75t_SL g13403 ( 
.A(n_13098),
.Y(n_13403)
);

AOI22xp33_ASAP7_75t_L g13404 ( 
.A1(n_13369),
.A2(n_2171),
.B1(n_2169),
.B2(n_2170),
.Y(n_13404)
);

AOI21xp5_ASAP7_75t_L g13405 ( 
.A1(n_13291),
.A2(n_2170),
.B(n_2171),
.Y(n_13405)
);

OAI22xp33_ASAP7_75t_SL g13406 ( 
.A1(n_13349),
.A2(n_2174),
.B1(n_2172),
.B2(n_2173),
.Y(n_13406)
);

OAI221xp5_ASAP7_75t_L g13407 ( 
.A1(n_13239),
.A2(n_2174),
.B1(n_2172),
.B2(n_2173),
.C(n_2175),
.Y(n_13407)
);

AND2x2_ASAP7_75t_L g13408 ( 
.A(n_13101),
.B(n_2175),
.Y(n_13408)
);

BUFx3_ASAP7_75t_L g13409 ( 
.A(n_13086),
.Y(n_13409)
);

OAI22xp5_ASAP7_75t_L g13410 ( 
.A1(n_13142),
.A2(n_2178),
.B1(n_2176),
.B2(n_2177),
.Y(n_13410)
);

AOI221xp5_ASAP7_75t_L g13411 ( 
.A1(n_13042),
.A2(n_2178),
.B1(n_2176),
.B2(n_2177),
.C(n_2179),
.Y(n_13411)
);

OAI21x1_ASAP7_75t_L g13412 ( 
.A1(n_13067),
.A2(n_2179),
.B(n_2180),
.Y(n_13412)
);

AOI21xp5_ASAP7_75t_L g13413 ( 
.A1(n_13307),
.A2(n_2181),
.B(n_2182),
.Y(n_13413)
);

HB1xp67_ASAP7_75t_L g13414 ( 
.A(n_13046),
.Y(n_13414)
);

AOI22xp33_ASAP7_75t_SL g13415 ( 
.A1(n_13189),
.A2(n_2183),
.B1(n_2181),
.B2(n_2182),
.Y(n_13415)
);

AND2x2_ASAP7_75t_L g13416 ( 
.A(n_13045),
.B(n_2183),
.Y(n_13416)
);

INVx1_ASAP7_75t_L g13417 ( 
.A(n_13097),
.Y(n_13417)
);

OAI31xp33_ASAP7_75t_SL g13418 ( 
.A1(n_13247),
.A2(n_2186),
.A3(n_2184),
.B(n_2185),
.Y(n_13418)
);

OR2x2_ASAP7_75t_L g13419 ( 
.A(n_13187),
.B(n_2185),
.Y(n_13419)
);

OAI22xp5_ASAP7_75t_L g13420 ( 
.A1(n_13371),
.A2(n_2189),
.B1(n_2187),
.B2(n_2188),
.Y(n_13420)
);

INVx1_ASAP7_75t_L g13421 ( 
.A(n_13162),
.Y(n_13421)
);

AOI22xp33_ASAP7_75t_L g13422 ( 
.A1(n_13384),
.A2(n_2190),
.B1(n_2188),
.B2(n_2189),
.Y(n_13422)
);

INVx2_ASAP7_75t_SL g13423 ( 
.A(n_13319),
.Y(n_13423)
);

AOI22xp5_ASAP7_75t_L g13424 ( 
.A1(n_13256),
.A2(n_2192),
.B1(n_2190),
.B2(n_2191),
.Y(n_13424)
);

INVx1_ASAP7_75t_L g13425 ( 
.A(n_13124),
.Y(n_13425)
);

OR2x2_ASAP7_75t_L g13426 ( 
.A(n_13172),
.B(n_2191),
.Y(n_13426)
);

INVx1_ASAP7_75t_L g13427 ( 
.A(n_13104),
.Y(n_13427)
);

OAI22xp33_ASAP7_75t_L g13428 ( 
.A1(n_13225),
.A2(n_2196),
.B1(n_2193),
.B2(n_2195),
.Y(n_13428)
);

NAND2xp5_ASAP7_75t_L g13429 ( 
.A(n_13365),
.B(n_2193),
.Y(n_13429)
);

AOI22xp33_ASAP7_75t_SL g13430 ( 
.A1(n_13164),
.A2(n_2197),
.B1(n_2195),
.B2(n_2196),
.Y(n_13430)
);

AO31x2_ASAP7_75t_L g13431 ( 
.A1(n_13146),
.A2(n_2201),
.A3(n_2198),
.B(n_2200),
.Y(n_13431)
);

INVx2_ASAP7_75t_L g13432 ( 
.A(n_13161),
.Y(n_13432)
);

AOI22xp33_ASAP7_75t_L g13433 ( 
.A1(n_13360),
.A2(n_2201),
.B1(n_2198),
.B2(n_2200),
.Y(n_13433)
);

AOI22xp33_ASAP7_75t_SL g13434 ( 
.A1(n_13167),
.A2(n_13145),
.B1(n_13137),
.B2(n_13223),
.Y(n_13434)
);

AND2x4_ASAP7_75t_L g13435 ( 
.A(n_13088),
.B(n_2202),
.Y(n_13435)
);

OAI22xp5_ASAP7_75t_L g13436 ( 
.A1(n_13366),
.A2(n_2204),
.B1(n_2202),
.B2(n_2203),
.Y(n_13436)
);

OAI211xp5_ASAP7_75t_SL g13437 ( 
.A1(n_13328),
.A2(n_2205),
.B(n_2203),
.C(n_2204),
.Y(n_13437)
);

AND2x2_ASAP7_75t_L g13438 ( 
.A(n_13070),
.B(n_2205),
.Y(n_13438)
);

AOI22xp33_ASAP7_75t_L g13439 ( 
.A1(n_13222),
.A2(n_2208),
.B1(n_2206),
.B2(n_2207),
.Y(n_13439)
);

AOI222xp33_ASAP7_75t_L g13440 ( 
.A1(n_13119),
.A2(n_2208),
.B1(n_2210),
.B2(n_2206),
.C1(n_2207),
.C2(n_2209),
.Y(n_13440)
);

AOI22xp33_ASAP7_75t_L g13441 ( 
.A1(n_13065),
.A2(n_2212),
.B1(n_2209),
.B2(n_2211),
.Y(n_13441)
);

OA21x2_ASAP7_75t_L g13442 ( 
.A1(n_13149),
.A2(n_13209),
.B(n_13200),
.Y(n_13442)
);

OAI211xp5_ASAP7_75t_SL g13443 ( 
.A1(n_13170),
.A2(n_13071),
.B(n_13094),
.C(n_13263),
.Y(n_13443)
);

AND2x2_ASAP7_75t_L g13444 ( 
.A(n_13122),
.B(n_2211),
.Y(n_13444)
);

AOI21xp5_ASAP7_75t_SL g13445 ( 
.A1(n_13099),
.A2(n_2212),
.B(n_2213),
.Y(n_13445)
);

AOI22xp33_ASAP7_75t_L g13446 ( 
.A1(n_13188),
.A2(n_2215),
.B1(n_2213),
.B2(n_2214),
.Y(n_13446)
);

CKINVDCx20_ASAP7_75t_R g13447 ( 
.A(n_13117),
.Y(n_13447)
);

OAI221xp5_ASAP7_75t_L g13448 ( 
.A1(n_13044),
.A2(n_2217),
.B1(n_2214),
.B2(n_2216),
.C(n_2218),
.Y(n_13448)
);

AND2x2_ASAP7_75t_L g13449 ( 
.A(n_13230),
.B(n_13072),
.Y(n_13449)
);

OAI221xp5_ASAP7_75t_SL g13450 ( 
.A1(n_13225),
.A2(n_2220),
.B1(n_2218),
.B2(n_2219),
.C(n_2221),
.Y(n_13450)
);

AND2x4_ASAP7_75t_SL g13451 ( 
.A(n_13110),
.B(n_2219),
.Y(n_13451)
);

INVx1_ASAP7_75t_L g13452 ( 
.A(n_13108),
.Y(n_13452)
);

OAI22xp5_ASAP7_75t_L g13453 ( 
.A1(n_13163),
.A2(n_2223),
.B1(n_2221),
.B2(n_2222),
.Y(n_13453)
);

NAND3xp33_ASAP7_75t_L g13454 ( 
.A(n_13388),
.B(n_2222),
.C(n_2224),
.Y(n_13454)
);

INVx1_ASAP7_75t_L g13455 ( 
.A(n_13112),
.Y(n_13455)
);

OAI22xp5_ASAP7_75t_L g13456 ( 
.A1(n_13127),
.A2(n_2227),
.B1(n_2225),
.B2(n_2226),
.Y(n_13456)
);

OR2x2_ASAP7_75t_L g13457 ( 
.A(n_13320),
.B(n_2225),
.Y(n_13457)
);

AOI221xp5_ASAP7_75t_SL g13458 ( 
.A1(n_13214),
.A2(n_2228),
.B1(n_2226),
.B2(n_2227),
.C(n_2229),
.Y(n_13458)
);

OA21x2_ASAP7_75t_L g13459 ( 
.A1(n_13358),
.A2(n_2228),
.B(n_2230),
.Y(n_13459)
);

INVx1_ASAP7_75t_L g13460 ( 
.A(n_13114),
.Y(n_13460)
);

OR2x6_ASAP7_75t_L g13461 ( 
.A(n_13041),
.B(n_2231),
.Y(n_13461)
);

INVx1_ASAP7_75t_L g13462 ( 
.A(n_13157),
.Y(n_13462)
);

INVx1_ASAP7_75t_L g13463 ( 
.A(n_13125),
.Y(n_13463)
);

NOR2x1_ASAP7_75t_L g13464 ( 
.A(n_13048),
.B(n_2231),
.Y(n_13464)
);

AND2x2_ASAP7_75t_L g13465 ( 
.A(n_13053),
.B(n_2232),
.Y(n_13465)
);

OAI211xp5_ASAP7_75t_SL g13466 ( 
.A1(n_13264),
.A2(n_2235),
.B(n_2233),
.C(n_2234),
.Y(n_13466)
);

INVx1_ASAP7_75t_L g13467 ( 
.A(n_13069),
.Y(n_13467)
);

BUFx6f_ASAP7_75t_L g13468 ( 
.A(n_13140),
.Y(n_13468)
);

INVx1_ASAP7_75t_L g13469 ( 
.A(n_13171),
.Y(n_13469)
);

AOI22xp33_ASAP7_75t_L g13470 ( 
.A1(n_13194),
.A2(n_2236),
.B1(n_2233),
.B2(n_2234),
.Y(n_13470)
);

OA21x2_ASAP7_75t_L g13471 ( 
.A1(n_13156),
.A2(n_2236),
.B(n_2237),
.Y(n_13471)
);

AOI22xp33_ASAP7_75t_L g13472 ( 
.A1(n_13261),
.A2(n_2240),
.B1(n_2238),
.B2(n_2239),
.Y(n_13472)
);

CKINVDCx5p33_ASAP7_75t_R g13473 ( 
.A(n_13212),
.Y(n_13473)
);

OAI22xp5_ASAP7_75t_L g13474 ( 
.A1(n_13324),
.A2(n_2241),
.B1(n_2238),
.B2(n_2240),
.Y(n_13474)
);

OAI22xp5_ASAP7_75t_L g13475 ( 
.A1(n_13303),
.A2(n_2243),
.B1(n_2241),
.B2(n_2242),
.Y(n_13475)
);

AOI222xp33_ASAP7_75t_L g13476 ( 
.A1(n_13047),
.A2(n_2246),
.B1(n_2248),
.B2(n_2244),
.C1(n_2245),
.C2(n_2247),
.Y(n_13476)
);

AND2x2_ASAP7_75t_L g13477 ( 
.A(n_13043),
.B(n_2244),
.Y(n_13477)
);

AOI22xp5_ASAP7_75t_SL g13478 ( 
.A1(n_13385),
.A2(n_2248),
.B1(n_2245),
.B2(n_2246),
.Y(n_13478)
);

AOI22xp33_ASAP7_75t_L g13479 ( 
.A1(n_13158),
.A2(n_2252),
.B1(n_2249),
.B2(n_2250),
.Y(n_13479)
);

AOI22xp33_ASAP7_75t_L g13480 ( 
.A1(n_13160),
.A2(n_2253),
.B1(n_2249),
.B2(n_2252),
.Y(n_13480)
);

NOR2xp33_ASAP7_75t_L g13481 ( 
.A(n_13356),
.B(n_2253),
.Y(n_13481)
);

OR2x2_ASAP7_75t_L g13482 ( 
.A(n_13267),
.B(n_2254),
.Y(n_13482)
);

INVx1_ASAP7_75t_L g13483 ( 
.A(n_13176),
.Y(n_13483)
);

A2O1A1Ixp33_ASAP7_75t_L g13484 ( 
.A1(n_13289),
.A2(n_2256),
.B(n_2254),
.C(n_2255),
.Y(n_13484)
);

OAI22xp5_ASAP7_75t_L g13485 ( 
.A1(n_13343),
.A2(n_2257),
.B1(n_2255),
.B2(n_2256),
.Y(n_13485)
);

HB1xp67_ASAP7_75t_L g13486 ( 
.A(n_13346),
.Y(n_13486)
);

BUFx5_ASAP7_75t_L g13487 ( 
.A(n_13285),
.Y(n_13487)
);

CKINVDCx20_ASAP7_75t_R g13488 ( 
.A(n_13281),
.Y(n_13488)
);

AOI21xp5_ASAP7_75t_L g13489 ( 
.A1(n_13255),
.A2(n_2258),
.B(n_2259),
.Y(n_13489)
);

NOR3xp33_ASAP7_75t_L g13490 ( 
.A(n_13089),
.B(n_2258),
.C(n_2260),
.Y(n_13490)
);

OAI221xp5_ASAP7_75t_L g13491 ( 
.A1(n_13305),
.A2(n_2262),
.B1(n_2260),
.B2(n_2261),
.C(n_2263),
.Y(n_13491)
);

AND2x2_ASAP7_75t_L g13492 ( 
.A(n_13143),
.B(n_2261),
.Y(n_13492)
);

INVx2_ASAP7_75t_L g13493 ( 
.A(n_13259),
.Y(n_13493)
);

O2A1O1Ixp33_ASAP7_75t_L g13494 ( 
.A1(n_13363),
.A2(n_2266),
.B(n_2264),
.C(n_2265),
.Y(n_13494)
);

AOI211xp5_ASAP7_75t_L g13495 ( 
.A1(n_13128),
.A2(n_2267),
.B(n_2264),
.C(n_2266),
.Y(n_13495)
);

AND2x2_ASAP7_75t_L g13496 ( 
.A(n_13096),
.B(n_2268),
.Y(n_13496)
);

NOR2xp33_ASAP7_75t_SL g13497 ( 
.A(n_13243),
.B(n_2268),
.Y(n_13497)
);

CKINVDCx5p33_ASAP7_75t_R g13498 ( 
.A(n_13049),
.Y(n_13498)
);

AOI22xp33_ASAP7_75t_SL g13499 ( 
.A1(n_13288),
.A2(n_2271),
.B1(n_2269),
.B2(n_2270),
.Y(n_13499)
);

OAI221xp5_ASAP7_75t_L g13500 ( 
.A1(n_13302),
.A2(n_2271),
.B1(n_2269),
.B2(n_2270),
.C(n_2272),
.Y(n_13500)
);

INVx3_ASAP7_75t_L g13501 ( 
.A(n_13242),
.Y(n_13501)
);

BUFx2_ASAP7_75t_L g13502 ( 
.A(n_13287),
.Y(n_13502)
);

OAI221xp5_ASAP7_75t_L g13503 ( 
.A1(n_13370),
.A2(n_2274),
.B1(n_2272),
.B2(n_2273),
.C(n_2275),
.Y(n_13503)
);

OAI21x1_ASAP7_75t_L g13504 ( 
.A1(n_13153),
.A2(n_2273),
.B(n_2274),
.Y(n_13504)
);

OAI211xp5_ASAP7_75t_L g13505 ( 
.A1(n_13275),
.A2(n_2277),
.B(n_2275),
.C(n_2276),
.Y(n_13505)
);

INVx2_ASAP7_75t_L g13506 ( 
.A(n_13151),
.Y(n_13506)
);

INVx1_ASAP7_75t_L g13507 ( 
.A(n_13056),
.Y(n_13507)
);

INVx1_ASAP7_75t_L g13508 ( 
.A(n_13058),
.Y(n_13508)
);

OAI22xp5_ASAP7_75t_L g13509 ( 
.A1(n_13283),
.A2(n_2278),
.B1(n_2276),
.B2(n_2277),
.Y(n_13509)
);

AND2x2_ASAP7_75t_L g13510 ( 
.A(n_13109),
.B(n_13111),
.Y(n_13510)
);

INVx1_ASAP7_75t_L g13511 ( 
.A(n_13061),
.Y(n_13511)
);

AND2x2_ASAP7_75t_L g13512 ( 
.A(n_13085),
.B(n_2278),
.Y(n_13512)
);

OAI21x1_ASAP7_75t_L g13513 ( 
.A1(n_13190),
.A2(n_2279),
.B(n_2280),
.Y(n_13513)
);

OAI22xp5_ASAP7_75t_L g13514 ( 
.A1(n_13378),
.A2(n_2281),
.B1(n_2279),
.B2(n_2280),
.Y(n_13514)
);

AOI22xp33_ASAP7_75t_L g13515 ( 
.A1(n_13165),
.A2(n_2283),
.B1(n_2281),
.B2(n_2282),
.Y(n_13515)
);

AOI22xp33_ASAP7_75t_L g13516 ( 
.A1(n_13273),
.A2(n_2285),
.B1(n_2283),
.B2(n_2284),
.Y(n_13516)
);

AND2x2_ASAP7_75t_L g13517 ( 
.A(n_13103),
.B(n_2286),
.Y(n_13517)
);

AOI22xp33_ASAP7_75t_L g13518 ( 
.A1(n_13237),
.A2(n_2289),
.B1(n_2286),
.B2(n_2287),
.Y(n_13518)
);

OR2x2_ASAP7_75t_L g13519 ( 
.A(n_13201),
.B(n_2289),
.Y(n_13519)
);

AOI22xp33_ASAP7_75t_L g13520 ( 
.A1(n_13240),
.A2(n_13241),
.B1(n_13257),
.B2(n_13244),
.Y(n_13520)
);

OAI221xp5_ASAP7_75t_SL g13521 ( 
.A1(n_13318),
.A2(n_2292),
.B1(n_2290),
.B2(n_2291),
.C(n_2293),
.Y(n_13521)
);

OAI22xp33_ASAP7_75t_L g13522 ( 
.A1(n_13318),
.A2(n_2292),
.B1(n_2290),
.B2(n_2291),
.Y(n_13522)
);

INVx2_ASAP7_75t_SL g13523 ( 
.A(n_13345),
.Y(n_13523)
);

AND2x2_ASAP7_75t_L g13524 ( 
.A(n_13367),
.B(n_2293),
.Y(n_13524)
);

AOI22xp5_ASAP7_75t_L g13525 ( 
.A1(n_13350),
.A2(n_13379),
.B1(n_13380),
.B2(n_13376),
.Y(n_13525)
);

INVx2_ASAP7_75t_L g13526 ( 
.A(n_13253),
.Y(n_13526)
);

INVx3_ASAP7_75t_L g13527 ( 
.A(n_13242),
.Y(n_13527)
);

INVx3_ASAP7_75t_L g13528 ( 
.A(n_13166),
.Y(n_13528)
);

NOR2xp33_ASAP7_75t_L g13529 ( 
.A(n_13177),
.B(n_2295),
.Y(n_13529)
);

OAI21xp5_ASAP7_75t_L g13530 ( 
.A1(n_13280),
.A2(n_2295),
.B(n_2296),
.Y(n_13530)
);

AOI221xp5_ASAP7_75t_L g13531 ( 
.A1(n_13250),
.A2(n_2298),
.B1(n_2296),
.B2(n_2297),
.C(n_2299),
.Y(n_13531)
);

INVx1_ASAP7_75t_L g13532 ( 
.A(n_13075),
.Y(n_13532)
);

BUFx2_ASAP7_75t_L g13533 ( 
.A(n_13367),
.Y(n_13533)
);

AOI222xp33_ASAP7_75t_L g13534 ( 
.A1(n_13051),
.A2(n_2300),
.B1(n_2302),
.B2(n_2297),
.C1(n_2299),
.C2(n_2301),
.Y(n_13534)
);

NAND3xp33_ASAP7_75t_L g13535 ( 
.A(n_13357),
.B(n_2300),
.C(n_2302),
.Y(n_13535)
);

OAI21xp33_ASAP7_75t_L g13536 ( 
.A1(n_13387),
.A2(n_13183),
.B(n_13181),
.Y(n_13536)
);

BUFx2_ASAP7_75t_L g13537 ( 
.A(n_13246),
.Y(n_13537)
);

AOI22xp33_ASAP7_75t_SL g13538 ( 
.A1(n_13359),
.A2(n_2305),
.B1(n_2303),
.B2(n_2304),
.Y(n_13538)
);

AOI22xp5_ASAP7_75t_L g13539 ( 
.A1(n_13380),
.A2(n_2306),
.B1(n_2303),
.B2(n_2305),
.Y(n_13539)
);

OAI221xp5_ASAP7_75t_L g13540 ( 
.A1(n_13272),
.A2(n_2308),
.B1(n_2306),
.B2(n_2307),
.C(n_2309),
.Y(n_13540)
);

AOI21xp5_ASAP7_75t_L g13541 ( 
.A1(n_13178),
.A2(n_2307),
.B(n_2308),
.Y(n_13541)
);

NAND2xp5_ASAP7_75t_L g13542 ( 
.A(n_13344),
.B(n_13152),
.Y(n_13542)
);

BUFx2_ASAP7_75t_L g13543 ( 
.A(n_13284),
.Y(n_13543)
);

AOI22xp33_ASAP7_75t_L g13544 ( 
.A1(n_13312),
.A2(n_2312),
.B1(n_2310),
.B2(n_2311),
.Y(n_13544)
);

AOI22xp33_ASAP7_75t_L g13545 ( 
.A1(n_13091),
.A2(n_13052),
.B1(n_13054),
.B2(n_13316),
.Y(n_13545)
);

INVx2_ASAP7_75t_L g13546 ( 
.A(n_13278),
.Y(n_13546)
);

INVx6_ASAP7_75t_L g13547 ( 
.A(n_13130),
.Y(n_13547)
);

INVx1_ASAP7_75t_L g13548 ( 
.A(n_13077),
.Y(n_13548)
);

AOI21xp5_ASAP7_75t_L g13549 ( 
.A1(n_13258),
.A2(n_2311),
.B(n_2312),
.Y(n_13549)
);

OAI221xp5_ASAP7_75t_L g13550 ( 
.A1(n_13374),
.A2(n_2315),
.B1(n_2313),
.B2(n_2314),
.C(n_2316),
.Y(n_13550)
);

AOI21xp5_ASAP7_75t_L g13551 ( 
.A1(n_13286),
.A2(n_2314),
.B(n_2315),
.Y(n_13551)
);

OAI21xp5_ASAP7_75t_SL g13552 ( 
.A1(n_13184),
.A2(n_2316),
.B(n_2317),
.Y(n_13552)
);

INVx1_ASAP7_75t_L g13553 ( 
.A(n_13079),
.Y(n_13553)
);

AND2x2_ASAP7_75t_L g13554 ( 
.A(n_13248),
.B(n_2318),
.Y(n_13554)
);

OAI22xp33_ASAP7_75t_L g13555 ( 
.A1(n_13340),
.A2(n_2321),
.B1(n_2319),
.B2(n_2320),
.Y(n_13555)
);

INVx1_ASAP7_75t_L g13556 ( 
.A(n_13080),
.Y(n_13556)
);

AO21x2_ASAP7_75t_L g13557 ( 
.A1(n_13311),
.A2(n_2320),
.B(n_2321),
.Y(n_13557)
);

OAI211xp5_ASAP7_75t_SL g13558 ( 
.A1(n_13055),
.A2(n_2324),
.B(n_2322),
.C(n_2323),
.Y(n_13558)
);

AOI222xp33_ASAP7_75t_L g13559 ( 
.A1(n_13373),
.A2(n_2325),
.B1(n_2327),
.B2(n_2322),
.C1(n_2324),
.C2(n_2326),
.Y(n_13559)
);

INVx2_ASAP7_75t_L g13560 ( 
.A(n_13297),
.Y(n_13560)
);

AOI22xp33_ASAP7_75t_L g13561 ( 
.A1(n_13262),
.A2(n_2327),
.B1(n_2325),
.B2(n_2326),
.Y(n_13561)
);

AOI22xp33_ASAP7_75t_L g13562 ( 
.A1(n_13265),
.A2(n_2331),
.B1(n_2328),
.B2(n_2329),
.Y(n_13562)
);

AOI22xp33_ASAP7_75t_L g13563 ( 
.A1(n_13364),
.A2(n_2332),
.B1(n_2329),
.B2(n_2331),
.Y(n_13563)
);

AOI211xp5_ASAP7_75t_L g13564 ( 
.A1(n_13271),
.A2(n_2335),
.B(n_2333),
.C(n_2334),
.Y(n_13564)
);

INVx2_ASAP7_75t_L g13565 ( 
.A(n_13345),
.Y(n_13565)
);

AOI22xp33_ASAP7_75t_L g13566 ( 
.A1(n_13106),
.A2(n_2337),
.B1(n_2333),
.B2(n_2336),
.Y(n_13566)
);

INVx2_ASAP7_75t_L g13567 ( 
.A(n_13148),
.Y(n_13567)
);

OAI22xp5_ASAP7_75t_L g13568 ( 
.A1(n_13333),
.A2(n_2339),
.B1(n_2336),
.B2(n_2338),
.Y(n_13568)
);

AO21x2_ASAP7_75t_L g13569 ( 
.A1(n_13290),
.A2(n_2338),
.B(n_2339),
.Y(n_13569)
);

NAND2xp5_ASAP7_75t_L g13570 ( 
.A(n_13327),
.B(n_2340),
.Y(n_13570)
);

INVx1_ASAP7_75t_L g13571 ( 
.A(n_13081),
.Y(n_13571)
);

OAI22xp5_ASAP7_75t_L g13572 ( 
.A1(n_13076),
.A2(n_2342),
.B1(n_2340),
.B2(n_2341),
.Y(n_13572)
);

CKINVDCx20_ASAP7_75t_R g13573 ( 
.A(n_13310),
.Y(n_13573)
);

INVx1_ASAP7_75t_L g13574 ( 
.A(n_13083),
.Y(n_13574)
);

INVx2_ASAP7_75t_L g13575 ( 
.A(n_13057),
.Y(n_13575)
);

AOI22xp5_ASAP7_75t_SL g13576 ( 
.A1(n_13386),
.A2(n_2343),
.B1(n_2341),
.B2(n_2342),
.Y(n_13576)
);

A2O1A1Ixp33_ASAP7_75t_L g13577 ( 
.A1(n_13353),
.A2(n_2345),
.B(n_2343),
.C(n_2344),
.Y(n_13577)
);

AOI22xp33_ASAP7_75t_L g13578 ( 
.A1(n_13231),
.A2(n_2347),
.B1(n_2344),
.B2(n_2346),
.Y(n_13578)
);

INVx2_ASAP7_75t_L g13579 ( 
.A(n_13068),
.Y(n_13579)
);

OAI22xp33_ASAP7_75t_L g13580 ( 
.A1(n_13341),
.A2(n_2349),
.B1(n_2347),
.B2(n_2348),
.Y(n_13580)
);

AOI22xp33_ASAP7_75t_L g13581 ( 
.A1(n_13169),
.A2(n_2350),
.B1(n_2348),
.B2(n_2349),
.Y(n_13581)
);

AOI22xp33_ASAP7_75t_L g13582 ( 
.A1(n_13173),
.A2(n_2352),
.B1(n_2350),
.B2(n_2351),
.Y(n_13582)
);

INVx1_ASAP7_75t_L g13583 ( 
.A(n_13084),
.Y(n_13583)
);

AOI22xp33_ASAP7_75t_L g13584 ( 
.A1(n_13211),
.A2(n_13292),
.B1(n_13199),
.B2(n_13204),
.Y(n_13584)
);

AOI221xp5_ASAP7_75t_L g13585 ( 
.A1(n_13180),
.A2(n_2353),
.B1(n_2351),
.B2(n_2352),
.C(n_2354),
.Y(n_13585)
);

OAI221xp5_ASAP7_75t_L g13586 ( 
.A1(n_13206),
.A2(n_2355),
.B1(n_2353),
.B2(n_2354),
.C(n_2356),
.Y(n_13586)
);

BUFx6f_ASAP7_75t_L g13587 ( 
.A(n_13218),
.Y(n_13587)
);

AOI22xp5_ASAP7_75t_L g13588 ( 
.A1(n_13381),
.A2(n_2357),
.B1(n_2355),
.B2(n_2356),
.Y(n_13588)
);

INVx2_ASAP7_75t_L g13589 ( 
.A(n_13313),
.Y(n_13589)
);

AOI21xp5_ASAP7_75t_L g13590 ( 
.A1(n_13306),
.A2(n_13123),
.B(n_13338),
.Y(n_13590)
);

OAI22xp5_ASAP7_75t_L g13591 ( 
.A1(n_13347),
.A2(n_2359),
.B1(n_2357),
.B2(n_2358),
.Y(n_13591)
);

OR2x2_ASAP7_75t_L g13592 ( 
.A(n_13174),
.B(n_2358),
.Y(n_13592)
);

AOI211xp5_ASAP7_75t_L g13593 ( 
.A1(n_13227),
.A2(n_2361),
.B(n_2359),
.C(n_2360),
.Y(n_13593)
);

OAI22xp33_ASAP7_75t_L g13594 ( 
.A1(n_13269),
.A2(n_2363),
.B1(n_2360),
.B2(n_2362),
.Y(n_13594)
);

AOI22xp33_ASAP7_75t_L g13595 ( 
.A1(n_13238),
.A2(n_2366),
.B1(n_2362),
.B2(n_2365),
.Y(n_13595)
);

NOR2xp33_ASAP7_75t_L g13596 ( 
.A(n_13249),
.B(n_2366),
.Y(n_13596)
);

INVx2_ASAP7_75t_L g13597 ( 
.A(n_13330),
.Y(n_13597)
);

AND2x4_ASAP7_75t_L g13598 ( 
.A(n_13294),
.B(n_2367),
.Y(n_13598)
);

INVx8_ASAP7_75t_L g13599 ( 
.A(n_13136),
.Y(n_13599)
);

INVx2_ASAP7_75t_L g13600 ( 
.A(n_13334),
.Y(n_13600)
);

OAI22xp5_ASAP7_75t_L g13601 ( 
.A1(n_13221),
.A2(n_2369),
.B1(n_2367),
.B2(n_2368),
.Y(n_13601)
);

AOI21xp5_ASAP7_75t_L g13602 ( 
.A1(n_13296),
.A2(n_2369),
.B(n_2370),
.Y(n_13602)
);

AND2x2_ASAP7_75t_L g13603 ( 
.A(n_13059),
.B(n_2370),
.Y(n_13603)
);

OAI211xp5_ASAP7_75t_SL g13604 ( 
.A1(n_13375),
.A2(n_2374),
.B(n_2371),
.C(n_2372),
.Y(n_13604)
);

AND2x4_ASAP7_75t_L g13605 ( 
.A(n_13100),
.B(n_2371),
.Y(n_13605)
);

AND2x6_ASAP7_75t_L g13606 ( 
.A(n_13219),
.B(n_2372),
.Y(n_13606)
);

OAI22xp5_ASAP7_75t_L g13607 ( 
.A1(n_13195),
.A2(n_2377),
.B1(n_2375),
.B2(n_2376),
.Y(n_13607)
);

INVx4_ASAP7_75t_SL g13608 ( 
.A(n_13095),
.Y(n_13608)
);

NOR2xp33_ASAP7_75t_L g13609 ( 
.A(n_13159),
.B(n_2376),
.Y(n_13609)
);

INVxp67_ASAP7_75t_L g13610 ( 
.A(n_13368),
.Y(n_13610)
);

AOI22xp33_ASAP7_75t_SL g13611 ( 
.A1(n_13182),
.A2(n_2380),
.B1(n_2377),
.B2(n_2378),
.Y(n_13611)
);

OA21x2_ASAP7_75t_L g13612 ( 
.A1(n_13060),
.A2(n_2380),
.B(n_2381),
.Y(n_13612)
);

OA21x2_ASAP7_75t_L g13613 ( 
.A1(n_13064),
.A2(n_2381),
.B(n_2382),
.Y(n_13613)
);

AOI22xp33_ASAP7_75t_L g13614 ( 
.A1(n_13198),
.A2(n_2384),
.B1(n_2382),
.B2(n_2383),
.Y(n_13614)
);

OAI221xp5_ASAP7_75t_SL g13615 ( 
.A1(n_13348),
.A2(n_2386),
.B1(n_2384),
.B2(n_2385),
.C(n_2387),
.Y(n_13615)
);

INVx2_ASAP7_75t_L g13616 ( 
.A(n_13202),
.Y(n_13616)
);

OAI211xp5_ASAP7_75t_L g13617 ( 
.A1(n_13315),
.A2(n_2387),
.B(n_2385),
.C(n_2386),
.Y(n_13617)
);

OAI22xp5_ASAP7_75t_L g13618 ( 
.A1(n_13207),
.A2(n_13208),
.B1(n_13205),
.B2(n_13203),
.Y(n_13618)
);

AOI22xp33_ASAP7_75t_L g13619 ( 
.A1(n_13298),
.A2(n_2390),
.B1(n_2388),
.B2(n_2389),
.Y(n_13619)
);

AOI21xp5_ASAP7_75t_L g13620 ( 
.A1(n_13175),
.A2(n_2388),
.B(n_2389),
.Y(n_13620)
);

AOI22xp33_ASAP7_75t_L g13621 ( 
.A1(n_13093),
.A2(n_2393),
.B1(n_2391),
.B2(n_2392),
.Y(n_13621)
);

AOI221xp5_ASAP7_75t_L g13622 ( 
.A1(n_13192),
.A2(n_2394),
.B1(n_2392),
.B2(n_2393),
.C(n_2395),
.Y(n_13622)
);

NAND2xp5_ASAP7_75t_L g13623 ( 
.A(n_13116),
.B(n_2395),
.Y(n_13623)
);

CKINVDCx5p33_ASAP7_75t_R g13624 ( 
.A(n_13213),
.Y(n_13624)
);

AOI222xp33_ASAP7_75t_L g13625 ( 
.A1(n_13325),
.A2(n_2398),
.B1(n_2400),
.B2(n_2396),
.C1(n_2397),
.C2(n_2399),
.Y(n_13625)
);

AOI22xp33_ASAP7_75t_L g13626 ( 
.A1(n_13102),
.A2(n_2398),
.B1(n_2396),
.B2(n_2397),
.Y(n_13626)
);

INVx2_ASAP7_75t_L g13627 ( 
.A(n_13132),
.Y(n_13627)
);

NAND2xp5_ASAP7_75t_L g13628 ( 
.A(n_13118),
.B(n_2400),
.Y(n_13628)
);

INVx2_ASAP7_75t_L g13629 ( 
.A(n_13361),
.Y(n_13629)
);

INVx1_ASAP7_75t_SL g13630 ( 
.A(n_13276),
.Y(n_13630)
);

AND2x2_ASAP7_75t_SL g13631 ( 
.A(n_13050),
.B(n_2401),
.Y(n_13631)
);

OAI21xp5_ASAP7_75t_L g13632 ( 
.A1(n_13082),
.A2(n_2401),
.B(n_2402),
.Y(n_13632)
);

AOI222xp33_ASAP7_75t_L g13633 ( 
.A1(n_13228),
.A2(n_2404),
.B1(n_2406),
.B2(n_2402),
.C1(n_2403),
.C2(n_2405),
.Y(n_13633)
);

OAI22xp5_ASAP7_75t_L g13634 ( 
.A1(n_13073),
.A2(n_2406),
.B1(n_2404),
.B2(n_2405),
.Y(n_13634)
);

AOI221xp5_ASAP7_75t_L g13635 ( 
.A1(n_13233),
.A2(n_2409),
.B1(n_2407),
.B2(n_2408),
.C(n_2410),
.Y(n_13635)
);

AOI22xp33_ASAP7_75t_L g13636 ( 
.A1(n_13342),
.A2(n_13236),
.B1(n_13235),
.B2(n_13217),
.Y(n_13636)
);

AOI221xp5_ASAP7_75t_L g13637 ( 
.A1(n_13186),
.A2(n_2411),
.B1(n_2409),
.B2(n_2410),
.C(n_2412),
.Y(n_13637)
);

OAI322xp33_ASAP7_75t_L g13638 ( 
.A1(n_13216),
.A2(n_2416),
.A3(n_2415),
.B1(n_2413),
.B2(n_2411),
.C1(n_2412),
.C2(n_2414),
.Y(n_13638)
);

OAI21x1_ASAP7_75t_L g13639 ( 
.A1(n_13293),
.A2(n_13260),
.B(n_13066),
.Y(n_13639)
);

INVx3_ASAP7_75t_L g13640 ( 
.A(n_13063),
.Y(n_13640)
);

AND2x2_ASAP7_75t_L g13641 ( 
.A(n_13121),
.B(n_2413),
.Y(n_13641)
);

BUFx3_ASAP7_75t_L g13642 ( 
.A(n_13268),
.Y(n_13642)
);

AOI22xp33_ASAP7_75t_L g13643 ( 
.A1(n_13215),
.A2(n_2416),
.B1(n_2414),
.B2(n_2415),
.Y(n_13643)
);

AND2x2_ASAP7_75t_L g13644 ( 
.A(n_13115),
.B(n_2417),
.Y(n_13644)
);

OAI21x1_ASAP7_75t_L g13645 ( 
.A1(n_13331),
.A2(n_13332),
.B(n_13226),
.Y(n_13645)
);

AND2x2_ASAP7_75t_L g13646 ( 
.A(n_13074),
.B(n_2417),
.Y(n_13646)
);

AND2x2_ASAP7_75t_L g13647 ( 
.A(n_13409),
.B(n_13131),
.Y(n_13647)
);

NAND2xp5_ASAP7_75t_L g13648 ( 
.A(n_13630),
.B(n_13120),
.Y(n_13648)
);

OR2x2_ASAP7_75t_L g13649 ( 
.A(n_13414),
.B(n_13135),
.Y(n_13649)
);

INVx2_ASAP7_75t_L g13650 ( 
.A(n_13393),
.Y(n_13650)
);

NOR2xp33_ASAP7_75t_L g13651 ( 
.A(n_13396),
.B(n_13351),
.Y(n_13651)
);

NAND2xp5_ASAP7_75t_L g13652 ( 
.A(n_13609),
.B(n_13133),
.Y(n_13652)
);

INVxp67_ASAP7_75t_L g13653 ( 
.A(n_13423),
.Y(n_13653)
);

BUFx3_ASAP7_75t_L g13654 ( 
.A(n_13447),
.Y(n_13654)
);

AND2x2_ASAP7_75t_L g13655 ( 
.A(n_13449),
.B(n_13141),
.Y(n_13655)
);

INVx1_ASAP7_75t_L g13656 ( 
.A(n_13431),
.Y(n_13656)
);

NAND2xp5_ASAP7_75t_L g13657 ( 
.A(n_13418),
.B(n_13459),
.Y(n_13657)
);

OR2x2_ASAP7_75t_L g13658 ( 
.A(n_13417),
.B(n_13144),
.Y(n_13658)
);

INVx3_ASAP7_75t_L g13659 ( 
.A(n_13468),
.Y(n_13659)
);

AND2x2_ASAP7_75t_L g13660 ( 
.A(n_13502),
.B(n_13543),
.Y(n_13660)
);

NOR2x1_ASAP7_75t_R g13661 ( 
.A(n_13473),
.B(n_13252),
.Y(n_13661)
);

AND2x2_ASAP7_75t_L g13662 ( 
.A(n_13528),
.B(n_13087),
.Y(n_13662)
);

INVx2_ASAP7_75t_L g13663 ( 
.A(n_13587),
.Y(n_13663)
);

OR2x2_ASAP7_75t_L g13664 ( 
.A(n_13421),
.B(n_13210),
.Y(n_13664)
);

HB1xp67_ASAP7_75t_L g13665 ( 
.A(n_13399),
.Y(n_13665)
);

OR2x2_ASAP7_75t_L g13666 ( 
.A(n_13567),
.B(n_13295),
.Y(n_13666)
);

BUFx2_ASAP7_75t_L g13667 ( 
.A(n_13573),
.Y(n_13667)
);

INVx2_ASAP7_75t_L g13668 ( 
.A(n_13587),
.Y(n_13668)
);

INVx3_ASAP7_75t_L g13669 ( 
.A(n_13468),
.Y(n_13669)
);

AOI222xp33_ASAP7_75t_L g13670 ( 
.A1(n_13542),
.A2(n_13299),
.B1(n_13274),
.B2(n_13304),
.C1(n_13301),
.C2(n_13300),
.Y(n_13670)
);

INVx1_ASAP7_75t_L g13671 ( 
.A(n_13431),
.Y(n_13671)
);

INVx2_ASAP7_75t_L g13672 ( 
.A(n_13642),
.Y(n_13672)
);

INVx1_ASAP7_75t_L g13673 ( 
.A(n_13442),
.Y(n_13673)
);

AND2x2_ASAP7_75t_L g13674 ( 
.A(n_13537),
.B(n_13090),
.Y(n_13674)
);

BUFx6f_ASAP7_75t_L g13675 ( 
.A(n_13524),
.Y(n_13675)
);

NAND2xp5_ASAP7_75t_L g13676 ( 
.A(n_13590),
.B(n_13155),
.Y(n_13676)
);

CKINVDCx11_ASAP7_75t_R g13677 ( 
.A(n_13488),
.Y(n_13677)
);

NAND2xp5_ASAP7_75t_L g13678 ( 
.A(n_13406),
.B(n_13321),
.Y(n_13678)
);

INVx1_ASAP7_75t_L g13679 ( 
.A(n_13486),
.Y(n_13679)
);

AND2x2_ASAP7_75t_L g13680 ( 
.A(n_13501),
.B(n_13092),
.Y(n_13680)
);

AND2x2_ASAP7_75t_L g13681 ( 
.A(n_13527),
.B(n_13510),
.Y(n_13681)
);

HB1xp67_ASAP7_75t_L g13682 ( 
.A(n_13432),
.Y(n_13682)
);

INVx2_ASAP7_75t_L g13683 ( 
.A(n_13547),
.Y(n_13683)
);

OR2x2_ASAP7_75t_L g13684 ( 
.A(n_13533),
.B(n_13335),
.Y(n_13684)
);

AND2x2_ASAP7_75t_L g13685 ( 
.A(n_13560),
.B(n_13138),
.Y(n_13685)
);

INVx2_ASAP7_75t_SL g13686 ( 
.A(n_13599),
.Y(n_13686)
);

BUFx2_ASAP7_75t_L g13687 ( 
.A(n_13624),
.Y(n_13687)
);

NAND2xp5_ASAP7_75t_L g13688 ( 
.A(n_13602),
.B(n_13326),
.Y(n_13688)
);

INVx3_ASAP7_75t_L g13689 ( 
.A(n_13599),
.Y(n_13689)
);

OR2x2_ASAP7_75t_L g13690 ( 
.A(n_13506),
.B(n_13339),
.Y(n_13690)
);

INVx2_ASAP7_75t_L g13691 ( 
.A(n_13547),
.Y(n_13691)
);

INVx3_ASAP7_75t_SL g13692 ( 
.A(n_13498),
.Y(n_13692)
);

INVx1_ASAP7_75t_L g13693 ( 
.A(n_13457),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_13429),
.Y(n_13694)
);

OR2x2_ASAP7_75t_L g13695 ( 
.A(n_13526),
.B(n_13323),
.Y(n_13695)
);

AND2x2_ASAP7_75t_L g13696 ( 
.A(n_13523),
.B(n_13337),
.Y(n_13696)
);

INVx2_ASAP7_75t_L g13697 ( 
.A(n_13461),
.Y(n_13697)
);

INVx2_ASAP7_75t_L g13698 ( 
.A(n_13461),
.Y(n_13698)
);

AND2x4_ASAP7_75t_L g13699 ( 
.A(n_13608),
.B(n_13234),
.Y(n_13699)
);

INVx2_ASAP7_75t_L g13700 ( 
.A(n_13487),
.Y(n_13700)
);

AND2x2_ASAP7_75t_L g13701 ( 
.A(n_13565),
.B(n_13185),
.Y(n_13701)
);

INVx2_ASAP7_75t_L g13702 ( 
.A(n_13487),
.Y(n_13702)
);

BUFx3_ASAP7_75t_L g13703 ( 
.A(n_13606),
.Y(n_13703)
);

INVx1_ASAP7_75t_L g13704 ( 
.A(n_13570),
.Y(n_13704)
);

INVx3_ASAP7_75t_L g13705 ( 
.A(n_13402),
.Y(n_13705)
);

INVx2_ASAP7_75t_L g13706 ( 
.A(n_13487),
.Y(n_13706)
);

HB1xp67_ASAP7_75t_L g13707 ( 
.A(n_13610),
.Y(n_13707)
);

INVx1_ASAP7_75t_L g13708 ( 
.A(n_13416),
.Y(n_13708)
);

INVx2_ASAP7_75t_L g13709 ( 
.A(n_13487),
.Y(n_13709)
);

INVx2_ASAP7_75t_L g13710 ( 
.A(n_13605),
.Y(n_13710)
);

INVx1_ASAP7_75t_L g13711 ( 
.A(n_13438),
.Y(n_13711)
);

INVx2_ASAP7_75t_L g13712 ( 
.A(n_13631),
.Y(n_13712)
);

BUFx6f_ASAP7_75t_L g13713 ( 
.A(n_13517),
.Y(n_13713)
);

INVx2_ASAP7_75t_L g13714 ( 
.A(n_13608),
.Y(n_13714)
);

AND2x2_ASAP7_75t_L g13715 ( 
.A(n_13444),
.B(n_13266),
.Y(n_13715)
);

BUFx2_ASAP7_75t_L g13716 ( 
.A(n_13403),
.Y(n_13716)
);

AND2x4_ASAP7_75t_L g13717 ( 
.A(n_13640),
.B(n_13229),
.Y(n_13717)
);

INVx1_ASAP7_75t_L g13718 ( 
.A(n_13427),
.Y(n_13718)
);

INVx1_ASAP7_75t_L g13719 ( 
.A(n_13452),
.Y(n_13719)
);

OAI22xp5_ASAP7_75t_SL g13720 ( 
.A1(n_13434),
.A2(n_13254),
.B1(n_13191),
.B2(n_13279),
.Y(n_13720)
);

INVx3_ASAP7_75t_L g13721 ( 
.A(n_13451),
.Y(n_13721)
);

NAND2xp5_ASAP7_75t_L g13722 ( 
.A(n_13549),
.B(n_13352),
.Y(n_13722)
);

INVx2_ASAP7_75t_SL g13723 ( 
.A(n_13435),
.Y(n_13723)
);

INVx1_ASAP7_75t_L g13724 ( 
.A(n_13455),
.Y(n_13724)
);

CKINVDCx20_ASAP7_75t_R g13725 ( 
.A(n_13408),
.Y(n_13725)
);

AND2x4_ASAP7_75t_SL g13726 ( 
.A(n_13598),
.B(n_13282),
.Y(n_13726)
);

INVxp67_ASAP7_75t_SL g13727 ( 
.A(n_13464),
.Y(n_13727)
);

AND2x2_ASAP7_75t_L g13728 ( 
.A(n_13546),
.B(n_13134),
.Y(n_13728)
);

INVx3_ASAP7_75t_L g13729 ( 
.A(n_13493),
.Y(n_13729)
);

AND2x2_ASAP7_75t_L g13730 ( 
.A(n_13554),
.B(n_13126),
.Y(n_13730)
);

NAND2xp5_ASAP7_75t_L g13731 ( 
.A(n_13551),
.B(n_13354),
.Y(n_13731)
);

AND2x2_ASAP7_75t_L g13732 ( 
.A(n_13641),
.B(n_13105),
.Y(n_13732)
);

HB1xp67_ASAP7_75t_L g13733 ( 
.A(n_13600),
.Y(n_13733)
);

HB1xp67_ASAP7_75t_L g13734 ( 
.A(n_13467),
.Y(n_13734)
);

BUFx3_ASAP7_75t_L g13735 ( 
.A(n_13606),
.Y(n_13735)
);

NAND2xp5_ASAP7_75t_L g13736 ( 
.A(n_13541),
.B(n_13329),
.Y(n_13736)
);

OR2x2_ASAP7_75t_L g13737 ( 
.A(n_13426),
.B(n_13362),
.Y(n_13737)
);

INVx3_ASAP7_75t_L g13738 ( 
.A(n_13603),
.Y(n_13738)
);

INVx2_ASAP7_75t_L g13739 ( 
.A(n_13492),
.Y(n_13739)
);

BUFx3_ASAP7_75t_L g13740 ( 
.A(n_13606),
.Y(n_13740)
);

NOR2xp33_ASAP7_75t_L g13741 ( 
.A(n_13552),
.B(n_13179),
.Y(n_13741)
);

AND2x2_ASAP7_75t_L g13742 ( 
.A(n_13496),
.B(n_13596),
.Y(n_13742)
);

INVx1_ASAP7_75t_L g13743 ( 
.A(n_13460),
.Y(n_13743)
);

INVx2_ASAP7_75t_L g13744 ( 
.A(n_13612),
.Y(n_13744)
);

INVx2_ASAP7_75t_L g13745 ( 
.A(n_13613),
.Y(n_13745)
);

INVx2_ASAP7_75t_L g13746 ( 
.A(n_13482),
.Y(n_13746)
);

INVx2_ASAP7_75t_L g13747 ( 
.A(n_13557),
.Y(n_13747)
);

AND2x2_ASAP7_75t_L g13748 ( 
.A(n_13512),
.B(n_13232),
.Y(n_13748)
);

AND2x2_ASAP7_75t_L g13749 ( 
.A(n_13481),
.B(n_13317),
.Y(n_13749)
);

AND2x2_ASAP7_75t_L g13750 ( 
.A(n_13477),
.B(n_13322),
.Y(n_13750)
);

AND2x2_ASAP7_75t_L g13751 ( 
.A(n_13465),
.B(n_13308),
.Y(n_13751)
);

OR2x2_ASAP7_75t_L g13752 ( 
.A(n_13618),
.B(n_13309),
.Y(n_13752)
);

INVx1_ASAP7_75t_L g13753 ( 
.A(n_13519),
.Y(n_13753)
);

HB1xp67_ASAP7_75t_L g13754 ( 
.A(n_13645),
.Y(n_13754)
);

HB1xp67_ASAP7_75t_L g13755 ( 
.A(n_13410),
.Y(n_13755)
);

INVx1_ASAP7_75t_L g13756 ( 
.A(n_13425),
.Y(n_13756)
);

AND2x2_ASAP7_75t_L g13757 ( 
.A(n_13463),
.B(n_13314),
.Y(n_13757)
);

AND2x2_ASAP7_75t_L g13758 ( 
.A(n_13644),
.B(n_13382),
.Y(n_13758)
);

AND2x2_ASAP7_75t_L g13759 ( 
.A(n_13646),
.B(n_13062),
.Y(n_13759)
);

INVx3_ASAP7_75t_L g13760 ( 
.A(n_13419),
.Y(n_13760)
);

AND2x2_ASAP7_75t_L g13761 ( 
.A(n_13462),
.B(n_13372),
.Y(n_13761)
);

INVx1_ASAP7_75t_L g13762 ( 
.A(n_13469),
.Y(n_13762)
);

AND2x2_ASAP7_75t_L g13763 ( 
.A(n_13507),
.B(n_13224),
.Y(n_13763)
);

AND2x2_ASAP7_75t_L g13764 ( 
.A(n_13508),
.B(n_13193),
.Y(n_13764)
);

BUFx2_ASAP7_75t_L g13765 ( 
.A(n_13632),
.Y(n_13765)
);

BUFx12f_ASAP7_75t_L g13766 ( 
.A(n_13592),
.Y(n_13766)
);

INVx1_ASAP7_75t_L g13767 ( 
.A(n_13483),
.Y(n_13767)
);

INVx1_ASAP7_75t_L g13768 ( 
.A(n_13511),
.Y(n_13768)
);

BUFx2_ASAP7_75t_L g13769 ( 
.A(n_13577),
.Y(n_13769)
);

INVx2_ASAP7_75t_L g13770 ( 
.A(n_13471),
.Y(n_13770)
);

AND2x2_ASAP7_75t_L g13771 ( 
.A(n_13532),
.B(n_13139),
.Y(n_13771)
);

AND2x2_ASAP7_75t_L g13772 ( 
.A(n_13548),
.B(n_13245),
.Y(n_13772)
);

NAND2xp5_ASAP7_75t_L g13773 ( 
.A(n_13489),
.B(n_13197),
.Y(n_13773)
);

AND2x2_ASAP7_75t_L g13774 ( 
.A(n_13553),
.B(n_13270),
.Y(n_13774)
);

NAND2xp5_ASAP7_75t_L g13775 ( 
.A(n_13538),
.B(n_13355),
.Y(n_13775)
);

INVx2_ASAP7_75t_L g13776 ( 
.A(n_13569),
.Y(n_13776)
);

AND2x2_ASAP7_75t_L g13777 ( 
.A(n_13556),
.B(n_13078),
.Y(n_13777)
);

INVx1_ASAP7_75t_L g13778 ( 
.A(n_13571),
.Y(n_13778)
);

NAND2xp5_ASAP7_75t_L g13779 ( 
.A(n_13478),
.B(n_2418),
.Y(n_13779)
);

HB1xp67_ASAP7_75t_L g13780 ( 
.A(n_13629),
.Y(n_13780)
);

AOI22xp33_ASAP7_75t_L g13781 ( 
.A1(n_13589),
.A2(n_2420),
.B1(n_2418),
.B2(n_2419),
.Y(n_13781)
);

INVx2_ASAP7_75t_L g13782 ( 
.A(n_13412),
.Y(n_13782)
);

INVx2_ASAP7_75t_L g13783 ( 
.A(n_13401),
.Y(n_13783)
);

INVx2_ASAP7_75t_SL g13784 ( 
.A(n_13576),
.Y(n_13784)
);

INVx3_ASAP7_75t_SL g13785 ( 
.A(n_13575),
.Y(n_13785)
);

AND2x2_ASAP7_75t_L g13786 ( 
.A(n_13574),
.B(n_2420),
.Y(n_13786)
);

AND2x2_ASAP7_75t_L g13787 ( 
.A(n_13583),
.B(n_2421),
.Y(n_13787)
);

AND2x2_ASAP7_75t_L g13788 ( 
.A(n_13536),
.B(n_13520),
.Y(n_13788)
);

OR2x2_ASAP7_75t_L g13789 ( 
.A(n_13514),
.B(n_2422),
.Y(n_13789)
);

INVx2_ASAP7_75t_L g13790 ( 
.A(n_13504),
.Y(n_13790)
);

INVx1_ASAP7_75t_L g13791 ( 
.A(n_13623),
.Y(n_13791)
);

INVx2_ASAP7_75t_SL g13792 ( 
.A(n_13474),
.Y(n_13792)
);

AND2x2_ASAP7_75t_L g13793 ( 
.A(n_13490),
.B(n_2422),
.Y(n_13793)
);

AND2x2_ASAP7_75t_L g13794 ( 
.A(n_13430),
.B(n_2423),
.Y(n_13794)
);

INVx4_ASAP7_75t_L g13795 ( 
.A(n_13579),
.Y(n_13795)
);

AND2x2_ASAP7_75t_L g13796 ( 
.A(n_13389),
.B(n_13525),
.Y(n_13796)
);

INVxp67_ASAP7_75t_SL g13797 ( 
.A(n_13494),
.Y(n_13797)
);

NAND2xp5_ASAP7_75t_L g13798 ( 
.A(n_13441),
.B(n_2423),
.Y(n_13798)
);

OR2x2_ASAP7_75t_L g13799 ( 
.A(n_13568),
.B(n_13509),
.Y(n_13799)
);

INVx2_ASAP7_75t_L g13800 ( 
.A(n_13513),
.Y(n_13800)
);

INVx2_ASAP7_75t_L g13801 ( 
.A(n_13627),
.Y(n_13801)
);

AND2x2_ASAP7_75t_L g13802 ( 
.A(n_13394),
.B(n_2424),
.Y(n_13802)
);

INVx2_ASAP7_75t_L g13803 ( 
.A(n_13597),
.Y(n_13803)
);

AND2x2_ASAP7_75t_L g13804 ( 
.A(n_13529),
.B(n_2424),
.Y(n_13804)
);

INVx1_ASAP7_75t_L g13805 ( 
.A(n_13628),
.Y(n_13805)
);

INVx2_ASAP7_75t_L g13806 ( 
.A(n_13616),
.Y(n_13806)
);

AND2x2_ASAP7_75t_L g13807 ( 
.A(n_13397),
.B(n_2426),
.Y(n_13807)
);

AND2x2_ASAP7_75t_L g13808 ( 
.A(n_13499),
.B(n_2426),
.Y(n_13808)
);

NAND2xp5_ASAP7_75t_L g13809 ( 
.A(n_13415),
.B(n_2427),
.Y(n_13809)
);

INVx2_ASAP7_75t_L g13810 ( 
.A(n_13639),
.Y(n_13810)
);

AND2x2_ASAP7_75t_L g13811 ( 
.A(n_13530),
.B(n_2427),
.Y(n_13811)
);

HB1xp67_ASAP7_75t_L g13812 ( 
.A(n_13634),
.Y(n_13812)
);

CKINVDCx8_ASAP7_75t_R g13813 ( 
.A(n_13450),
.Y(n_13813)
);

AND2x2_ASAP7_75t_L g13814 ( 
.A(n_13611),
.B(n_2428),
.Y(n_13814)
);

INVx2_ASAP7_75t_L g13815 ( 
.A(n_13445),
.Y(n_13815)
);

AND2x2_ASAP7_75t_L g13816 ( 
.A(n_13456),
.B(n_2428),
.Y(n_13816)
);

AND2x4_ASAP7_75t_L g13817 ( 
.A(n_13454),
.B(n_2429),
.Y(n_13817)
);

INVx1_ASAP7_75t_L g13818 ( 
.A(n_13607),
.Y(n_13818)
);

AND2x4_ASAP7_75t_SL g13819 ( 
.A(n_13424),
.B(n_2429),
.Y(n_13819)
);

INVx2_ASAP7_75t_L g13820 ( 
.A(n_13550),
.Y(n_13820)
);

INVx1_ASAP7_75t_L g13821 ( 
.A(n_13601),
.Y(n_13821)
);

HB1xp67_ASAP7_75t_L g13822 ( 
.A(n_13420),
.Y(n_13822)
);

AND2x2_ASAP7_75t_L g13823 ( 
.A(n_13422),
.B(n_2430),
.Y(n_13823)
);

INVx2_ASAP7_75t_L g13824 ( 
.A(n_13407),
.Y(n_13824)
);

AND2x4_ASAP7_75t_SL g13825 ( 
.A(n_13539),
.B(n_2430),
.Y(n_13825)
);

OR2x2_ASAP7_75t_L g13826 ( 
.A(n_13485),
.B(n_2431),
.Y(n_13826)
);

INVxp67_ASAP7_75t_SL g13827 ( 
.A(n_13428),
.Y(n_13827)
);

HB1xp67_ASAP7_75t_L g13828 ( 
.A(n_13491),
.Y(n_13828)
);

INVx2_ASAP7_75t_L g13829 ( 
.A(n_13588),
.Y(n_13829)
);

AND2x2_ASAP7_75t_L g13830 ( 
.A(n_13625),
.B(n_2432),
.Y(n_13830)
);

BUFx2_ASAP7_75t_L g13831 ( 
.A(n_13411),
.Y(n_13831)
);

BUFx6f_ASAP7_75t_L g13832 ( 
.A(n_13535),
.Y(n_13832)
);

INVx2_ASAP7_75t_L g13833 ( 
.A(n_13448),
.Y(n_13833)
);

INVx2_ASAP7_75t_L g13834 ( 
.A(n_13503),
.Y(n_13834)
);

AND2x2_ASAP7_75t_L g13835 ( 
.A(n_13458),
.B(n_2432),
.Y(n_13835)
);

INVx1_ASAP7_75t_L g13836 ( 
.A(n_13436),
.Y(n_13836)
);

OAI22xp5_ASAP7_75t_L g13837 ( 
.A1(n_13584),
.A2(n_2437),
.B1(n_2433),
.B2(n_2435),
.Y(n_13837)
);

OR2x2_ASAP7_75t_L g13838 ( 
.A(n_13540),
.B(n_2433),
.Y(n_13838)
);

OR2x2_ASAP7_75t_L g13839 ( 
.A(n_13617),
.B(n_2435),
.Y(n_13839)
);

AND2x2_ASAP7_75t_L g13840 ( 
.A(n_13559),
.B(n_2437),
.Y(n_13840)
);

INVx1_ASAP7_75t_L g13841 ( 
.A(n_13591),
.Y(n_13841)
);

INVx2_ASAP7_75t_L g13842 ( 
.A(n_13500),
.Y(n_13842)
);

INVx1_ASAP7_75t_L g13843 ( 
.A(n_13545),
.Y(n_13843)
);

INVx1_ASAP7_75t_L g13844 ( 
.A(n_13475),
.Y(n_13844)
);

AND2x4_ASAP7_75t_L g13845 ( 
.A(n_13484),
.B(n_2438),
.Y(n_13845)
);

INVx1_ASAP7_75t_L g13846 ( 
.A(n_13594),
.Y(n_13846)
);

AND2x4_ASAP7_75t_L g13847 ( 
.A(n_13405),
.B(n_2438),
.Y(n_13847)
);

NAND2xp5_ASAP7_75t_L g13848 ( 
.A(n_13440),
.B(n_2439),
.Y(n_13848)
);

BUFx3_ASAP7_75t_L g13849 ( 
.A(n_13453),
.Y(n_13849)
);

INVx1_ASAP7_75t_L g13850 ( 
.A(n_13667),
.Y(n_13850)
);

NAND2xp5_ASAP7_75t_L g13851 ( 
.A(n_13738),
.B(n_13413),
.Y(n_13851)
);

INVx1_ASAP7_75t_L g13852 ( 
.A(n_13780),
.Y(n_13852)
);

INVx1_ASAP7_75t_L g13853 ( 
.A(n_13707),
.Y(n_13853)
);

INVx2_ASAP7_75t_L g13854 ( 
.A(n_13677),
.Y(n_13854)
);

OR2x6_ASAP7_75t_SL g13855 ( 
.A(n_13683),
.B(n_13572),
.Y(n_13855)
);

AND2x2_ASAP7_75t_L g13856 ( 
.A(n_13654),
.B(n_13497),
.Y(n_13856)
);

INVx1_ASAP7_75t_L g13857 ( 
.A(n_13665),
.Y(n_13857)
);

AND2x2_ASAP7_75t_L g13858 ( 
.A(n_13716),
.B(n_13563),
.Y(n_13858)
);

INVx2_ASAP7_75t_L g13859 ( 
.A(n_13725),
.Y(n_13859)
);

INVx2_ASAP7_75t_L g13860 ( 
.A(n_13713),
.Y(n_13860)
);

BUFx2_ASAP7_75t_L g13861 ( 
.A(n_13661),
.Y(n_13861)
);

INVx2_ASAP7_75t_L g13862 ( 
.A(n_13713),
.Y(n_13862)
);

INVx1_ASAP7_75t_L g13863 ( 
.A(n_13682),
.Y(n_13863)
);

INVx1_ASAP7_75t_L g13864 ( 
.A(n_13734),
.Y(n_13864)
);

OR2x2_ASAP7_75t_L g13865 ( 
.A(n_13649),
.B(n_13615),
.Y(n_13865)
);

OR2x2_ASAP7_75t_L g13866 ( 
.A(n_13708),
.B(n_13505),
.Y(n_13866)
);

AND2x2_ASAP7_75t_L g13867 ( 
.A(n_13692),
.B(n_13398),
.Y(n_13867)
);

INVx1_ASAP7_75t_L g13868 ( 
.A(n_13656),
.Y(n_13868)
);

NAND2xp5_ASAP7_75t_L g13869 ( 
.A(n_13739),
.B(n_13620),
.Y(n_13869)
);

INVx1_ASAP7_75t_L g13870 ( 
.A(n_13671),
.Y(n_13870)
);

AND2x2_ASAP7_75t_L g13871 ( 
.A(n_13660),
.B(n_13495),
.Y(n_13871)
);

AND2x4_ASAP7_75t_L g13872 ( 
.A(n_13699),
.B(n_13687),
.Y(n_13872)
);

AND2x4_ASAP7_75t_L g13873 ( 
.A(n_13715),
.B(n_13433),
.Y(n_13873)
);

INVx1_ASAP7_75t_L g13874 ( 
.A(n_13693),
.Y(n_13874)
);

INVx1_ASAP7_75t_L g13875 ( 
.A(n_13673),
.Y(n_13875)
);

INVx1_ASAP7_75t_L g13876 ( 
.A(n_13679),
.Y(n_13876)
);

NOR2xp33_ASAP7_75t_L g13877 ( 
.A(n_13653),
.B(n_13443),
.Y(n_13877)
);

AND2x2_ASAP7_75t_L g13878 ( 
.A(n_13721),
.B(n_13659),
.Y(n_13878)
);

OR2x2_ASAP7_75t_L g13879 ( 
.A(n_13711),
.B(n_13580),
.Y(n_13879)
);

INVx1_ASAP7_75t_L g13880 ( 
.A(n_13753),
.Y(n_13880)
);

INVx1_ASAP7_75t_L g13881 ( 
.A(n_13757),
.Y(n_13881)
);

OR2x2_ASAP7_75t_L g13882 ( 
.A(n_13666),
.B(n_13695),
.Y(n_13882)
);

INVx2_ASAP7_75t_L g13883 ( 
.A(n_13675),
.Y(n_13883)
);

INVx1_ASAP7_75t_L g13884 ( 
.A(n_13786),
.Y(n_13884)
);

AND2x2_ASAP7_75t_L g13885 ( 
.A(n_13669),
.B(n_13392),
.Y(n_13885)
);

AND2x2_ASAP7_75t_L g13886 ( 
.A(n_13689),
.B(n_13390),
.Y(n_13886)
);

NAND2xp5_ASAP7_75t_L g13887 ( 
.A(n_13758),
.B(n_13476),
.Y(n_13887)
);

OR2x2_ASAP7_75t_L g13888 ( 
.A(n_13650),
.B(n_13521),
.Y(n_13888)
);

INVx3_ASAP7_75t_L g13889 ( 
.A(n_13717),
.Y(n_13889)
);

BUFx2_ASAP7_75t_L g13890 ( 
.A(n_13714),
.Y(n_13890)
);

AOI22xp33_ASAP7_75t_L g13891 ( 
.A1(n_13829),
.A2(n_13636),
.B1(n_13604),
.B2(n_13391),
.Y(n_13891)
);

INVx1_ASAP7_75t_L g13892 ( 
.A(n_13787),
.Y(n_13892)
);

INVx1_ASAP7_75t_L g13893 ( 
.A(n_13664),
.Y(n_13893)
);

OR2x2_ASAP7_75t_L g13894 ( 
.A(n_13657),
.B(n_13446),
.Y(n_13894)
);

INVx1_ASAP7_75t_L g13895 ( 
.A(n_13658),
.Y(n_13895)
);

OR2x2_ASAP7_75t_L g13896 ( 
.A(n_13672),
.B(n_13470),
.Y(n_13896)
);

INVx1_ASAP7_75t_L g13897 ( 
.A(n_13746),
.Y(n_13897)
);

OR2x2_ASAP7_75t_L g13898 ( 
.A(n_13690),
.B(n_13555),
.Y(n_13898)
);

INVx1_ASAP7_75t_L g13899 ( 
.A(n_13835),
.Y(n_13899)
);

INVx1_ASAP7_75t_L g13900 ( 
.A(n_13694),
.Y(n_13900)
);

BUFx2_ASAP7_75t_L g13901 ( 
.A(n_13705),
.Y(n_13901)
);

INVx1_ASAP7_75t_L g13902 ( 
.A(n_13674),
.Y(n_13902)
);

AND2x2_ASAP7_75t_L g13903 ( 
.A(n_13681),
.B(n_13593),
.Y(n_13903)
);

NAND2xp5_ASAP7_75t_L g13904 ( 
.A(n_13830),
.B(n_13534),
.Y(n_13904)
);

INVx2_ASAP7_75t_L g13905 ( 
.A(n_13675),
.Y(n_13905)
);

INVx2_ASAP7_75t_L g13906 ( 
.A(n_13703),
.Y(n_13906)
);

INVx2_ASAP7_75t_L g13907 ( 
.A(n_13735),
.Y(n_13907)
);

INVx2_ASAP7_75t_L g13908 ( 
.A(n_13740),
.Y(n_13908)
);

AND2x2_ASAP7_75t_L g13909 ( 
.A(n_13655),
.B(n_13564),
.Y(n_13909)
);

INVx1_ASAP7_75t_L g13910 ( 
.A(n_13801),
.Y(n_13910)
);

AND2x2_ASAP7_75t_L g13911 ( 
.A(n_13701),
.B(n_13633),
.Y(n_13911)
);

INVx2_ASAP7_75t_L g13912 ( 
.A(n_13732),
.Y(n_13912)
);

AND2x4_ASAP7_75t_L g13913 ( 
.A(n_13723),
.B(n_13518),
.Y(n_13913)
);

AND2x2_ASAP7_75t_L g13914 ( 
.A(n_13686),
.B(n_13531),
.Y(n_13914)
);

BUFx3_ASAP7_75t_L g13915 ( 
.A(n_13766),
.Y(n_13915)
);

OR2x2_ASAP7_75t_L g13916 ( 
.A(n_13684),
.B(n_13400),
.Y(n_13916)
);

INVx1_ASAP7_75t_L g13917 ( 
.A(n_13803),
.Y(n_13917)
);

AND2x2_ASAP7_75t_L g13918 ( 
.A(n_13647),
.B(n_13395),
.Y(n_13918)
);

INVx2_ASAP7_75t_L g13919 ( 
.A(n_13712),
.Y(n_13919)
);

HB1xp67_ASAP7_75t_L g13920 ( 
.A(n_13697),
.Y(n_13920)
);

INVx1_ASAP7_75t_L g13921 ( 
.A(n_13806),
.Y(n_13921)
);

AND2x2_ASAP7_75t_L g13922 ( 
.A(n_13691),
.B(n_13566),
.Y(n_13922)
);

NAND2xp5_ASAP7_75t_L g13923 ( 
.A(n_13797),
.B(n_13522),
.Y(n_13923)
);

INVx2_ASAP7_75t_L g13924 ( 
.A(n_13726),
.Y(n_13924)
);

INVx2_ASAP7_75t_L g13925 ( 
.A(n_13685),
.Y(n_13925)
);

INVx1_ASAP7_75t_L g13926 ( 
.A(n_13718),
.Y(n_13926)
);

INVx1_ASAP7_75t_L g13927 ( 
.A(n_13719),
.Y(n_13927)
);

AND2x2_ASAP7_75t_L g13928 ( 
.A(n_13662),
.B(n_13439),
.Y(n_13928)
);

INVx2_ASAP7_75t_L g13929 ( 
.A(n_13729),
.Y(n_13929)
);

AND2x2_ASAP7_75t_L g13930 ( 
.A(n_13651),
.B(n_13696),
.Y(n_13930)
);

INVx1_ASAP7_75t_L g13931 ( 
.A(n_13724),
.Y(n_13931)
);

INVx2_ASAP7_75t_L g13932 ( 
.A(n_13759),
.Y(n_13932)
);

AND2x2_ASAP7_75t_L g13933 ( 
.A(n_13663),
.B(n_13585),
.Y(n_13933)
);

NAND2x1p5_ASAP7_75t_L g13934 ( 
.A(n_13793),
.B(n_13466),
.Y(n_13934)
);

HB1xp67_ASAP7_75t_L g13935 ( 
.A(n_13698),
.Y(n_13935)
);

INVx1_ASAP7_75t_L g13936 ( 
.A(n_13743),
.Y(n_13936)
);

INVx1_ASAP7_75t_L g13937 ( 
.A(n_13756),
.Y(n_13937)
);

INVx2_ASAP7_75t_L g13938 ( 
.A(n_13742),
.Y(n_13938)
);

NAND2xp5_ASAP7_75t_L g13939 ( 
.A(n_13755),
.B(n_13622),
.Y(n_13939)
);

OR2x2_ASAP7_75t_L g13940 ( 
.A(n_13792),
.B(n_13648),
.Y(n_13940)
);

INVx1_ASAP7_75t_L g13941 ( 
.A(n_13762),
.Y(n_13941)
);

INVx2_ASAP7_75t_L g13942 ( 
.A(n_13737),
.Y(n_13942)
);

AND2x2_ASAP7_75t_L g13943 ( 
.A(n_13668),
.B(n_13578),
.Y(n_13943)
);

INVx2_ASAP7_75t_L g13944 ( 
.A(n_13760),
.Y(n_13944)
);

AND2x2_ASAP7_75t_L g13945 ( 
.A(n_13680),
.B(n_13621),
.Y(n_13945)
);

OR2x2_ASAP7_75t_L g13946 ( 
.A(n_13733),
.B(n_13472),
.Y(n_13946)
);

INVx1_ASAP7_75t_L g13947 ( 
.A(n_13767),
.Y(n_13947)
);

BUFx2_ASAP7_75t_L g13948 ( 
.A(n_13727),
.Y(n_13948)
);

INVx1_ASAP7_75t_L g13949 ( 
.A(n_13768),
.Y(n_13949)
);

AND2x2_ASAP7_75t_L g13950 ( 
.A(n_13788),
.B(n_13626),
.Y(n_13950)
);

HB1xp67_ASAP7_75t_L g13951 ( 
.A(n_13754),
.Y(n_13951)
);

INVx1_ASAP7_75t_L g13952 ( 
.A(n_13778),
.Y(n_13952)
);

INVx1_ASAP7_75t_L g13953 ( 
.A(n_13804),
.Y(n_13953)
);

AND2x2_ASAP7_75t_L g13954 ( 
.A(n_13761),
.B(n_13480),
.Y(n_13954)
);

AND2x2_ASAP7_75t_L g13955 ( 
.A(n_13777),
.B(n_13515),
.Y(n_13955)
);

OAI22xp5_ASAP7_75t_L g13956 ( 
.A1(n_13769),
.A2(n_13516),
.B1(n_13404),
.B2(n_13561),
.Y(n_13956)
);

INVx1_ASAP7_75t_L g13957 ( 
.A(n_13704),
.Y(n_13957)
);

AND2x2_ASAP7_75t_L g13958 ( 
.A(n_13728),
.B(n_13479),
.Y(n_13958)
);

AND2x4_ASAP7_75t_L g13959 ( 
.A(n_13710),
.B(n_13643),
.Y(n_13959)
);

OR2x2_ASAP7_75t_L g13960 ( 
.A(n_13676),
.B(n_13562),
.Y(n_13960)
);

INVx1_ASAP7_75t_L g13961 ( 
.A(n_13838),
.Y(n_13961)
);

INVx2_ASAP7_75t_L g13962 ( 
.A(n_13748),
.Y(n_13962)
);

NAND2xp5_ASAP7_75t_L g13963 ( 
.A(n_13784),
.B(n_13544),
.Y(n_13963)
);

INVx1_ASAP7_75t_L g13964 ( 
.A(n_13791),
.Y(n_13964)
);

AND2x2_ASAP7_75t_L g13965 ( 
.A(n_13700),
.B(n_13702),
.Y(n_13965)
);

NAND2xp5_ASAP7_75t_L g13966 ( 
.A(n_13765),
.B(n_13635),
.Y(n_13966)
);

AND2x2_ASAP7_75t_L g13967 ( 
.A(n_13706),
.B(n_13709),
.Y(n_13967)
);

INVx1_ASAP7_75t_SL g13968 ( 
.A(n_13785),
.Y(n_13968)
);

INVx2_ASAP7_75t_L g13969 ( 
.A(n_13744),
.Y(n_13969)
);

AOI22xp33_ASAP7_75t_SL g13970 ( 
.A1(n_13741),
.A2(n_13843),
.B1(n_13822),
.B2(n_13722),
.Y(n_13970)
);

OAI22xp5_ASAP7_75t_L g13971 ( 
.A1(n_13799),
.A2(n_13619),
.B1(n_13581),
.B2(n_13595),
.Y(n_13971)
);

INVx2_ASAP7_75t_L g13972 ( 
.A(n_13745),
.Y(n_13972)
);

AND2x4_ASAP7_75t_L g13973 ( 
.A(n_13730),
.B(n_13582),
.Y(n_13973)
);

INVx2_ASAP7_75t_L g13974 ( 
.A(n_13815),
.Y(n_13974)
);

OR2x2_ASAP7_75t_L g13975 ( 
.A(n_13844),
.B(n_13614),
.Y(n_13975)
);

INVx2_ASAP7_75t_L g13976 ( 
.A(n_13770),
.Y(n_13976)
);

INVx1_ASAP7_75t_L g13977 ( 
.A(n_13805),
.Y(n_13977)
);

AND2x2_ASAP7_75t_L g13978 ( 
.A(n_13849),
.B(n_13637),
.Y(n_13978)
);

NAND2xp5_ASAP7_75t_L g13979 ( 
.A(n_13827),
.B(n_13840),
.Y(n_13979)
);

NAND2x1_ASAP7_75t_L g13980 ( 
.A(n_13795),
.B(n_13437),
.Y(n_13980)
);

BUFx2_ASAP7_75t_L g13981 ( 
.A(n_13764),
.Y(n_13981)
);

AND2x2_ASAP7_75t_L g13982 ( 
.A(n_13818),
.B(n_2439),
.Y(n_13982)
);

AND2x2_ASAP7_75t_L g13983 ( 
.A(n_13821),
.B(n_2440),
.Y(n_13983)
);

OR2x2_ASAP7_75t_L g13984 ( 
.A(n_13688),
.B(n_13586),
.Y(n_13984)
);

INVx4_ASAP7_75t_L g13985 ( 
.A(n_13832),
.Y(n_13985)
);

AND2x2_ASAP7_75t_L g13986 ( 
.A(n_13841),
.B(n_2440),
.Y(n_13986)
);

AND2x2_ASAP7_75t_L g13987 ( 
.A(n_13751),
.B(n_2441),
.Y(n_13987)
);

BUFx3_ASAP7_75t_L g13988 ( 
.A(n_13832),
.Y(n_13988)
);

INVx3_ASAP7_75t_L g13989 ( 
.A(n_13825),
.Y(n_13989)
);

INVx2_ASAP7_75t_L g13990 ( 
.A(n_13747),
.Y(n_13990)
);

INVx1_ASAP7_75t_L g13991 ( 
.A(n_13839),
.Y(n_13991)
);

INVx1_ASAP7_75t_L g13992 ( 
.A(n_13763),
.Y(n_13992)
);

INVx2_ASAP7_75t_L g13993 ( 
.A(n_13750),
.Y(n_13993)
);

AOI22xp33_ASAP7_75t_L g13994 ( 
.A1(n_13776),
.A2(n_13828),
.B1(n_13831),
.B2(n_13824),
.Y(n_13994)
);

AND2x2_ASAP7_75t_L g13995 ( 
.A(n_13811),
.B(n_2441),
.Y(n_13995)
);

AND2x2_ASAP7_75t_L g13996 ( 
.A(n_13812),
.B(n_13771),
.Y(n_13996)
);

OAI22xp5_ASAP7_75t_L g13997 ( 
.A1(n_13775),
.A2(n_13558),
.B1(n_13638),
.B2(n_2444),
.Y(n_13997)
);

INVx1_ASAP7_75t_L g13998 ( 
.A(n_13772),
.Y(n_13998)
);

AND2x2_ASAP7_75t_L g13999 ( 
.A(n_13774),
.B(n_2442),
.Y(n_13999)
);

NAND2xp5_ASAP7_75t_L g14000 ( 
.A(n_13779),
.B(n_13817),
.Y(n_14000)
);

INVx2_ASAP7_75t_L g14001 ( 
.A(n_13847),
.Y(n_14001)
);

AOI22xp33_ASAP7_75t_L g14002 ( 
.A1(n_13833),
.A2(n_2444),
.B1(n_2442),
.B2(n_2443),
.Y(n_14002)
);

INVx1_ASAP7_75t_L g14003 ( 
.A(n_13848),
.Y(n_14003)
);

INVx1_ASAP7_75t_L g14004 ( 
.A(n_13810),
.Y(n_14004)
);

INVx1_ASAP7_75t_L g14005 ( 
.A(n_13678),
.Y(n_14005)
);

NAND2xp5_ASAP7_75t_L g14006 ( 
.A(n_13859),
.B(n_13845),
.Y(n_14006)
);

INVx1_ASAP7_75t_L g14007 ( 
.A(n_13920),
.Y(n_14007)
);

INVx2_ASAP7_75t_L g14008 ( 
.A(n_13854),
.Y(n_14008)
);

AND2x2_ASAP7_75t_L g14009 ( 
.A(n_13872),
.B(n_13796),
.Y(n_14009)
);

AND2x2_ASAP7_75t_L g14010 ( 
.A(n_13901),
.B(n_13836),
.Y(n_14010)
);

INVx4_ASAP7_75t_L g14011 ( 
.A(n_13915),
.Y(n_14011)
);

NOR2xp33_ASAP7_75t_L g14012 ( 
.A(n_13856),
.B(n_13813),
.Y(n_14012)
);

INVx2_ASAP7_75t_L g14013 ( 
.A(n_13889),
.Y(n_14013)
);

INVx2_ASAP7_75t_L g14014 ( 
.A(n_13987),
.Y(n_14014)
);

OR2x2_ASAP7_75t_L g14015 ( 
.A(n_13850),
.B(n_13752),
.Y(n_14015)
);

NOR2xp33_ASAP7_75t_SL g14016 ( 
.A(n_13985),
.B(n_13814),
.Y(n_14016)
);

INVx1_ASAP7_75t_L g14017 ( 
.A(n_13935),
.Y(n_14017)
);

INVx3_ASAP7_75t_L g14018 ( 
.A(n_13989),
.Y(n_14018)
);

INVx1_ASAP7_75t_L g14019 ( 
.A(n_13948),
.Y(n_14019)
);

OR2x2_ASAP7_75t_L g14020 ( 
.A(n_13912),
.B(n_13736),
.Y(n_14020)
);

INVx2_ASAP7_75t_L g14021 ( 
.A(n_13995),
.Y(n_14021)
);

AND2x4_ASAP7_75t_L g14022 ( 
.A(n_13878),
.B(n_13749),
.Y(n_14022)
);

OR2x2_ASAP7_75t_L g14023 ( 
.A(n_13857),
.B(n_13731),
.Y(n_14023)
);

INVx1_ASAP7_75t_L g14024 ( 
.A(n_13863),
.Y(n_14024)
);

AND2x4_ASAP7_75t_L g14025 ( 
.A(n_13925),
.B(n_13820),
.Y(n_14025)
);

OR2x2_ASAP7_75t_L g14026 ( 
.A(n_13942),
.B(n_13846),
.Y(n_14026)
);

INVx2_ASAP7_75t_SL g14027 ( 
.A(n_13938),
.Y(n_14027)
);

INVx1_ASAP7_75t_L g14028 ( 
.A(n_13919),
.Y(n_14028)
);

OR2x2_ASAP7_75t_L g14029 ( 
.A(n_13981),
.B(n_13773),
.Y(n_14029)
);

AND2x4_ASAP7_75t_L g14030 ( 
.A(n_13924),
.B(n_13794),
.Y(n_14030)
);

INVx1_ASAP7_75t_L g14031 ( 
.A(n_13969),
.Y(n_14031)
);

INVx1_ASAP7_75t_L g14032 ( 
.A(n_13972),
.Y(n_14032)
);

AOI21xp33_ASAP7_75t_L g14033 ( 
.A1(n_13979),
.A2(n_13652),
.B(n_13670),
.Y(n_14033)
);

INVx1_ASAP7_75t_L g14034 ( 
.A(n_13976),
.Y(n_14034)
);

AND2x2_ASAP7_75t_L g14035 ( 
.A(n_13861),
.B(n_13816),
.Y(n_14035)
);

NAND2xp5_ASAP7_75t_L g14036 ( 
.A(n_13999),
.B(n_13802),
.Y(n_14036)
);

AND2x2_ASAP7_75t_L g14037 ( 
.A(n_13930),
.B(n_13968),
.Y(n_14037)
);

INVx2_ASAP7_75t_L g14038 ( 
.A(n_13890),
.Y(n_14038)
);

OR2x2_ASAP7_75t_L g14039 ( 
.A(n_13899),
.B(n_13837),
.Y(n_14039)
);

NAND2xp5_ASAP7_75t_L g14040 ( 
.A(n_13953),
.B(n_13808),
.Y(n_14040)
);

INVxp67_ASAP7_75t_SL g14041 ( 
.A(n_13877),
.Y(n_14041)
);

AND2x4_ASAP7_75t_L g14042 ( 
.A(n_13988),
.B(n_13826),
.Y(n_14042)
);

AND2x2_ASAP7_75t_L g14043 ( 
.A(n_13902),
.B(n_13819),
.Y(n_14043)
);

AND2x2_ASAP7_75t_L g14044 ( 
.A(n_13871),
.B(n_13842),
.Y(n_14044)
);

INVx1_ASAP7_75t_L g14045 ( 
.A(n_13982),
.Y(n_14045)
);

NAND2xp5_ASAP7_75t_L g14046 ( 
.A(n_13911),
.B(n_13823),
.Y(n_14046)
);

OR2x2_ASAP7_75t_L g14047 ( 
.A(n_13853),
.B(n_13809),
.Y(n_14047)
);

INVx1_ASAP7_75t_L g14048 ( 
.A(n_13983),
.Y(n_14048)
);

AND2x2_ASAP7_75t_L g14049 ( 
.A(n_13883),
.B(n_13789),
.Y(n_14049)
);

HB1xp67_ASAP7_75t_L g14050 ( 
.A(n_13929),
.Y(n_14050)
);

HB1xp67_ASAP7_75t_L g14051 ( 
.A(n_13882),
.Y(n_14051)
);

AND3x1_ASAP7_75t_L g14052 ( 
.A(n_13962),
.B(n_13834),
.C(n_13790),
.Y(n_14052)
);

INVx1_ASAP7_75t_L g14053 ( 
.A(n_13986),
.Y(n_14053)
);

INVx2_ASAP7_75t_L g14054 ( 
.A(n_14001),
.Y(n_14054)
);

INVx1_ASAP7_75t_L g14055 ( 
.A(n_13868),
.Y(n_14055)
);

AND2x4_ASAP7_75t_L g14056 ( 
.A(n_13905),
.B(n_13782),
.Y(n_14056)
);

AND2x2_ASAP7_75t_L g14057 ( 
.A(n_13860),
.B(n_13798),
.Y(n_14057)
);

OR2x2_ASAP7_75t_L g14058 ( 
.A(n_13944),
.B(n_13720),
.Y(n_14058)
);

NAND2xp5_ASAP7_75t_L g14059 ( 
.A(n_13909),
.B(n_13781),
.Y(n_14059)
);

INVx1_ASAP7_75t_L g14060 ( 
.A(n_13870),
.Y(n_14060)
);

INVx3_ASAP7_75t_L g14061 ( 
.A(n_13862),
.Y(n_14061)
);

INVx1_ASAP7_75t_L g14062 ( 
.A(n_13852),
.Y(n_14062)
);

INVxp67_ASAP7_75t_L g14063 ( 
.A(n_13855),
.Y(n_14063)
);

INVx2_ASAP7_75t_L g14064 ( 
.A(n_13934),
.Y(n_14064)
);

NAND2xp5_ASAP7_75t_L g14065 ( 
.A(n_13970),
.B(n_13807),
.Y(n_14065)
);

AND2x2_ASAP7_75t_L g14066 ( 
.A(n_13867),
.B(n_13800),
.Y(n_14066)
);

AND2x2_ASAP7_75t_L g14067 ( 
.A(n_13881),
.B(n_13783),
.Y(n_14067)
);

OR2x2_ASAP7_75t_L g14068 ( 
.A(n_13893),
.B(n_2443),
.Y(n_14068)
);

NOR2x1_ASAP7_75t_L g14069 ( 
.A(n_13864),
.B(n_2445),
.Y(n_14069)
);

INVx2_ASAP7_75t_SL g14070 ( 
.A(n_13906),
.Y(n_14070)
);

INVx3_ASAP7_75t_L g14071 ( 
.A(n_13907),
.Y(n_14071)
);

NAND2xp5_ASAP7_75t_L g14072 ( 
.A(n_13884),
.B(n_2446),
.Y(n_14072)
);

AND2x2_ASAP7_75t_L g14073 ( 
.A(n_13903),
.B(n_2446),
.Y(n_14073)
);

AND2x2_ASAP7_75t_L g14074 ( 
.A(n_13895),
.B(n_2447),
.Y(n_14074)
);

INVx1_ASAP7_75t_L g14075 ( 
.A(n_13951),
.Y(n_14075)
);

INVx1_ASAP7_75t_L g14076 ( 
.A(n_13892),
.Y(n_14076)
);

HB1xp67_ASAP7_75t_L g14077 ( 
.A(n_13996),
.Y(n_14077)
);

INVx2_ASAP7_75t_L g14078 ( 
.A(n_13993),
.Y(n_14078)
);

AND2x6_ASAP7_75t_SL g14079 ( 
.A(n_14000),
.B(n_2447),
.Y(n_14079)
);

INVx1_ASAP7_75t_L g14080 ( 
.A(n_13961),
.Y(n_14080)
);

INVx1_ASAP7_75t_L g14081 ( 
.A(n_14004),
.Y(n_14081)
);

OR2x2_ASAP7_75t_L g14082 ( 
.A(n_13865),
.B(n_2448),
.Y(n_14082)
);

AND2x4_ASAP7_75t_L g14083 ( 
.A(n_13908),
.B(n_2449),
.Y(n_14083)
);

AND2x2_ASAP7_75t_L g14084 ( 
.A(n_13914),
.B(n_2449),
.Y(n_14084)
);

BUFx2_ASAP7_75t_L g14085 ( 
.A(n_13932),
.Y(n_14085)
);

INVxp67_ASAP7_75t_SL g14086 ( 
.A(n_13980),
.Y(n_14086)
);

INVx3_ASAP7_75t_L g14087 ( 
.A(n_13965),
.Y(n_14087)
);

INVx1_ASAP7_75t_L g14088 ( 
.A(n_13991),
.Y(n_14088)
);

INVx1_ASAP7_75t_L g14089 ( 
.A(n_13990),
.Y(n_14089)
);

INVx1_ASAP7_75t_L g14090 ( 
.A(n_13875),
.Y(n_14090)
);

NAND2xp5_ASAP7_75t_L g14091 ( 
.A(n_13955),
.B(n_2450),
.Y(n_14091)
);

OR2x2_ASAP7_75t_L g14092 ( 
.A(n_13992),
.B(n_13998),
.Y(n_14092)
);

INVx1_ASAP7_75t_L g14093 ( 
.A(n_13869),
.Y(n_14093)
);

INVx1_ASAP7_75t_L g14094 ( 
.A(n_13897),
.Y(n_14094)
);

INVx2_ASAP7_75t_L g14095 ( 
.A(n_13898),
.Y(n_14095)
);

AND2x4_ASAP7_75t_L g14096 ( 
.A(n_13858),
.B(n_2450),
.Y(n_14096)
);

AND2x2_ASAP7_75t_L g14097 ( 
.A(n_13885),
.B(n_2451),
.Y(n_14097)
);

INVx2_ASAP7_75t_L g14098 ( 
.A(n_13873),
.Y(n_14098)
);

NAND2xp5_ASAP7_75t_SL g14099 ( 
.A(n_13913),
.B(n_2451),
.Y(n_14099)
);

INVx2_ASAP7_75t_L g14100 ( 
.A(n_13959),
.Y(n_14100)
);

AND2x2_ASAP7_75t_L g14101 ( 
.A(n_13945),
.B(n_2452),
.Y(n_14101)
);

INVx2_ASAP7_75t_L g14102 ( 
.A(n_13896),
.Y(n_14102)
);

INVx2_ASAP7_75t_L g14103 ( 
.A(n_13879),
.Y(n_14103)
);

AOI22x1_ASAP7_75t_L g14104 ( 
.A1(n_13876),
.A2(n_2455),
.B1(n_2453),
.B2(n_2454),
.Y(n_14104)
);

AOI22xp33_ASAP7_75t_L g14105 ( 
.A1(n_14005),
.A2(n_2456),
.B1(n_2453),
.B2(n_2454),
.Y(n_14105)
);

AND2x4_ASAP7_75t_L g14106 ( 
.A(n_13874),
.B(n_2456),
.Y(n_14106)
);

NAND2xp5_ASAP7_75t_L g14107 ( 
.A(n_13918),
.B(n_2457),
.Y(n_14107)
);

OR2x2_ASAP7_75t_L g14108 ( 
.A(n_13940),
.B(n_2457),
.Y(n_14108)
);

AND2x4_ASAP7_75t_L g14109 ( 
.A(n_13886),
.B(n_2458),
.Y(n_14109)
);

INVx1_ASAP7_75t_L g14110 ( 
.A(n_13851),
.Y(n_14110)
);

INVx2_ASAP7_75t_L g14111 ( 
.A(n_13922),
.Y(n_14111)
);

AND2x2_ASAP7_75t_L g14112 ( 
.A(n_13928),
.B(n_2458),
.Y(n_14112)
);

INVx1_ASAP7_75t_L g14113 ( 
.A(n_13910),
.Y(n_14113)
);

INVx1_ASAP7_75t_L g14114 ( 
.A(n_13917),
.Y(n_14114)
);

INVx1_ASAP7_75t_L g14115 ( 
.A(n_13921),
.Y(n_14115)
);

NAND2xp5_ASAP7_75t_L g14116 ( 
.A(n_13978),
.B(n_2459),
.Y(n_14116)
);

INVx1_ASAP7_75t_L g14117 ( 
.A(n_13866),
.Y(n_14117)
);

INVx1_ASAP7_75t_L g14118 ( 
.A(n_13880),
.Y(n_14118)
);

AND2x2_ASAP7_75t_L g14119 ( 
.A(n_13964),
.B(n_2459),
.Y(n_14119)
);

AND2x2_ASAP7_75t_L g14120 ( 
.A(n_13977),
.B(n_2460),
.Y(n_14120)
);

AND2x2_ASAP7_75t_L g14121 ( 
.A(n_13967),
.B(n_2460),
.Y(n_14121)
);

INVx2_ASAP7_75t_L g14122 ( 
.A(n_13974),
.Y(n_14122)
);

NAND2xp5_ASAP7_75t_L g14123 ( 
.A(n_13973),
.B(n_2461),
.Y(n_14123)
);

INVx1_ASAP7_75t_L g14124 ( 
.A(n_13888),
.Y(n_14124)
);

AND2x4_ASAP7_75t_L g14125 ( 
.A(n_13900),
.B(n_2461),
.Y(n_14125)
);

INVxp67_ASAP7_75t_SL g14126 ( 
.A(n_13939),
.Y(n_14126)
);

AND2x2_ASAP7_75t_L g14127 ( 
.A(n_13933),
.B(n_2463),
.Y(n_14127)
);

INVx2_ASAP7_75t_SL g14128 ( 
.A(n_13916),
.Y(n_14128)
);

NAND2xp5_ASAP7_75t_L g14129 ( 
.A(n_14003),
.B(n_13950),
.Y(n_14129)
);

NAND2xp5_ASAP7_75t_L g14130 ( 
.A(n_13954),
.B(n_2463),
.Y(n_14130)
);

NAND2xp5_ASAP7_75t_L g14131 ( 
.A(n_13958),
.B(n_2464),
.Y(n_14131)
);

OR2x2_ASAP7_75t_L g14132 ( 
.A(n_13957),
.B(n_2464),
.Y(n_14132)
);

INVx1_ASAP7_75t_L g14133 ( 
.A(n_13975),
.Y(n_14133)
);

INVx2_ASAP7_75t_L g14134 ( 
.A(n_13943),
.Y(n_14134)
);

AND2x2_ASAP7_75t_L g14135 ( 
.A(n_13926),
.B(n_2465),
.Y(n_14135)
);

INVx2_ASAP7_75t_L g14136 ( 
.A(n_13946),
.Y(n_14136)
);

AND2x2_ASAP7_75t_L g14137 ( 
.A(n_13927),
.B(n_2465),
.Y(n_14137)
);

INVx1_ASAP7_75t_L g14138 ( 
.A(n_13931),
.Y(n_14138)
);

AND2x4_ASAP7_75t_L g14139 ( 
.A(n_14037),
.B(n_13936),
.Y(n_14139)
);

NOR2x1p5_ASAP7_75t_L g14140 ( 
.A(n_14018),
.B(n_13923),
.Y(n_14140)
);

AND2x2_ASAP7_75t_L g14141 ( 
.A(n_14009),
.B(n_13937),
.Y(n_14141)
);

HB1xp67_ASAP7_75t_L g14142 ( 
.A(n_14051),
.Y(n_14142)
);

NOR2xp33_ASAP7_75t_R g14143 ( 
.A(n_14071),
.B(n_13941),
.Y(n_14143)
);

INVxp67_ASAP7_75t_L g14144 ( 
.A(n_14077),
.Y(n_14144)
);

OAI211xp5_ASAP7_75t_L g14145 ( 
.A1(n_14086),
.A2(n_13949),
.B(n_13952),
.C(n_13947),
.Y(n_14145)
);

AND2x2_ASAP7_75t_L g14146 ( 
.A(n_14038),
.B(n_13997),
.Y(n_14146)
);

INVx1_ASAP7_75t_L g14147 ( 
.A(n_14010),
.Y(n_14147)
);

INVx1_ASAP7_75t_L g14148 ( 
.A(n_14085),
.Y(n_14148)
);

AOI22xp5_ASAP7_75t_L g14149 ( 
.A1(n_14128),
.A2(n_13887),
.B1(n_13904),
.B2(n_13960),
.Y(n_14149)
);

AND2x4_ASAP7_75t_L g14150 ( 
.A(n_14022),
.B(n_14011),
.Y(n_14150)
);

AND2x2_ASAP7_75t_L g14151 ( 
.A(n_14035),
.B(n_13894),
.Y(n_14151)
);

NAND2xp5_ASAP7_75t_L g14152 ( 
.A(n_14083),
.B(n_14002),
.Y(n_14152)
);

NAND2xp5_ASAP7_75t_L g14153 ( 
.A(n_14084),
.B(n_13891),
.Y(n_14153)
);

OR2x2_ASAP7_75t_L g14154 ( 
.A(n_14029),
.B(n_13984),
.Y(n_14154)
);

INVx2_ASAP7_75t_L g14155 ( 
.A(n_14127),
.Y(n_14155)
);

INVx2_ASAP7_75t_L g14156 ( 
.A(n_14104),
.Y(n_14156)
);

HB1xp67_ASAP7_75t_L g14157 ( 
.A(n_14063),
.Y(n_14157)
);

AND2x2_ASAP7_75t_L g14158 ( 
.A(n_14008),
.B(n_14013),
.Y(n_14158)
);

OR2x6_ASAP7_75t_L g14159 ( 
.A(n_14064),
.B(n_14007),
.Y(n_14159)
);

HB1xp67_ASAP7_75t_L g14160 ( 
.A(n_14017),
.Y(n_14160)
);

AND2x4_ASAP7_75t_L g14161 ( 
.A(n_14027),
.B(n_13963),
.Y(n_14161)
);

BUFx3_ASAP7_75t_L g14162 ( 
.A(n_14042),
.Y(n_14162)
);

INVx2_ASAP7_75t_L g14163 ( 
.A(n_14109),
.Y(n_14163)
);

INVx2_ASAP7_75t_L g14164 ( 
.A(n_14097),
.Y(n_14164)
);

INVx2_ASAP7_75t_SL g14165 ( 
.A(n_14087),
.Y(n_14165)
);

OAI22xp5_ASAP7_75t_L g14166 ( 
.A1(n_14015),
.A2(n_14041),
.B1(n_14020),
.B2(n_14023),
.Y(n_14166)
);

AND2x4_ASAP7_75t_L g14167 ( 
.A(n_14070),
.B(n_13966),
.Y(n_14167)
);

AOI221xp5_ASAP7_75t_L g14168 ( 
.A1(n_14033),
.A2(n_13994),
.B1(n_13956),
.B2(n_13971),
.C(n_2468),
.Y(n_14168)
);

AND2x2_ASAP7_75t_L g14169 ( 
.A(n_14050),
.B(n_2466),
.Y(n_14169)
);

AND2x2_ASAP7_75t_L g14170 ( 
.A(n_14043),
.B(n_2466),
.Y(n_14170)
);

INVx2_ASAP7_75t_L g14171 ( 
.A(n_14096),
.Y(n_14171)
);

INVx1_ASAP7_75t_L g14172 ( 
.A(n_14026),
.Y(n_14172)
);

NAND2xp5_ASAP7_75t_L g14173 ( 
.A(n_14121),
.B(n_2467),
.Y(n_14173)
);

NOR2xp33_ASAP7_75t_L g14174 ( 
.A(n_14016),
.B(n_2467),
.Y(n_14174)
);

AND2x2_ASAP7_75t_L g14175 ( 
.A(n_14061),
.B(n_2468),
.Y(n_14175)
);

AND2x2_ASAP7_75t_L g14176 ( 
.A(n_14117),
.B(n_2469),
.Y(n_14176)
);

INVx1_ASAP7_75t_L g14177 ( 
.A(n_14103),
.Y(n_14177)
);

INVx3_ASAP7_75t_L g14178 ( 
.A(n_14106),
.Y(n_14178)
);

AND2x4_ASAP7_75t_L g14179 ( 
.A(n_14078),
.B(n_2470),
.Y(n_14179)
);

AOI221xp5_ASAP7_75t_L g14180 ( 
.A1(n_14052),
.A2(n_14065),
.B1(n_14032),
.B2(n_14034),
.C(n_14031),
.Y(n_14180)
);

INVx5_ASAP7_75t_L g14181 ( 
.A(n_14125),
.Y(n_14181)
);

INVx3_ASAP7_75t_L g14182 ( 
.A(n_14030),
.Y(n_14182)
);

HB1xp67_ASAP7_75t_L g14183 ( 
.A(n_14069),
.Y(n_14183)
);

INVx1_ASAP7_75t_SL g14184 ( 
.A(n_14112),
.Y(n_14184)
);

BUFx2_ASAP7_75t_L g14185 ( 
.A(n_14049),
.Y(n_14185)
);

NAND2xp5_ASAP7_75t_L g14186 ( 
.A(n_14021),
.B(n_2470),
.Y(n_14186)
);

HB1xp67_ASAP7_75t_L g14187 ( 
.A(n_14073),
.Y(n_14187)
);

BUFx2_ASAP7_75t_L g14188 ( 
.A(n_14019),
.Y(n_14188)
);

AND2x2_ASAP7_75t_SL g14189 ( 
.A(n_14025),
.B(n_2471),
.Y(n_14189)
);

OAI32xp33_ASAP7_75t_L g14190 ( 
.A1(n_14058),
.A2(n_2473),
.A3(n_2471),
.B1(n_2472),
.B2(n_2474),
.Y(n_14190)
);

AND2x2_ASAP7_75t_L g14191 ( 
.A(n_14076),
.B(n_2472),
.Y(n_14191)
);

INVx1_ASAP7_75t_L g14192 ( 
.A(n_14098),
.Y(n_14192)
);

NOR2x1_ASAP7_75t_L g14193 ( 
.A(n_14088),
.B(n_2473),
.Y(n_14193)
);

OAI211xp5_ASAP7_75t_L g14194 ( 
.A1(n_14075),
.A2(n_2476),
.B(n_2474),
.C(n_2475),
.Y(n_14194)
);

NOR2xp33_ASAP7_75t_L g14195 ( 
.A(n_14079),
.B(n_14108),
.Y(n_14195)
);

INVx1_ASAP7_75t_L g14196 ( 
.A(n_14101),
.Y(n_14196)
);

NAND3xp33_ASAP7_75t_L g14197 ( 
.A(n_14012),
.B(n_2475),
.C(n_2477),
.Y(n_14197)
);

OR2x2_ASAP7_75t_L g14198 ( 
.A(n_14092),
.B(n_2477),
.Y(n_14198)
);

NAND2xp5_ASAP7_75t_L g14199 ( 
.A(n_14014),
.B(n_2478),
.Y(n_14199)
);

NOR2xp33_ASAP7_75t_L g14200 ( 
.A(n_14082),
.B(n_2478),
.Y(n_14200)
);

INVx1_ASAP7_75t_L g14201 ( 
.A(n_14074),
.Y(n_14201)
);

INVx1_ASAP7_75t_L g14202 ( 
.A(n_14091),
.Y(n_14202)
);

INVx3_ASAP7_75t_L g14203 ( 
.A(n_14056),
.Y(n_14203)
);

INVx1_ASAP7_75t_SL g14204 ( 
.A(n_14066),
.Y(n_14204)
);

NOR2xp33_ASAP7_75t_L g14205 ( 
.A(n_14036),
.B(n_2479),
.Y(n_14205)
);

BUFx3_ASAP7_75t_L g14206 ( 
.A(n_14028),
.Y(n_14206)
);

INVx1_ASAP7_75t_L g14207 ( 
.A(n_14107),
.Y(n_14207)
);

OR2x2_ASAP7_75t_L g14208 ( 
.A(n_14040),
.B(n_2479),
.Y(n_14208)
);

OR2x2_ASAP7_75t_L g14209 ( 
.A(n_14047),
.B(n_2480),
.Y(n_14209)
);

INVx1_ASAP7_75t_L g14210 ( 
.A(n_14068),
.Y(n_14210)
);

INVx2_ASAP7_75t_L g14211 ( 
.A(n_14111),
.Y(n_14211)
);

OR2x2_ASAP7_75t_L g14212 ( 
.A(n_14080),
.B(n_2480),
.Y(n_14212)
);

INVx1_ASAP7_75t_L g14213 ( 
.A(n_14135),
.Y(n_14213)
);

AOI22xp33_ASAP7_75t_L g14214 ( 
.A1(n_14126),
.A2(n_2483),
.B1(n_2481),
.B2(n_2482),
.Y(n_14214)
);

CKINVDCx5p33_ASAP7_75t_R g14215 ( 
.A(n_14116),
.Y(n_14215)
);

INVx1_ASAP7_75t_L g14216 ( 
.A(n_14137),
.Y(n_14216)
);

AND2x2_ASAP7_75t_L g14217 ( 
.A(n_14110),
.B(n_2481),
.Y(n_14217)
);

OR2x2_ASAP7_75t_L g14218 ( 
.A(n_14094),
.B(n_2482),
.Y(n_14218)
);

INVx1_ASAP7_75t_L g14219 ( 
.A(n_14131),
.Y(n_14219)
);

INVx1_ASAP7_75t_L g14220 ( 
.A(n_14119),
.Y(n_14220)
);

OR2x2_ASAP7_75t_L g14221 ( 
.A(n_14039),
.B(n_2483),
.Y(n_14221)
);

AND2x2_ASAP7_75t_L g14222 ( 
.A(n_14067),
.B(n_2484),
.Y(n_14222)
);

INVx2_ASAP7_75t_L g14223 ( 
.A(n_14134),
.Y(n_14223)
);

NAND2xp5_ASAP7_75t_L g14224 ( 
.A(n_14045),
.B(n_14048),
.Y(n_14224)
);

INVx2_ASAP7_75t_L g14225 ( 
.A(n_14102),
.Y(n_14225)
);

INVx1_ASAP7_75t_L g14226 ( 
.A(n_14120),
.Y(n_14226)
);

BUFx2_ASAP7_75t_L g14227 ( 
.A(n_14006),
.Y(n_14227)
);

AND2x2_ASAP7_75t_L g14228 ( 
.A(n_14024),
.B(n_2484),
.Y(n_14228)
);

INVx2_ASAP7_75t_L g14229 ( 
.A(n_14100),
.Y(n_14229)
);

INVxp67_ASAP7_75t_SL g14230 ( 
.A(n_14129),
.Y(n_14230)
);

OR2x2_ASAP7_75t_L g14231 ( 
.A(n_14124),
.B(n_2485),
.Y(n_14231)
);

INVxp67_ASAP7_75t_SL g14232 ( 
.A(n_14099),
.Y(n_14232)
);

INVxp67_ASAP7_75t_SL g14233 ( 
.A(n_14130),
.Y(n_14233)
);

INVx2_ASAP7_75t_L g14234 ( 
.A(n_14132),
.Y(n_14234)
);

NAND2xp5_ASAP7_75t_L g14235 ( 
.A(n_14053),
.B(n_2486),
.Y(n_14235)
);

INVx2_ASAP7_75t_L g14236 ( 
.A(n_14095),
.Y(n_14236)
);

INVx1_ASAP7_75t_L g14237 ( 
.A(n_14123),
.Y(n_14237)
);

AND2x2_ASAP7_75t_L g14238 ( 
.A(n_14062),
.B(n_2486),
.Y(n_14238)
);

AND2x2_ASAP7_75t_L g14239 ( 
.A(n_14057),
.B(n_2487),
.Y(n_14239)
);

NAND2xp5_ASAP7_75t_L g14240 ( 
.A(n_14093),
.B(n_14054),
.Y(n_14240)
);

NAND3xp33_ASAP7_75t_SL g14241 ( 
.A(n_14133),
.B(n_2487),
.C(n_2488),
.Y(n_14241)
);

BUFx2_ASAP7_75t_L g14242 ( 
.A(n_14113),
.Y(n_14242)
);

OAI22xp5_ASAP7_75t_SL g14243 ( 
.A1(n_14118),
.A2(n_14059),
.B1(n_14090),
.B2(n_14138),
.Y(n_14243)
);

NAND2xp5_ASAP7_75t_L g14244 ( 
.A(n_14044),
.B(n_14105),
.Y(n_14244)
);

AND2x2_ASAP7_75t_L g14245 ( 
.A(n_14114),
.B(n_2489),
.Y(n_14245)
);

AND2x2_ASAP7_75t_L g14246 ( 
.A(n_14115),
.B(n_2489),
.Y(n_14246)
);

INVx1_ASAP7_75t_L g14247 ( 
.A(n_14136),
.Y(n_14247)
);

OAI22xp5_ASAP7_75t_L g14248 ( 
.A1(n_14072),
.A2(n_2492),
.B1(n_2490),
.B2(n_2491),
.Y(n_14248)
);

NOR3xp33_ASAP7_75t_SL g14249 ( 
.A(n_14081),
.B(n_2490),
.C(n_2491),
.Y(n_14249)
);

INVx1_ASAP7_75t_L g14250 ( 
.A(n_14122),
.Y(n_14250)
);

BUFx3_ASAP7_75t_L g14251 ( 
.A(n_14089),
.Y(n_14251)
);

AOI222xp33_ASAP7_75t_L g14252 ( 
.A1(n_14046),
.A2(n_2495),
.B1(n_2497),
.B2(n_2493),
.C1(n_2494),
.C2(n_2496),
.Y(n_14252)
);

AND2x2_ASAP7_75t_L g14253 ( 
.A(n_14055),
.B(n_2493),
.Y(n_14253)
);

INVx1_ASAP7_75t_L g14254 ( 
.A(n_14185),
.Y(n_14254)
);

NAND2xp5_ASAP7_75t_L g14255 ( 
.A(n_14187),
.B(n_14060),
.Y(n_14255)
);

INVx1_ASAP7_75t_L g14256 ( 
.A(n_14142),
.Y(n_14256)
);

INVx1_ASAP7_75t_L g14257 ( 
.A(n_14151),
.Y(n_14257)
);

NAND2xp5_ASAP7_75t_L g14258 ( 
.A(n_14195),
.B(n_2495),
.Y(n_14258)
);

OR2x2_ASAP7_75t_L g14259 ( 
.A(n_14154),
.B(n_2496),
.Y(n_14259)
);

INVx1_ASAP7_75t_L g14260 ( 
.A(n_14167),
.Y(n_14260)
);

AND2x2_ASAP7_75t_L g14261 ( 
.A(n_14150),
.B(n_2497),
.Y(n_14261)
);

INVx4_ASAP7_75t_L g14262 ( 
.A(n_14162),
.Y(n_14262)
);

NAND2xp5_ASAP7_75t_L g14263 ( 
.A(n_14204),
.B(n_2498),
.Y(n_14263)
);

NOR2x1_ASAP7_75t_L g14264 ( 
.A(n_14140),
.B(n_14166),
.Y(n_14264)
);

AND2x2_ASAP7_75t_L g14265 ( 
.A(n_14141),
.B(n_2498),
.Y(n_14265)
);

INVx1_ASAP7_75t_L g14266 ( 
.A(n_14236),
.Y(n_14266)
);

NAND2xp5_ASAP7_75t_L g14267 ( 
.A(n_14184),
.B(n_2499),
.Y(n_14267)
);

AND2x2_ASAP7_75t_L g14268 ( 
.A(n_14158),
.B(n_2499),
.Y(n_14268)
);

NAND2x1p5_ASAP7_75t_L g14269 ( 
.A(n_14181),
.B(n_2500),
.Y(n_14269)
);

INVx1_ASAP7_75t_L g14270 ( 
.A(n_14225),
.Y(n_14270)
);

AND2x2_ASAP7_75t_L g14271 ( 
.A(n_14147),
.B(n_2501),
.Y(n_14271)
);

INVx1_ASAP7_75t_L g14272 ( 
.A(n_14169),
.Y(n_14272)
);

OR2x2_ASAP7_75t_L g14273 ( 
.A(n_14148),
.B(n_2501),
.Y(n_14273)
);

NAND2xp5_ASAP7_75t_L g14274 ( 
.A(n_14239),
.B(n_14183),
.Y(n_14274)
);

AND2x2_ASAP7_75t_L g14275 ( 
.A(n_14139),
.B(n_2502),
.Y(n_14275)
);

INVx1_ASAP7_75t_L g14276 ( 
.A(n_14172),
.Y(n_14276)
);

INVx1_ASAP7_75t_L g14277 ( 
.A(n_14221),
.Y(n_14277)
);

NAND2xp5_ASAP7_75t_L g14278 ( 
.A(n_14179),
.B(n_2502),
.Y(n_14278)
);

AND2x2_ASAP7_75t_L g14279 ( 
.A(n_14182),
.B(n_2503),
.Y(n_14279)
);

AND2x2_ASAP7_75t_L g14280 ( 
.A(n_14230),
.B(n_2503),
.Y(n_14280)
);

OR2x2_ASAP7_75t_L g14281 ( 
.A(n_14165),
.B(n_2504),
.Y(n_14281)
);

INVx1_ASAP7_75t_L g14282 ( 
.A(n_14198),
.Y(n_14282)
);

INVx4_ASAP7_75t_L g14283 ( 
.A(n_14159),
.Y(n_14283)
);

NAND2xp5_ASAP7_75t_L g14284 ( 
.A(n_14181),
.B(n_2504),
.Y(n_14284)
);

INVx1_ASAP7_75t_SL g14285 ( 
.A(n_14143),
.Y(n_14285)
);

NAND2xp5_ASAP7_75t_L g14286 ( 
.A(n_14222),
.B(n_2505),
.Y(n_14286)
);

AND2x2_ASAP7_75t_L g14287 ( 
.A(n_14159),
.B(n_2505),
.Y(n_14287)
);

INVx1_ASAP7_75t_L g14288 ( 
.A(n_14177),
.Y(n_14288)
);

INVx1_ASAP7_75t_L g14289 ( 
.A(n_14161),
.Y(n_14289)
);

NAND2x1p5_ASAP7_75t_L g14290 ( 
.A(n_14203),
.B(n_2506),
.Y(n_14290)
);

AND2x2_ASAP7_75t_L g14291 ( 
.A(n_14170),
.B(n_2506),
.Y(n_14291)
);

AND2x2_ASAP7_75t_L g14292 ( 
.A(n_14157),
.B(n_2507),
.Y(n_14292)
);

INVx2_ASAP7_75t_SL g14293 ( 
.A(n_14175),
.Y(n_14293)
);

INVx2_ASAP7_75t_L g14294 ( 
.A(n_14189),
.Y(n_14294)
);

AND2x4_ASAP7_75t_L g14295 ( 
.A(n_14178),
.B(n_2507),
.Y(n_14295)
);

INVxp67_ASAP7_75t_L g14296 ( 
.A(n_14200),
.Y(n_14296)
);

OR2x2_ASAP7_75t_L g14297 ( 
.A(n_14144),
.B(n_2508),
.Y(n_14297)
);

INVxp67_ASAP7_75t_SL g14298 ( 
.A(n_14193),
.Y(n_14298)
);

INVx1_ASAP7_75t_L g14299 ( 
.A(n_14247),
.Y(n_14299)
);

INVx1_ASAP7_75t_L g14300 ( 
.A(n_14231),
.Y(n_14300)
);

INVx1_ASAP7_75t_L g14301 ( 
.A(n_14227),
.Y(n_14301)
);

AND2x2_ASAP7_75t_L g14302 ( 
.A(n_14188),
.B(n_2508),
.Y(n_14302)
);

NAND2xp5_ASAP7_75t_L g14303 ( 
.A(n_14196),
.B(n_2509),
.Y(n_14303)
);

INVx1_ASAP7_75t_L g14304 ( 
.A(n_14229),
.Y(n_14304)
);

AND2x2_ASAP7_75t_L g14305 ( 
.A(n_14146),
.B(n_2509),
.Y(n_14305)
);

INVx1_ASAP7_75t_L g14306 ( 
.A(n_14176),
.Y(n_14306)
);

NAND2xp5_ASAP7_75t_L g14307 ( 
.A(n_14249),
.B(n_2510),
.Y(n_14307)
);

AND2x2_ASAP7_75t_L g14308 ( 
.A(n_14160),
.B(n_2511),
.Y(n_14308)
);

AND2x2_ASAP7_75t_L g14309 ( 
.A(n_14156),
.B(n_2511),
.Y(n_14309)
);

INVx1_ASAP7_75t_SL g14310 ( 
.A(n_14209),
.Y(n_14310)
);

NAND2xp5_ASAP7_75t_L g14311 ( 
.A(n_14217),
.B(n_2512),
.Y(n_14311)
);

INVx1_ASAP7_75t_L g14312 ( 
.A(n_14211),
.Y(n_14312)
);

INVx2_ASAP7_75t_L g14313 ( 
.A(n_14155),
.Y(n_14313)
);

AND2x2_ASAP7_75t_L g14314 ( 
.A(n_14242),
.B(n_2512),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_14223),
.Y(n_14315)
);

NAND2xp5_ASAP7_75t_L g14316 ( 
.A(n_14215),
.B(n_2513),
.Y(n_14316)
);

HB1xp67_ASAP7_75t_L g14317 ( 
.A(n_14206),
.Y(n_14317)
);

AND2x2_ASAP7_75t_L g14318 ( 
.A(n_14251),
.B(n_2513),
.Y(n_14318)
);

AND2x2_ASAP7_75t_L g14319 ( 
.A(n_14174),
.B(n_14228),
.Y(n_14319)
);

AND2x2_ASAP7_75t_L g14320 ( 
.A(n_14238),
.B(n_2514),
.Y(n_14320)
);

INVx1_ASAP7_75t_L g14321 ( 
.A(n_14173),
.Y(n_14321)
);

AND2x2_ASAP7_75t_L g14322 ( 
.A(n_14191),
.B(n_2514),
.Y(n_14322)
);

AND2x2_ASAP7_75t_L g14323 ( 
.A(n_14224),
.B(n_2515),
.Y(n_14323)
);

NAND2xp5_ASAP7_75t_L g14324 ( 
.A(n_14201),
.B(n_2515),
.Y(n_14324)
);

AND2x4_ASAP7_75t_L g14325 ( 
.A(n_14232),
.B(n_2516),
.Y(n_14325)
);

AND2x4_ASAP7_75t_L g14326 ( 
.A(n_14253),
.B(n_2516),
.Y(n_14326)
);

OR2x2_ASAP7_75t_L g14327 ( 
.A(n_14240),
.B(n_2517),
.Y(n_14327)
);

INVx1_ASAP7_75t_L g14328 ( 
.A(n_14164),
.Y(n_14328)
);

AND2x2_ASAP7_75t_L g14329 ( 
.A(n_14205),
.B(n_2517),
.Y(n_14329)
);

NAND2xp5_ASAP7_75t_L g14330 ( 
.A(n_14245),
.B(n_2518),
.Y(n_14330)
);

AND2x4_ASAP7_75t_L g14331 ( 
.A(n_14213),
.B(n_2518),
.Y(n_14331)
);

OR2x2_ASAP7_75t_L g14332 ( 
.A(n_14208),
.B(n_2519),
.Y(n_14332)
);

NAND2xp5_ASAP7_75t_L g14333 ( 
.A(n_14246),
.B(n_2519),
.Y(n_14333)
);

NOR2xp33_ASAP7_75t_L g14334 ( 
.A(n_14241),
.B(n_2520),
.Y(n_14334)
);

INVx2_ASAP7_75t_L g14335 ( 
.A(n_14163),
.Y(n_14335)
);

INVx1_ASAP7_75t_L g14336 ( 
.A(n_14192),
.Y(n_14336)
);

INVx1_ASAP7_75t_L g14337 ( 
.A(n_14233),
.Y(n_14337)
);

OR2x2_ASAP7_75t_L g14338 ( 
.A(n_14212),
.B(n_2520),
.Y(n_14338)
);

AND2x2_ASAP7_75t_L g14339 ( 
.A(n_14216),
.B(n_2521),
.Y(n_14339)
);

AND2x4_ASAP7_75t_L g14340 ( 
.A(n_14220),
.B(n_2521),
.Y(n_14340)
);

INVx1_ASAP7_75t_L g14341 ( 
.A(n_14218),
.Y(n_14341)
);

AND2x4_ASAP7_75t_L g14342 ( 
.A(n_14226),
.B(n_14250),
.Y(n_14342)
);

AND2x2_ASAP7_75t_L g14343 ( 
.A(n_14252),
.B(n_2522),
.Y(n_14343)
);

NAND2xp5_ASAP7_75t_L g14344 ( 
.A(n_14234),
.B(n_2522),
.Y(n_14344)
);

INVx1_ASAP7_75t_L g14345 ( 
.A(n_14210),
.Y(n_14345)
);

OR2x2_ASAP7_75t_L g14346 ( 
.A(n_14235),
.B(n_2523),
.Y(n_14346)
);

AND2x4_ASAP7_75t_L g14347 ( 
.A(n_14171),
.B(n_2523),
.Y(n_14347)
);

INVx2_ASAP7_75t_L g14348 ( 
.A(n_14207),
.Y(n_14348)
);

NAND2xp5_ASAP7_75t_L g14349 ( 
.A(n_14202),
.B(n_2525),
.Y(n_14349)
);

AND2x2_ASAP7_75t_L g14350 ( 
.A(n_14180),
.B(n_14145),
.Y(n_14350)
);

AND2x2_ASAP7_75t_L g14351 ( 
.A(n_14219),
.B(n_2525),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_14243),
.Y(n_14352)
);

NAND2xp5_ASAP7_75t_L g14353 ( 
.A(n_14214),
.B(n_2526),
.Y(n_14353)
);

INVx1_ASAP7_75t_L g14354 ( 
.A(n_14186),
.Y(n_14354)
);

NAND2x1_ASAP7_75t_L g14355 ( 
.A(n_14199),
.B(n_2526),
.Y(n_14355)
);

AND2x2_ASAP7_75t_L g14356 ( 
.A(n_14149),
.B(n_2527),
.Y(n_14356)
);

HB1xp67_ASAP7_75t_L g14357 ( 
.A(n_14244),
.Y(n_14357)
);

INVx1_ASAP7_75t_L g14358 ( 
.A(n_14153),
.Y(n_14358)
);

AND2x2_ASAP7_75t_L g14359 ( 
.A(n_14237),
.B(n_2527),
.Y(n_14359)
);

AND3x2_ASAP7_75t_L g14360 ( 
.A(n_14168),
.B(n_14152),
.C(n_14194),
.Y(n_14360)
);

AND2x2_ASAP7_75t_L g14361 ( 
.A(n_14248),
.B(n_2528),
.Y(n_14361)
);

NAND2xp5_ASAP7_75t_L g14362 ( 
.A(n_14197),
.B(n_2528),
.Y(n_14362)
);

NAND2xp5_ASAP7_75t_L g14363 ( 
.A(n_14190),
.B(n_2529),
.Y(n_14363)
);

INVx1_ASAP7_75t_L g14364 ( 
.A(n_14185),
.Y(n_14364)
);

AND2x4_ASAP7_75t_L g14365 ( 
.A(n_14150),
.B(n_2529),
.Y(n_14365)
);

NAND2xp5_ASAP7_75t_L g14366 ( 
.A(n_14185),
.B(n_2530),
.Y(n_14366)
);

NOR2xp33_ASAP7_75t_L g14367 ( 
.A(n_14181),
.B(n_2530),
.Y(n_14367)
);

OR2x2_ASAP7_75t_L g14368 ( 
.A(n_14185),
.B(n_2531),
.Y(n_14368)
);

AND2x2_ASAP7_75t_L g14369 ( 
.A(n_14150),
.B(n_2531),
.Y(n_14369)
);

INVx1_ASAP7_75t_L g14370 ( 
.A(n_14185),
.Y(n_14370)
);

NAND2xp5_ASAP7_75t_L g14371 ( 
.A(n_14185),
.B(n_2532),
.Y(n_14371)
);

INVx1_ASAP7_75t_L g14372 ( 
.A(n_14185),
.Y(n_14372)
);

INVx2_ASAP7_75t_L g14373 ( 
.A(n_14185),
.Y(n_14373)
);

AND2x2_ASAP7_75t_L g14374 ( 
.A(n_14150),
.B(n_2535),
.Y(n_14374)
);

INVx2_ASAP7_75t_L g14375 ( 
.A(n_14185),
.Y(n_14375)
);

INVx1_ASAP7_75t_L g14376 ( 
.A(n_14185),
.Y(n_14376)
);

AND2x4_ASAP7_75t_L g14377 ( 
.A(n_14150),
.B(n_2535),
.Y(n_14377)
);

INVx1_ASAP7_75t_L g14378 ( 
.A(n_14185),
.Y(n_14378)
);

INVx2_ASAP7_75t_SL g14379 ( 
.A(n_14283),
.Y(n_14379)
);

AOI22xp5_ASAP7_75t_L g14380 ( 
.A1(n_14298),
.A2(n_2538),
.B1(n_2536),
.B2(n_2537),
.Y(n_14380)
);

NAND2xp5_ASAP7_75t_L g14381 ( 
.A(n_14257),
.B(n_2536),
.Y(n_14381)
);

INVx1_ASAP7_75t_SL g14382 ( 
.A(n_14264),
.Y(n_14382)
);

INVx1_ASAP7_75t_L g14383 ( 
.A(n_14317),
.Y(n_14383)
);

AND2x2_ASAP7_75t_L g14384 ( 
.A(n_14262),
.B(n_2538),
.Y(n_14384)
);

OR2x2_ASAP7_75t_L g14385 ( 
.A(n_14373),
.B(n_2539),
.Y(n_14385)
);

AND2x2_ASAP7_75t_L g14386 ( 
.A(n_14375),
.B(n_2539),
.Y(n_14386)
);

INVx1_ASAP7_75t_L g14387 ( 
.A(n_14259),
.Y(n_14387)
);

INVx2_ASAP7_75t_L g14388 ( 
.A(n_14269),
.Y(n_14388)
);

NAND2xp5_ASAP7_75t_L g14389 ( 
.A(n_14291),
.B(n_2540),
.Y(n_14389)
);

AND2x2_ASAP7_75t_L g14390 ( 
.A(n_14289),
.B(n_2540),
.Y(n_14390)
);

OR2x2_ASAP7_75t_L g14391 ( 
.A(n_14260),
.B(n_2541),
.Y(n_14391)
);

AND2x2_ASAP7_75t_L g14392 ( 
.A(n_14254),
.B(n_2542),
.Y(n_14392)
);

INVx1_ASAP7_75t_L g14393 ( 
.A(n_14302),
.Y(n_14393)
);

OAI22xp33_ASAP7_75t_R g14394 ( 
.A1(n_14352),
.A2(n_2544),
.B1(n_2542),
.B2(n_2543),
.Y(n_14394)
);

NOR2xp33_ASAP7_75t_L g14395 ( 
.A(n_14285),
.B(n_2543),
.Y(n_14395)
);

NAND2xp5_ASAP7_75t_L g14396 ( 
.A(n_14265),
.B(n_2544),
.Y(n_14396)
);

OR2x2_ASAP7_75t_L g14397 ( 
.A(n_14364),
.B(n_2545),
.Y(n_14397)
);

INVx3_ASAP7_75t_L g14398 ( 
.A(n_14365),
.Y(n_14398)
);

NOR2x1_ASAP7_75t_L g14399 ( 
.A(n_14370),
.B(n_2545),
.Y(n_14399)
);

AOI21xp5_ASAP7_75t_L g14400 ( 
.A1(n_14350),
.A2(n_14274),
.B(n_14284),
.Y(n_14400)
);

AND2x2_ASAP7_75t_L g14401 ( 
.A(n_14372),
.B(n_2546),
.Y(n_14401)
);

INVx2_ASAP7_75t_L g14402 ( 
.A(n_14290),
.Y(n_14402)
);

NAND2xp5_ASAP7_75t_L g14403 ( 
.A(n_14326),
.B(n_2546),
.Y(n_14403)
);

AND2x4_ASAP7_75t_L g14404 ( 
.A(n_14301),
.B(n_2547),
.Y(n_14404)
);

NAND2xp5_ASAP7_75t_L g14405 ( 
.A(n_14268),
.B(n_2547),
.Y(n_14405)
);

INVx1_ASAP7_75t_SL g14406 ( 
.A(n_14368),
.Y(n_14406)
);

INVx1_ASAP7_75t_L g14407 ( 
.A(n_14357),
.Y(n_14407)
);

NAND2xp5_ASAP7_75t_L g14408 ( 
.A(n_14320),
.B(n_2548),
.Y(n_14408)
);

AND2x2_ASAP7_75t_L g14409 ( 
.A(n_14376),
.B(n_14378),
.Y(n_14409)
);

OR2x2_ASAP7_75t_L g14410 ( 
.A(n_14366),
.B(n_2549),
.Y(n_14410)
);

AND2x2_ASAP7_75t_L g14411 ( 
.A(n_14261),
.B(n_2550),
.Y(n_14411)
);

NAND2x1p5_ASAP7_75t_L g14412 ( 
.A(n_14377),
.B(n_14275),
.Y(n_14412)
);

OR2x2_ASAP7_75t_L g14413 ( 
.A(n_14371),
.B(n_2550),
.Y(n_14413)
);

OA211x2_ASAP7_75t_L g14414 ( 
.A1(n_14367),
.A2(n_2553),
.B(n_2551),
.C(n_2552),
.Y(n_14414)
);

OR2x2_ASAP7_75t_L g14415 ( 
.A(n_14255),
.B(n_14281),
.Y(n_14415)
);

AND2x2_ASAP7_75t_L g14416 ( 
.A(n_14369),
.B(n_2551),
.Y(n_14416)
);

INVxp67_ASAP7_75t_SL g14417 ( 
.A(n_14305),
.Y(n_14417)
);

AND2x2_ASAP7_75t_L g14418 ( 
.A(n_14374),
.B(n_2552),
.Y(n_14418)
);

AND2x2_ASAP7_75t_L g14419 ( 
.A(n_14342),
.B(n_2554),
.Y(n_14419)
);

AND2x2_ASAP7_75t_L g14420 ( 
.A(n_14323),
.B(n_2554),
.Y(n_14420)
);

INVxp67_ASAP7_75t_L g14421 ( 
.A(n_14287),
.Y(n_14421)
);

NAND2xp5_ASAP7_75t_L g14422 ( 
.A(n_14322),
.B(n_2555),
.Y(n_14422)
);

OR2x6_ASAP7_75t_L g14423 ( 
.A(n_14335),
.B(n_2555),
.Y(n_14423)
);

AND2x2_ASAP7_75t_L g14424 ( 
.A(n_14314),
.B(n_2556),
.Y(n_14424)
);

AND2x2_ASAP7_75t_L g14425 ( 
.A(n_14292),
.B(n_2556),
.Y(n_14425)
);

NAND3xp33_ASAP7_75t_L g14426 ( 
.A(n_14304),
.B(n_2557),
.C(n_2558),
.Y(n_14426)
);

INVx2_ASAP7_75t_L g14427 ( 
.A(n_14347),
.Y(n_14427)
);

INVx1_ASAP7_75t_L g14428 ( 
.A(n_14308),
.Y(n_14428)
);

NAND2x1p5_ASAP7_75t_L g14429 ( 
.A(n_14279),
.B(n_2557),
.Y(n_14429)
);

INVx1_ASAP7_75t_L g14430 ( 
.A(n_14332),
.Y(n_14430)
);

INVx1_ASAP7_75t_L g14431 ( 
.A(n_14286),
.Y(n_14431)
);

NAND2xp5_ASAP7_75t_L g14432 ( 
.A(n_14310),
.B(n_2559),
.Y(n_14432)
);

INVx1_ASAP7_75t_L g14433 ( 
.A(n_14338),
.Y(n_14433)
);

AND2x2_ASAP7_75t_L g14434 ( 
.A(n_14256),
.B(n_2559),
.Y(n_14434)
);

NOR2xp33_ASAP7_75t_L g14435 ( 
.A(n_14272),
.B(n_14306),
.Y(n_14435)
);

AND2x2_ASAP7_75t_L g14436 ( 
.A(n_14276),
.B(n_2560),
.Y(n_14436)
);

HB1xp67_ASAP7_75t_L g14437 ( 
.A(n_14280),
.Y(n_14437)
);

AND2x2_ASAP7_75t_L g14438 ( 
.A(n_14337),
.B(n_2560),
.Y(n_14438)
);

INVx1_ASAP7_75t_L g14439 ( 
.A(n_14356),
.Y(n_14439)
);

INVx2_ASAP7_75t_L g14440 ( 
.A(n_14329),
.Y(n_14440)
);

OR2x2_ASAP7_75t_L g14441 ( 
.A(n_14273),
.B(n_2561),
.Y(n_14441)
);

NOR2xp67_ASAP7_75t_L g14442 ( 
.A(n_14288),
.B(n_2561),
.Y(n_14442)
);

INVx1_ASAP7_75t_L g14443 ( 
.A(n_14318),
.Y(n_14443)
);

INVx1_ASAP7_75t_L g14444 ( 
.A(n_14311),
.Y(n_14444)
);

INVx2_ASAP7_75t_L g14445 ( 
.A(n_14295),
.Y(n_14445)
);

AND2x4_ASAP7_75t_L g14446 ( 
.A(n_14328),
.B(n_2562),
.Y(n_14446)
);

INVx1_ASAP7_75t_L g14447 ( 
.A(n_14316),
.Y(n_14447)
);

INVx2_ASAP7_75t_L g14448 ( 
.A(n_14355),
.Y(n_14448)
);

AND2x2_ASAP7_75t_L g14449 ( 
.A(n_14345),
.B(n_2563),
.Y(n_14449)
);

NAND2xp5_ASAP7_75t_L g14450 ( 
.A(n_14325),
.B(n_2563),
.Y(n_14450)
);

INVx1_ASAP7_75t_L g14451 ( 
.A(n_14330),
.Y(n_14451)
);

AO22x1_ASAP7_75t_L g14452 ( 
.A1(n_14266),
.A2(n_2567),
.B1(n_2564),
.B2(n_2566),
.Y(n_14452)
);

OR2x2_ASAP7_75t_L g14453 ( 
.A(n_14263),
.B(n_2566),
.Y(n_14453)
);

NAND2xp5_ASAP7_75t_L g14454 ( 
.A(n_14331),
.B(n_2567),
.Y(n_14454)
);

INVx1_ASAP7_75t_L g14455 ( 
.A(n_14333),
.Y(n_14455)
);

INVx1_ASAP7_75t_L g14456 ( 
.A(n_14271),
.Y(n_14456)
);

OR2x2_ASAP7_75t_L g14457 ( 
.A(n_14312),
.B(n_2568),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_14358),
.Y(n_14458)
);

INVxp67_ASAP7_75t_SL g14459 ( 
.A(n_14258),
.Y(n_14459)
);

INVx1_ASAP7_75t_L g14460 ( 
.A(n_14339),
.Y(n_14460)
);

NAND2x1p5_ASAP7_75t_L g14461 ( 
.A(n_14270),
.B(n_2568),
.Y(n_14461)
);

NAND2xp5_ASAP7_75t_L g14462 ( 
.A(n_14340),
.B(n_2569),
.Y(n_14462)
);

INVxp67_ASAP7_75t_L g14463 ( 
.A(n_14319),
.Y(n_14463)
);

AO221x1_ASAP7_75t_L g14464 ( 
.A1(n_14315),
.A2(n_2572),
.B1(n_2570),
.B2(n_2571),
.C(n_2573),
.Y(n_14464)
);

NAND2xp5_ASAP7_75t_L g14465 ( 
.A(n_14293),
.B(n_2570),
.Y(n_14465)
);

NOR2xp33_ASAP7_75t_L g14466 ( 
.A(n_14282),
.B(n_2571),
.Y(n_14466)
);

OR2x2_ASAP7_75t_L g14467 ( 
.A(n_14336),
.B(n_2572),
.Y(n_14467)
);

INVx1_ASAP7_75t_L g14468 ( 
.A(n_14351),
.Y(n_14468)
);

INVx1_ASAP7_75t_L g14469 ( 
.A(n_14359),
.Y(n_14469)
);

OR2x2_ASAP7_75t_L g14470 ( 
.A(n_14297),
.B(n_2573),
.Y(n_14470)
);

OR2x2_ASAP7_75t_L g14471 ( 
.A(n_14299),
.B(n_2574),
.Y(n_14471)
);

AND2x4_ASAP7_75t_L g14472 ( 
.A(n_14313),
.B(n_2574),
.Y(n_14472)
);

INVx1_ASAP7_75t_L g14473 ( 
.A(n_14307),
.Y(n_14473)
);

AND2x2_ASAP7_75t_L g14474 ( 
.A(n_14309),
.B(n_2575),
.Y(n_14474)
);

INVx1_ASAP7_75t_L g14475 ( 
.A(n_14327),
.Y(n_14475)
);

INVx1_ASAP7_75t_L g14476 ( 
.A(n_14277),
.Y(n_14476)
);

OR2x6_ASAP7_75t_L g14477 ( 
.A(n_14267),
.B(n_2575),
.Y(n_14477)
);

NOR2xp33_ASAP7_75t_SL g14478 ( 
.A(n_14334),
.B(n_2576),
.Y(n_14478)
);

HB1xp67_ASAP7_75t_L g14479 ( 
.A(n_14300),
.Y(n_14479)
);

NAND2xp5_ASAP7_75t_L g14480 ( 
.A(n_14360),
.B(n_2577),
.Y(n_14480)
);

AND2x2_ASAP7_75t_SL g14481 ( 
.A(n_14343),
.B(n_2577),
.Y(n_14481)
);

INVx1_ASAP7_75t_L g14482 ( 
.A(n_14278),
.Y(n_14482)
);

AND2x2_ASAP7_75t_L g14483 ( 
.A(n_14348),
.B(n_2578),
.Y(n_14483)
);

NAND2xp5_ASAP7_75t_SL g14484 ( 
.A(n_14363),
.B(n_2578),
.Y(n_14484)
);

NAND2xp5_ASAP7_75t_L g14485 ( 
.A(n_14341),
.B(n_2579),
.Y(n_14485)
);

INVx2_ASAP7_75t_SL g14486 ( 
.A(n_14346),
.Y(n_14486)
);

BUFx2_ASAP7_75t_L g14487 ( 
.A(n_14303),
.Y(n_14487)
);

INVx1_ASAP7_75t_L g14488 ( 
.A(n_14294),
.Y(n_14488)
);

INVx3_ASAP7_75t_L g14489 ( 
.A(n_14361),
.Y(n_14489)
);

HB1xp67_ASAP7_75t_L g14490 ( 
.A(n_14344),
.Y(n_14490)
);

OR2x2_ASAP7_75t_L g14491 ( 
.A(n_14324),
.B(n_2579),
.Y(n_14491)
);

AND2x2_ASAP7_75t_L g14492 ( 
.A(n_14354),
.B(n_2580),
.Y(n_14492)
);

INVx2_ASAP7_75t_L g14493 ( 
.A(n_14321),
.Y(n_14493)
);

NOR2x1p5_ASAP7_75t_L g14494 ( 
.A(n_14349),
.B(n_2581),
.Y(n_14494)
);

INVx1_ASAP7_75t_L g14495 ( 
.A(n_14362),
.Y(n_14495)
);

AOI22xp5_ASAP7_75t_L g14496 ( 
.A1(n_14353),
.A2(n_2583),
.B1(n_2581),
.B2(n_2582),
.Y(n_14496)
);

INVx1_ASAP7_75t_L g14497 ( 
.A(n_14296),
.Y(n_14497)
);

NAND2xp5_ASAP7_75t_L g14498 ( 
.A(n_14283),
.B(n_2582),
.Y(n_14498)
);

OR2x2_ASAP7_75t_L g14499 ( 
.A(n_14257),
.B(n_2583),
.Y(n_14499)
);

AND2x2_ASAP7_75t_L g14500 ( 
.A(n_14257),
.B(n_2584),
.Y(n_14500)
);

NAND2xp5_ASAP7_75t_L g14501 ( 
.A(n_14283),
.B(n_2585),
.Y(n_14501)
);

INVxp67_ASAP7_75t_L g14502 ( 
.A(n_14264),
.Y(n_14502)
);

INVx1_ASAP7_75t_L g14503 ( 
.A(n_14257),
.Y(n_14503)
);

AND2x4_ASAP7_75t_SL g14504 ( 
.A(n_14262),
.B(n_2585),
.Y(n_14504)
);

INVx1_ASAP7_75t_L g14505 ( 
.A(n_14257),
.Y(n_14505)
);

INVx1_ASAP7_75t_L g14506 ( 
.A(n_14257),
.Y(n_14506)
);

AND2x2_ASAP7_75t_SL g14507 ( 
.A(n_14283),
.B(n_2586),
.Y(n_14507)
);

INVx1_ASAP7_75t_L g14508 ( 
.A(n_14257),
.Y(n_14508)
);

INVx2_ASAP7_75t_L g14509 ( 
.A(n_14269),
.Y(n_14509)
);

INVx1_ASAP7_75t_L g14510 ( 
.A(n_14257),
.Y(n_14510)
);

NAND2xp5_ASAP7_75t_L g14511 ( 
.A(n_14283),
.B(n_2586),
.Y(n_14511)
);

OR2x2_ASAP7_75t_L g14512 ( 
.A(n_14257),
.B(n_2587),
.Y(n_14512)
);

NAND3xp33_ASAP7_75t_L g14513 ( 
.A(n_14283),
.B(n_2587),
.C(n_2588),
.Y(n_14513)
);

NOR2xp33_ASAP7_75t_L g14514 ( 
.A(n_14283),
.B(n_2589),
.Y(n_14514)
);

INVxp33_ASAP7_75t_L g14515 ( 
.A(n_14264),
.Y(n_14515)
);

AND2x2_ASAP7_75t_L g14516 ( 
.A(n_14257),
.B(n_2589),
.Y(n_14516)
);

OR2x2_ASAP7_75t_L g14517 ( 
.A(n_14257),
.B(n_2590),
.Y(n_14517)
);

INVx1_ASAP7_75t_L g14518 ( 
.A(n_14257),
.Y(n_14518)
);

INVx1_ASAP7_75t_L g14519 ( 
.A(n_14257),
.Y(n_14519)
);

OR2x2_ASAP7_75t_L g14520 ( 
.A(n_14257),
.B(n_2590),
.Y(n_14520)
);

NAND2xp5_ASAP7_75t_L g14521 ( 
.A(n_14283),
.B(n_2591),
.Y(n_14521)
);

AND2x2_ASAP7_75t_L g14522 ( 
.A(n_14257),
.B(n_2592),
.Y(n_14522)
);

OR2x2_ASAP7_75t_L g14523 ( 
.A(n_14257),
.B(n_2592),
.Y(n_14523)
);

INVx2_ASAP7_75t_L g14524 ( 
.A(n_14269),
.Y(n_14524)
);

AND2x4_ASAP7_75t_L g14525 ( 
.A(n_14283),
.B(n_2593),
.Y(n_14525)
);

INVx2_ASAP7_75t_L g14526 ( 
.A(n_14269),
.Y(n_14526)
);

NAND2xp5_ASAP7_75t_L g14527 ( 
.A(n_14283),
.B(n_2593),
.Y(n_14527)
);

INVx1_ASAP7_75t_L g14528 ( 
.A(n_14257),
.Y(n_14528)
);

INVx2_ASAP7_75t_L g14529 ( 
.A(n_14429),
.Y(n_14529)
);

INVx1_ASAP7_75t_L g14530 ( 
.A(n_14417),
.Y(n_14530)
);

INVx2_ASAP7_75t_L g14531 ( 
.A(n_14412),
.Y(n_14531)
);

NAND2xp5_ASAP7_75t_L g14532 ( 
.A(n_14464),
.B(n_2594),
.Y(n_14532)
);

NOR2xp33_ASAP7_75t_L g14533 ( 
.A(n_14515),
.B(n_2594),
.Y(n_14533)
);

INVx1_ASAP7_75t_L g14534 ( 
.A(n_14437),
.Y(n_14534)
);

INVx1_ASAP7_75t_L g14535 ( 
.A(n_14394),
.Y(n_14535)
);

INVx2_ASAP7_75t_L g14536 ( 
.A(n_14461),
.Y(n_14536)
);

AND2x4_ASAP7_75t_L g14537 ( 
.A(n_14379),
.B(n_2595),
.Y(n_14537)
);

BUFx2_ASAP7_75t_L g14538 ( 
.A(n_14502),
.Y(n_14538)
);

OR2x6_ASAP7_75t_L g14539 ( 
.A(n_14498),
.B(n_2595),
.Y(n_14539)
);

AND2x2_ASAP7_75t_L g14540 ( 
.A(n_14382),
.B(n_2596),
.Y(n_14540)
);

INVx2_ASAP7_75t_L g14541 ( 
.A(n_14423),
.Y(n_14541)
);

OR2x2_ASAP7_75t_L g14542 ( 
.A(n_14407),
.B(n_2597),
.Y(n_14542)
);

NAND3xp33_ASAP7_75t_L g14543 ( 
.A(n_14399),
.B(n_2598),
.C(n_2599),
.Y(n_14543)
);

INVx1_ASAP7_75t_L g14544 ( 
.A(n_14423),
.Y(n_14544)
);

OR2x2_ASAP7_75t_L g14545 ( 
.A(n_14415),
.B(n_2598),
.Y(n_14545)
);

OAI322xp33_ASAP7_75t_L g14546 ( 
.A1(n_14463),
.A2(n_2604),
.A3(n_2603),
.B1(n_2601),
.B2(n_2599),
.C1(n_2600),
.C2(n_2602),
.Y(n_14546)
);

INVx1_ASAP7_75t_L g14547 ( 
.A(n_14424),
.Y(n_14547)
);

OR2x2_ASAP7_75t_L g14548 ( 
.A(n_14479),
.B(n_2600),
.Y(n_14548)
);

INVx1_ASAP7_75t_L g14549 ( 
.A(n_14425),
.Y(n_14549)
);

INVx2_ASAP7_75t_L g14550 ( 
.A(n_14494),
.Y(n_14550)
);

AND2x2_ASAP7_75t_L g14551 ( 
.A(n_14419),
.B(n_2601),
.Y(n_14551)
);

NOR2x1_ASAP7_75t_L g14552 ( 
.A(n_14383),
.B(n_2602),
.Y(n_14552)
);

AND2x2_ASAP7_75t_L g14553 ( 
.A(n_14384),
.B(n_2603),
.Y(n_14553)
);

AND2x2_ASAP7_75t_L g14554 ( 
.A(n_14409),
.B(n_14503),
.Y(n_14554)
);

INVx2_ASAP7_75t_L g14555 ( 
.A(n_14507),
.Y(n_14555)
);

INVx1_ASAP7_75t_L g14556 ( 
.A(n_14420),
.Y(n_14556)
);

OAI21xp5_ASAP7_75t_L g14557 ( 
.A1(n_14400),
.A2(n_2605),
.B(n_2606),
.Y(n_14557)
);

INVx1_ASAP7_75t_L g14558 ( 
.A(n_14442),
.Y(n_14558)
);

OR2x2_ASAP7_75t_L g14559 ( 
.A(n_14397),
.B(n_2606),
.Y(n_14559)
);

INVx1_ASAP7_75t_SL g14560 ( 
.A(n_14504),
.Y(n_14560)
);

INVx2_ASAP7_75t_L g14561 ( 
.A(n_14411),
.Y(n_14561)
);

INVx1_ASAP7_75t_SL g14562 ( 
.A(n_14416),
.Y(n_14562)
);

INVx1_ASAP7_75t_L g14563 ( 
.A(n_14474),
.Y(n_14563)
);

INVx1_ASAP7_75t_L g14564 ( 
.A(n_14441),
.Y(n_14564)
);

INVx1_ASAP7_75t_L g14565 ( 
.A(n_14408),
.Y(n_14565)
);

NAND2xp5_ASAP7_75t_L g14566 ( 
.A(n_14452),
.B(n_2607),
.Y(n_14566)
);

OR2x2_ASAP7_75t_L g14567 ( 
.A(n_14458),
.B(n_2607),
.Y(n_14567)
);

INVx2_ASAP7_75t_L g14568 ( 
.A(n_14418),
.Y(n_14568)
);

NAND3xp33_ASAP7_75t_SL g14569 ( 
.A(n_14406),
.B(n_2608),
.C(n_2609),
.Y(n_14569)
);

INVxp67_ASAP7_75t_SL g14570 ( 
.A(n_14398),
.Y(n_14570)
);

INVx1_ASAP7_75t_L g14571 ( 
.A(n_14422),
.Y(n_14571)
);

AND2x2_ASAP7_75t_L g14572 ( 
.A(n_14505),
.B(n_2608),
.Y(n_14572)
);

AOI22xp33_ASAP7_75t_L g14573 ( 
.A1(n_14473),
.A2(n_2612),
.B1(n_2610),
.B2(n_2611),
.Y(n_14573)
);

INVx1_ASAP7_75t_L g14574 ( 
.A(n_14389),
.Y(n_14574)
);

INVx1_ASAP7_75t_L g14575 ( 
.A(n_14405),
.Y(n_14575)
);

NAND2xp5_ASAP7_75t_L g14576 ( 
.A(n_14472),
.B(n_2610),
.Y(n_14576)
);

INVxp67_ASAP7_75t_L g14577 ( 
.A(n_14514),
.Y(n_14577)
);

NAND2xp5_ASAP7_75t_L g14578 ( 
.A(n_14486),
.B(n_14446),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_14396),
.Y(n_14579)
);

INVxp67_ASAP7_75t_SL g14580 ( 
.A(n_14480),
.Y(n_14580)
);

INVx1_ASAP7_75t_L g14581 ( 
.A(n_14500),
.Y(n_14581)
);

INVx2_ASAP7_75t_L g14582 ( 
.A(n_14414),
.Y(n_14582)
);

HB1xp67_ASAP7_75t_L g14583 ( 
.A(n_14477),
.Y(n_14583)
);

OR2x2_ASAP7_75t_L g14584 ( 
.A(n_14506),
.B(n_2611),
.Y(n_14584)
);

INVx1_ASAP7_75t_L g14585 ( 
.A(n_14516),
.Y(n_14585)
);

INVx2_ASAP7_75t_SL g14586 ( 
.A(n_14522),
.Y(n_14586)
);

AND2x2_ASAP7_75t_L g14587 ( 
.A(n_14508),
.B(n_2612),
.Y(n_14587)
);

INVx1_ASAP7_75t_SL g14588 ( 
.A(n_14390),
.Y(n_14588)
);

INVx2_ASAP7_75t_L g14589 ( 
.A(n_14477),
.Y(n_14589)
);

AND2x2_ASAP7_75t_L g14590 ( 
.A(n_14510),
.B(n_2613),
.Y(n_14590)
);

INVx1_ASAP7_75t_L g14591 ( 
.A(n_14470),
.Y(n_14591)
);

NAND2xp5_ASAP7_75t_L g14592 ( 
.A(n_14525),
.B(n_2613),
.Y(n_14592)
);

INVx1_ASAP7_75t_L g14593 ( 
.A(n_14499),
.Y(n_14593)
);

INVx2_ASAP7_75t_SL g14594 ( 
.A(n_14392),
.Y(n_14594)
);

INVx1_ASAP7_75t_L g14595 ( 
.A(n_14512),
.Y(n_14595)
);

AND2x2_ASAP7_75t_L g14596 ( 
.A(n_14518),
.B(n_2614),
.Y(n_14596)
);

INVx1_ASAP7_75t_L g14597 ( 
.A(n_14517),
.Y(n_14597)
);

INVx1_ASAP7_75t_L g14598 ( 
.A(n_14520),
.Y(n_14598)
);

INVx1_ASAP7_75t_L g14599 ( 
.A(n_14523),
.Y(n_14599)
);

INVx1_ASAP7_75t_L g14600 ( 
.A(n_14487),
.Y(n_14600)
);

OAI21xp33_ASAP7_75t_L g14601 ( 
.A1(n_14435),
.A2(n_2614),
.B(n_2615),
.Y(n_14601)
);

INVx2_ASAP7_75t_L g14602 ( 
.A(n_14481),
.Y(n_14602)
);

INVx1_ASAP7_75t_L g14603 ( 
.A(n_14403),
.Y(n_14603)
);

NAND2xp5_ASAP7_75t_L g14604 ( 
.A(n_14388),
.B(n_2616),
.Y(n_14604)
);

OAI21xp5_ASAP7_75t_SL g14605 ( 
.A1(n_14488),
.A2(n_2616),
.B(n_2617),
.Y(n_14605)
);

NAND2xp5_ASAP7_75t_L g14606 ( 
.A(n_14509),
.B(n_2617),
.Y(n_14606)
);

INVx1_ASAP7_75t_L g14607 ( 
.A(n_14483),
.Y(n_14607)
);

INVx1_ASAP7_75t_SL g14608 ( 
.A(n_14391),
.Y(n_14608)
);

INVx1_ASAP7_75t_L g14609 ( 
.A(n_14440),
.Y(n_14609)
);

INVxp67_ASAP7_75t_SL g14610 ( 
.A(n_14395),
.Y(n_14610)
);

INVx1_ASAP7_75t_L g14611 ( 
.A(n_14436),
.Y(n_14611)
);

AND2x2_ASAP7_75t_L g14612 ( 
.A(n_14519),
.B(n_2618),
.Y(n_14612)
);

INVx1_ASAP7_75t_L g14613 ( 
.A(n_14449),
.Y(n_14613)
);

NAND2x1p5_ASAP7_75t_L g14614 ( 
.A(n_14524),
.B(n_2618),
.Y(n_14614)
);

INVx1_ASAP7_75t_L g14615 ( 
.A(n_14492),
.Y(n_14615)
);

AND2x2_ASAP7_75t_L g14616 ( 
.A(n_14528),
.B(n_2619),
.Y(n_14616)
);

INVxp67_ASAP7_75t_SL g14617 ( 
.A(n_14450),
.Y(n_14617)
);

INVx2_ASAP7_75t_L g14618 ( 
.A(n_14448),
.Y(n_14618)
);

INVx1_ASAP7_75t_L g14619 ( 
.A(n_14457),
.Y(n_14619)
);

INVx1_ASAP7_75t_L g14620 ( 
.A(n_14438),
.Y(n_14620)
);

AND2x2_ASAP7_75t_L g14621 ( 
.A(n_14401),
.B(n_2620),
.Y(n_14621)
);

INVx1_ASAP7_75t_L g14622 ( 
.A(n_14386),
.Y(n_14622)
);

OR2x2_ASAP7_75t_L g14623 ( 
.A(n_14385),
.B(n_2620),
.Y(n_14623)
);

INVx1_ASAP7_75t_L g14624 ( 
.A(n_14467),
.Y(n_14624)
);

INVx1_ASAP7_75t_L g14625 ( 
.A(n_14471),
.Y(n_14625)
);

AND2x2_ASAP7_75t_L g14626 ( 
.A(n_14476),
.B(n_2621),
.Y(n_14626)
);

AND2x4_ASAP7_75t_L g14627 ( 
.A(n_14404),
.B(n_2621),
.Y(n_14627)
);

INVx1_ASAP7_75t_L g14628 ( 
.A(n_14490),
.Y(n_14628)
);

NAND2xp5_ASAP7_75t_L g14629 ( 
.A(n_14526),
.B(n_14456),
.Y(n_14629)
);

INVx1_ASAP7_75t_L g14630 ( 
.A(n_14433),
.Y(n_14630)
);

INVx1_ASAP7_75t_L g14631 ( 
.A(n_14430),
.Y(n_14631)
);

INVx1_ASAP7_75t_L g14632 ( 
.A(n_14434),
.Y(n_14632)
);

OR2x2_ASAP7_75t_L g14633 ( 
.A(n_14381),
.B(n_2622),
.Y(n_14633)
);

NAND2xp5_ASAP7_75t_L g14634 ( 
.A(n_14460),
.B(n_2622),
.Y(n_14634)
);

INVx1_ASAP7_75t_L g14635 ( 
.A(n_14491),
.Y(n_14635)
);

INVxp67_ASAP7_75t_L g14636 ( 
.A(n_14466),
.Y(n_14636)
);

INVx1_ASAP7_75t_L g14637 ( 
.A(n_14387),
.Y(n_14637)
);

AND2x2_ASAP7_75t_L g14638 ( 
.A(n_14493),
.B(n_2624),
.Y(n_14638)
);

INVxp67_ASAP7_75t_L g14639 ( 
.A(n_14478),
.Y(n_14639)
);

AND2x4_ASAP7_75t_L g14640 ( 
.A(n_14402),
.B(n_2624),
.Y(n_14640)
);

INVx2_ASAP7_75t_L g14641 ( 
.A(n_14427),
.Y(n_14641)
);

NOR2x1_ASAP7_75t_L g14642 ( 
.A(n_14513),
.B(n_2625),
.Y(n_14642)
);

INVx1_ASAP7_75t_L g14643 ( 
.A(n_14454),
.Y(n_14643)
);

AND2x2_ASAP7_75t_L g14644 ( 
.A(n_14445),
.B(n_2625),
.Y(n_14644)
);

OR2x2_ASAP7_75t_L g14645 ( 
.A(n_14501),
.B(n_2626),
.Y(n_14645)
);

AND2x2_ASAP7_75t_L g14646 ( 
.A(n_14428),
.B(n_2627),
.Y(n_14646)
);

INVx1_ASAP7_75t_L g14647 ( 
.A(n_14462),
.Y(n_14647)
);

OR2x2_ASAP7_75t_L g14648 ( 
.A(n_14511),
.B(n_2628),
.Y(n_14648)
);

INVx1_ASAP7_75t_SL g14649 ( 
.A(n_14453),
.Y(n_14649)
);

INVx1_ASAP7_75t_L g14650 ( 
.A(n_14410),
.Y(n_14650)
);

INVx2_ASAP7_75t_L g14651 ( 
.A(n_14489),
.Y(n_14651)
);

NOR2x1p5_ASAP7_75t_L g14652 ( 
.A(n_14521),
.B(n_2628),
.Y(n_14652)
);

BUFx2_ASAP7_75t_L g14653 ( 
.A(n_14393),
.Y(n_14653)
);

INVx1_ASAP7_75t_SL g14654 ( 
.A(n_14413),
.Y(n_14654)
);

NAND2xp5_ASAP7_75t_L g14655 ( 
.A(n_14459),
.B(n_2629),
.Y(n_14655)
);

AND2x2_ASAP7_75t_L g14656 ( 
.A(n_14447),
.B(n_2629),
.Y(n_14656)
);

INVx1_ASAP7_75t_L g14657 ( 
.A(n_14468),
.Y(n_14657)
);

AOI22xp5_ASAP7_75t_L g14658 ( 
.A1(n_14484),
.A2(n_2633),
.B1(n_2631),
.B2(n_2632),
.Y(n_14658)
);

BUFx3_ASAP7_75t_L g14659 ( 
.A(n_14527),
.Y(n_14659)
);

AND2x2_ASAP7_75t_L g14660 ( 
.A(n_14475),
.B(n_2631),
.Y(n_14660)
);

AND2x2_ASAP7_75t_L g14661 ( 
.A(n_14469),
.B(n_2632),
.Y(n_14661)
);

INVx2_ASAP7_75t_L g14662 ( 
.A(n_14443),
.Y(n_14662)
);

INVx3_ASAP7_75t_L g14663 ( 
.A(n_14497),
.Y(n_14663)
);

OAI21xp33_ASAP7_75t_L g14664 ( 
.A1(n_14495),
.A2(n_2634),
.B(n_2635),
.Y(n_14664)
);

AND2x2_ASAP7_75t_L g14665 ( 
.A(n_14421),
.B(n_2634),
.Y(n_14665)
);

AND2x4_ASAP7_75t_L g14666 ( 
.A(n_14465),
.B(n_2635),
.Y(n_14666)
);

INVx1_ASAP7_75t_L g14667 ( 
.A(n_14432),
.Y(n_14667)
);

NOR2xp33_ASAP7_75t_L g14668 ( 
.A(n_14431),
.B(n_2636),
.Y(n_14668)
);

AND2x2_ASAP7_75t_L g14669 ( 
.A(n_14444),
.B(n_2636),
.Y(n_14669)
);

HB1xp67_ASAP7_75t_L g14670 ( 
.A(n_14439),
.Y(n_14670)
);

INVx1_ASAP7_75t_L g14671 ( 
.A(n_14485),
.Y(n_14671)
);

NAND2xp5_ASAP7_75t_L g14672 ( 
.A(n_14451),
.B(n_2637),
.Y(n_14672)
);

OAI21xp33_ASAP7_75t_L g14673 ( 
.A1(n_14570),
.A2(n_14455),
.B(n_14482),
.Y(n_14673)
);

AOI22xp5_ASAP7_75t_L g14674 ( 
.A1(n_14580),
.A2(n_14496),
.B1(n_14426),
.B2(n_14380),
.Y(n_14674)
);

INVx1_ASAP7_75t_L g14675 ( 
.A(n_14538),
.Y(n_14675)
);

INVx1_ASAP7_75t_L g14676 ( 
.A(n_14554),
.Y(n_14676)
);

OAI211xp5_ASAP7_75t_SL g14677 ( 
.A1(n_14534),
.A2(n_2640),
.B(n_2638),
.C(n_2639),
.Y(n_14677)
);

INVxp67_ASAP7_75t_SL g14678 ( 
.A(n_14552),
.Y(n_14678)
);

INVx1_ASAP7_75t_L g14679 ( 
.A(n_14583),
.Y(n_14679)
);

INVx1_ASAP7_75t_L g14680 ( 
.A(n_14621),
.Y(n_14680)
);

INVx3_ASAP7_75t_L g14681 ( 
.A(n_14537),
.Y(n_14681)
);

NAND2xp5_ASAP7_75t_L g14682 ( 
.A(n_14582),
.B(n_2638),
.Y(n_14682)
);

NOR2x1_ASAP7_75t_L g14683 ( 
.A(n_14531),
.B(n_2639),
.Y(n_14683)
);

OAI22xp33_ASAP7_75t_L g14684 ( 
.A1(n_14548),
.A2(n_2643),
.B1(n_2641),
.B2(n_2642),
.Y(n_14684)
);

NAND3xp33_ASAP7_75t_L g14685 ( 
.A(n_14533),
.B(n_2642),
.C(n_2643),
.Y(n_14685)
);

AOI22xp5_ASAP7_75t_L g14686 ( 
.A1(n_14560),
.A2(n_2646),
.B1(n_2644),
.B2(n_2645),
.Y(n_14686)
);

INVx1_ASAP7_75t_L g14687 ( 
.A(n_14670),
.Y(n_14687)
);

OR2x2_ASAP7_75t_L g14688 ( 
.A(n_14532),
.B(n_2645),
.Y(n_14688)
);

INVx1_ASAP7_75t_L g14689 ( 
.A(n_14553),
.Y(n_14689)
);

AOI211xp5_ASAP7_75t_L g14690 ( 
.A1(n_14530),
.A2(n_2648),
.B(n_2646),
.C(n_2647),
.Y(n_14690)
);

NOR2xp67_ASAP7_75t_SL g14691 ( 
.A(n_14663),
.B(n_2647),
.Y(n_14691)
);

NAND2xp5_ASAP7_75t_L g14692 ( 
.A(n_14627),
.B(n_2648),
.Y(n_14692)
);

OR2x2_ASAP7_75t_L g14693 ( 
.A(n_14653),
.B(n_2649),
.Y(n_14693)
);

O2A1O1Ixp33_ASAP7_75t_L g14694 ( 
.A1(n_14618),
.A2(n_2651),
.B(n_2649),
.C(n_2650),
.Y(n_14694)
);

OA21x2_ASAP7_75t_L g14695 ( 
.A1(n_14557),
.A2(n_2651),
.B(n_2652),
.Y(n_14695)
);

NAND2x1p5_ASAP7_75t_L g14696 ( 
.A(n_14600),
.B(n_2652),
.Y(n_14696)
);

INVx1_ASAP7_75t_L g14697 ( 
.A(n_14559),
.Y(n_14697)
);

NAND2xp5_ASAP7_75t_L g14698 ( 
.A(n_14551),
.B(n_2653),
.Y(n_14698)
);

AOI21xp33_ASAP7_75t_L g14699 ( 
.A1(n_14558),
.A2(n_2653),
.B(n_2654),
.Y(n_14699)
);

AND2x4_ASAP7_75t_L g14700 ( 
.A(n_14651),
.B(n_2654),
.Y(n_14700)
);

INVx1_ASAP7_75t_L g14701 ( 
.A(n_14652),
.Y(n_14701)
);

NAND2xp5_ASAP7_75t_SL g14702 ( 
.A(n_14609),
.B(n_2655),
.Y(n_14702)
);

INVx1_ASAP7_75t_L g14703 ( 
.A(n_14545),
.Y(n_14703)
);

INVx2_ASAP7_75t_SL g14704 ( 
.A(n_14540),
.Y(n_14704)
);

INVx1_ASAP7_75t_L g14705 ( 
.A(n_14623),
.Y(n_14705)
);

INVx2_ASAP7_75t_L g14706 ( 
.A(n_14614),
.Y(n_14706)
);

INVx1_ASAP7_75t_L g14707 ( 
.A(n_14535),
.Y(n_14707)
);

INVx1_ASAP7_75t_L g14708 ( 
.A(n_14566),
.Y(n_14708)
);

INVx1_ASAP7_75t_L g14709 ( 
.A(n_14660),
.Y(n_14709)
);

INVx1_ASAP7_75t_L g14710 ( 
.A(n_14644),
.Y(n_14710)
);

AOI22xp5_ASAP7_75t_L g14711 ( 
.A1(n_14617),
.A2(n_2657),
.B1(n_2655),
.B2(n_2656),
.Y(n_14711)
);

INVx1_ASAP7_75t_L g14712 ( 
.A(n_14556),
.Y(n_14712)
);

NAND2xp5_ASAP7_75t_L g14713 ( 
.A(n_14586),
.B(n_2656),
.Y(n_14713)
);

HB1xp67_ASAP7_75t_L g14714 ( 
.A(n_14539),
.Y(n_14714)
);

AND2x2_ASAP7_75t_L g14715 ( 
.A(n_14662),
.B(n_2657),
.Y(n_14715)
);

INVx1_ASAP7_75t_L g14716 ( 
.A(n_14572),
.Y(n_14716)
);

INVx1_ASAP7_75t_L g14717 ( 
.A(n_14587),
.Y(n_14717)
);

INVx2_ASAP7_75t_L g14718 ( 
.A(n_14539),
.Y(n_14718)
);

AOI222xp33_ASAP7_75t_L g14719 ( 
.A1(n_14562),
.A2(n_2660),
.B1(n_2662),
.B2(n_2658),
.C1(n_2659),
.C2(n_2661),
.Y(n_14719)
);

NAND2xp5_ASAP7_75t_L g14720 ( 
.A(n_14594),
.B(n_2658),
.Y(n_14720)
);

INVx1_ASAP7_75t_L g14721 ( 
.A(n_14590),
.Y(n_14721)
);

A2O1A1Ixp33_ASAP7_75t_L g14722 ( 
.A1(n_14630),
.A2(n_14631),
.B(n_14637),
.C(n_14543),
.Y(n_14722)
);

OR2x2_ASAP7_75t_L g14723 ( 
.A(n_14578),
.B(n_2659),
.Y(n_14723)
);

OR2x2_ASAP7_75t_L g14724 ( 
.A(n_14542),
.B(n_2660),
.Y(n_14724)
);

INVx1_ASAP7_75t_L g14725 ( 
.A(n_14596),
.Y(n_14725)
);

OAI21xp5_ASAP7_75t_L g14726 ( 
.A1(n_14605),
.A2(n_2661),
.B(n_2662),
.Y(n_14726)
);

INVx1_ASAP7_75t_L g14727 ( 
.A(n_14612),
.Y(n_14727)
);

NAND2xp5_ASAP7_75t_L g14728 ( 
.A(n_14640),
.B(n_2663),
.Y(n_14728)
);

AO22x1_ASAP7_75t_L g14729 ( 
.A1(n_14628),
.A2(n_2665),
.B1(n_2663),
.B2(n_2664),
.Y(n_14729)
);

INVx1_ASAP7_75t_SL g14730 ( 
.A(n_14616),
.Y(n_14730)
);

NAND2xp5_ASAP7_75t_L g14731 ( 
.A(n_14588),
.B(n_2664),
.Y(n_14731)
);

INVx2_ASAP7_75t_SL g14732 ( 
.A(n_14626),
.Y(n_14732)
);

OAI21xp33_ASAP7_75t_L g14733 ( 
.A1(n_14629),
.A2(n_2667),
.B(n_2668),
.Y(n_14733)
);

AOI21xp33_ASAP7_75t_SL g14734 ( 
.A1(n_14584),
.A2(n_2667),
.B(n_2668),
.Y(n_14734)
);

INVx1_ASAP7_75t_L g14735 ( 
.A(n_14638),
.Y(n_14735)
);

INVx1_ASAP7_75t_L g14736 ( 
.A(n_14656),
.Y(n_14736)
);

NAND2xp5_ASAP7_75t_L g14737 ( 
.A(n_14610),
.B(n_2669),
.Y(n_14737)
);

INVx1_ASAP7_75t_L g14738 ( 
.A(n_14561),
.Y(n_14738)
);

INVx1_ASAP7_75t_L g14739 ( 
.A(n_14568),
.Y(n_14739)
);

INVx1_ASAP7_75t_L g14740 ( 
.A(n_14661),
.Y(n_14740)
);

AND2x2_ASAP7_75t_L g14741 ( 
.A(n_14657),
.B(n_2669),
.Y(n_14741)
);

AOI21xp33_ASAP7_75t_SL g14742 ( 
.A1(n_14567),
.A2(n_2670),
.B(n_2671),
.Y(n_14742)
);

OR2x2_ASAP7_75t_L g14743 ( 
.A(n_14569),
.B(n_2672),
.Y(n_14743)
);

NAND2xp5_ASAP7_75t_L g14744 ( 
.A(n_14669),
.B(n_2672),
.Y(n_14744)
);

O2A1O1Ixp33_ASAP7_75t_L g14745 ( 
.A1(n_14536),
.A2(n_2676),
.B(n_2673),
.C(n_2675),
.Y(n_14745)
);

A2O1A1Ixp33_ASAP7_75t_L g14746 ( 
.A1(n_14664),
.A2(n_2676),
.B(n_2673),
.C(n_2675),
.Y(n_14746)
);

INVx2_ASAP7_75t_L g14747 ( 
.A(n_14529),
.Y(n_14747)
);

INVx1_ASAP7_75t_L g14748 ( 
.A(n_14576),
.Y(n_14748)
);

A2O1A1Ixp33_ASAP7_75t_L g14749 ( 
.A1(n_14668),
.A2(n_2679),
.B(n_2677),
.C(n_2678),
.Y(n_14749)
);

AND2x2_ASAP7_75t_L g14750 ( 
.A(n_14646),
.B(n_2677),
.Y(n_14750)
);

INVx1_ASAP7_75t_L g14751 ( 
.A(n_14563),
.Y(n_14751)
);

INVx1_ASAP7_75t_L g14752 ( 
.A(n_14547),
.Y(n_14752)
);

INVx1_ASAP7_75t_L g14753 ( 
.A(n_14549),
.Y(n_14753)
);

OR2x2_ASAP7_75t_L g14754 ( 
.A(n_14634),
.B(n_2678),
.Y(n_14754)
);

NAND3xp33_ASAP7_75t_L g14755 ( 
.A(n_14555),
.B(n_2680),
.C(n_2681),
.Y(n_14755)
);

NAND2xp5_ASAP7_75t_SL g14756 ( 
.A(n_14666),
.B(n_2680),
.Y(n_14756)
);

INVx1_ASAP7_75t_L g14757 ( 
.A(n_14592),
.Y(n_14757)
);

INVx1_ASAP7_75t_L g14758 ( 
.A(n_14550),
.Y(n_14758)
);

OAI222xp33_ASAP7_75t_L g14759 ( 
.A1(n_14642),
.A2(n_2683),
.B1(n_2685),
.B2(n_2681),
.C1(n_2682),
.C2(n_2684),
.Y(n_14759)
);

AOI32xp33_ASAP7_75t_L g14760 ( 
.A1(n_14620),
.A2(n_2686),
.A3(n_2682),
.B1(n_2683),
.B2(n_2687),
.Y(n_14760)
);

NAND2xp5_ASAP7_75t_L g14761 ( 
.A(n_14581),
.B(n_2686),
.Y(n_14761)
);

INVx1_ASAP7_75t_L g14762 ( 
.A(n_14602),
.Y(n_14762)
);

INVx1_ASAP7_75t_L g14763 ( 
.A(n_14564),
.Y(n_14763)
);

AOI211xp5_ASAP7_75t_L g14764 ( 
.A1(n_14601),
.A2(n_2689),
.B(n_2687),
.C(n_2688),
.Y(n_14764)
);

INVx1_ASAP7_75t_L g14765 ( 
.A(n_14633),
.Y(n_14765)
);

INVx1_ASAP7_75t_L g14766 ( 
.A(n_14591),
.Y(n_14766)
);

OAI21xp5_ASAP7_75t_L g14767 ( 
.A1(n_14655),
.A2(n_2688),
.B(n_2689),
.Y(n_14767)
);

AND2x4_ASAP7_75t_L g14768 ( 
.A(n_14665),
.B(n_2690),
.Y(n_14768)
);

INVx2_ASAP7_75t_L g14769 ( 
.A(n_14659),
.Y(n_14769)
);

AND2x2_ASAP7_75t_L g14770 ( 
.A(n_14632),
.B(n_2690),
.Y(n_14770)
);

INVx2_ASAP7_75t_L g14771 ( 
.A(n_14645),
.Y(n_14771)
);

INVx1_ASAP7_75t_L g14772 ( 
.A(n_14589),
.Y(n_14772)
);

AND2x4_ASAP7_75t_L g14773 ( 
.A(n_14585),
.B(n_2691),
.Y(n_14773)
);

INVx1_ASAP7_75t_L g14774 ( 
.A(n_14648),
.Y(n_14774)
);

NOR2xp33_ASAP7_75t_L g14775 ( 
.A(n_14611),
.B(n_2692),
.Y(n_14775)
);

INVx2_ASAP7_75t_SL g14776 ( 
.A(n_14604),
.Y(n_14776)
);

OAI22xp5_ASAP7_75t_L g14777 ( 
.A1(n_14658),
.A2(n_2694),
.B1(n_2692),
.B2(n_2693),
.Y(n_14777)
);

NAND2x1_ASAP7_75t_L g14778 ( 
.A(n_14613),
.B(n_2693),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_14593),
.Y(n_14779)
);

OAI22xp5_ASAP7_75t_L g14780 ( 
.A1(n_14573),
.A2(n_2696),
.B1(n_2694),
.B2(n_2695),
.Y(n_14780)
);

INVx1_ASAP7_75t_L g14781 ( 
.A(n_14595),
.Y(n_14781)
);

INVx1_ASAP7_75t_L g14782 ( 
.A(n_14597),
.Y(n_14782)
);

AND2x4_ASAP7_75t_L g14783 ( 
.A(n_14641),
.B(n_2696),
.Y(n_14783)
);

AND2x2_ASAP7_75t_L g14784 ( 
.A(n_14615),
.B(n_14598),
.Y(n_14784)
);

AND2x2_ASAP7_75t_L g14785 ( 
.A(n_14599),
.B(n_2697),
.Y(n_14785)
);

INVx2_ASAP7_75t_L g14786 ( 
.A(n_14635),
.Y(n_14786)
);

NAND3xp33_ASAP7_75t_L g14787 ( 
.A(n_14639),
.B(n_2697),
.C(n_2698),
.Y(n_14787)
);

NAND2xp5_ASAP7_75t_L g14788 ( 
.A(n_14654),
.B(n_2698),
.Y(n_14788)
);

NAND3xp33_ASAP7_75t_L g14789 ( 
.A(n_14650),
.B(n_2699),
.C(n_2700),
.Y(n_14789)
);

INVx1_ASAP7_75t_SL g14790 ( 
.A(n_14672),
.Y(n_14790)
);

INVx2_ASAP7_75t_SL g14791 ( 
.A(n_14606),
.Y(n_14791)
);

OR2x2_ASAP7_75t_L g14792 ( 
.A(n_14608),
.B(n_14622),
.Y(n_14792)
);

NAND2xp5_ASAP7_75t_L g14793 ( 
.A(n_14624),
.B(n_2699),
.Y(n_14793)
);

NOR2xp33_ASAP7_75t_L g14794 ( 
.A(n_14649),
.B(n_2700),
.Y(n_14794)
);

INVxp67_ASAP7_75t_L g14795 ( 
.A(n_14541),
.Y(n_14795)
);

INVx2_ASAP7_75t_L g14796 ( 
.A(n_14619),
.Y(n_14796)
);

INVx2_ASAP7_75t_SL g14797 ( 
.A(n_14625),
.Y(n_14797)
);

NAND2xp5_ASAP7_75t_L g14798 ( 
.A(n_14565),
.B(n_14571),
.Y(n_14798)
);

INVx2_ASAP7_75t_L g14799 ( 
.A(n_14607),
.Y(n_14799)
);

OAI32xp33_ASAP7_75t_L g14800 ( 
.A1(n_14671),
.A2(n_2703),
.A3(n_2701),
.B1(n_2702),
.B2(n_2704),
.Y(n_14800)
);

INVx1_ASAP7_75t_L g14801 ( 
.A(n_14544),
.Y(n_14801)
);

INVx1_ASAP7_75t_L g14802 ( 
.A(n_14574),
.Y(n_14802)
);

AOI21x1_ASAP7_75t_L g14803 ( 
.A1(n_14643),
.A2(n_2702),
.B(n_2703),
.Y(n_14803)
);

AND2x2_ASAP7_75t_L g14804 ( 
.A(n_14647),
.B(n_2704),
.Y(n_14804)
);

INVx1_ASAP7_75t_L g14805 ( 
.A(n_14575),
.Y(n_14805)
);

INVx1_ASAP7_75t_L g14806 ( 
.A(n_14579),
.Y(n_14806)
);

OR2x2_ASAP7_75t_L g14807 ( 
.A(n_14603),
.B(n_2705),
.Y(n_14807)
);

INVx1_ASAP7_75t_L g14808 ( 
.A(n_14546),
.Y(n_14808)
);

O2A1O1Ixp33_ASAP7_75t_L g14809 ( 
.A1(n_14675),
.A2(n_14636),
.B(n_14577),
.C(n_14667),
.Y(n_14809)
);

INVx2_ASAP7_75t_L g14810 ( 
.A(n_14696),
.Y(n_14810)
);

NOR2xp67_ASAP7_75t_SL g14811 ( 
.A(n_14714),
.B(n_2705),
.Y(n_14811)
);

OR2x2_ASAP7_75t_L g14812 ( 
.A(n_14693),
.B(n_2706),
.Y(n_14812)
);

NAND2xp5_ASAP7_75t_SL g14813 ( 
.A(n_14687),
.B(n_2706),
.Y(n_14813)
);

AND2x2_ASAP7_75t_L g14814 ( 
.A(n_14676),
.B(n_2707),
.Y(n_14814)
);

OR2x2_ASAP7_75t_L g14815 ( 
.A(n_14681),
.B(n_2707),
.Y(n_14815)
);

INVx2_ASAP7_75t_L g14816 ( 
.A(n_14803),
.Y(n_14816)
);

NAND2xp5_ASAP7_75t_L g14817 ( 
.A(n_14729),
.B(n_2708),
.Y(n_14817)
);

BUFx2_ASAP7_75t_L g14818 ( 
.A(n_14678),
.Y(n_14818)
);

AND2x4_ASAP7_75t_L g14819 ( 
.A(n_14797),
.B(n_2708),
.Y(n_14819)
);

AOI31xp33_ASAP7_75t_L g14820 ( 
.A1(n_14769),
.A2(n_2711),
.A3(n_2709),
.B(n_2710),
.Y(n_14820)
);

AND2x2_ASAP7_75t_L g14821 ( 
.A(n_14712),
.B(n_2709),
.Y(n_14821)
);

NOR4xp25_ASAP7_75t_L g14822 ( 
.A(n_14673),
.B(n_2712),
.C(n_2710),
.D(n_2711),
.Y(n_14822)
);

NAND2xp5_ASAP7_75t_L g14823 ( 
.A(n_14750),
.B(n_2712),
.Y(n_14823)
);

OR2x2_ASAP7_75t_L g14824 ( 
.A(n_14778),
.B(n_2713),
.Y(n_14824)
);

INVxp67_ASAP7_75t_L g14825 ( 
.A(n_14691),
.Y(n_14825)
);

AOI221xp5_ASAP7_75t_L g14826 ( 
.A1(n_14762),
.A2(n_2715),
.B1(n_2713),
.B2(n_2714),
.C(n_2716),
.Y(n_14826)
);

INVx1_ASAP7_75t_L g14827 ( 
.A(n_14683),
.Y(n_14827)
);

INVx1_ASAP7_75t_L g14828 ( 
.A(n_14724),
.Y(n_14828)
);

OAI22xp5_ASAP7_75t_L g14829 ( 
.A1(n_14722),
.A2(n_2717),
.B1(n_2715),
.B2(n_2716),
.Y(n_14829)
);

INVx2_ASAP7_75t_L g14830 ( 
.A(n_14783),
.Y(n_14830)
);

NOR2xp33_ASAP7_75t_L g14831 ( 
.A(n_14759),
.B(n_2717),
.Y(n_14831)
);

INVx1_ASAP7_75t_L g14832 ( 
.A(n_14743),
.Y(n_14832)
);

INVx1_ASAP7_75t_L g14833 ( 
.A(n_14698),
.Y(n_14833)
);

NAND2xp5_ASAP7_75t_L g14834 ( 
.A(n_14700),
.B(n_2718),
.Y(n_14834)
);

INVx1_ASAP7_75t_SL g14835 ( 
.A(n_14792),
.Y(n_14835)
);

CKINVDCx20_ASAP7_75t_R g14836 ( 
.A(n_14730),
.Y(n_14836)
);

NOR2xp33_ASAP7_75t_SL g14837 ( 
.A(n_14738),
.B(n_2719),
.Y(n_14837)
);

NAND2xp5_ASAP7_75t_L g14838 ( 
.A(n_14768),
.B(n_2719),
.Y(n_14838)
);

AOI22xp5_ASAP7_75t_L g14839 ( 
.A1(n_14708),
.A2(n_2722),
.B1(n_2720),
.B2(n_2721),
.Y(n_14839)
);

NAND4xp25_ASAP7_75t_SL g14840 ( 
.A(n_14751),
.B(n_2723),
.C(n_2720),
.D(n_2722),
.Y(n_14840)
);

NOR2xp33_ASAP7_75t_L g14841 ( 
.A(n_14677),
.B(n_2724),
.Y(n_14841)
);

INVx1_ASAP7_75t_L g14842 ( 
.A(n_14741),
.Y(n_14842)
);

INVx1_ASAP7_75t_L g14843 ( 
.A(n_14715),
.Y(n_14843)
);

AOI22xp5_ASAP7_75t_L g14844 ( 
.A1(n_14779),
.A2(n_2728),
.B1(n_2726),
.B2(n_2727),
.Y(n_14844)
);

INVx1_ASAP7_75t_L g14845 ( 
.A(n_14785),
.Y(n_14845)
);

INVx1_ASAP7_75t_L g14846 ( 
.A(n_14744),
.Y(n_14846)
);

INVxp67_ASAP7_75t_L g14847 ( 
.A(n_14794),
.Y(n_14847)
);

INVx1_ASAP7_75t_L g14848 ( 
.A(n_14770),
.Y(n_14848)
);

INVx2_ASAP7_75t_L g14849 ( 
.A(n_14695),
.Y(n_14849)
);

AOI31xp33_ASAP7_75t_SL g14850 ( 
.A1(n_14799),
.A2(n_14798),
.A3(n_14786),
.B(n_14796),
.Y(n_14850)
);

NOR2xp67_ASAP7_75t_L g14851 ( 
.A(n_14686),
.B(n_2727),
.Y(n_14851)
);

INVx2_ASAP7_75t_L g14852 ( 
.A(n_14695),
.Y(n_14852)
);

INVx1_ASAP7_75t_L g14853 ( 
.A(n_14728),
.Y(n_14853)
);

AOI322xp5_ASAP7_75t_L g14854 ( 
.A1(n_14790),
.A2(n_2733),
.A3(n_2732),
.B1(n_2730),
.B2(n_2728),
.C1(n_2729),
.C2(n_2731),
.Y(n_14854)
);

AOI32xp33_ASAP7_75t_L g14855 ( 
.A1(n_14752),
.A2(n_2732),
.A3(n_2730),
.B1(n_2731),
.B2(n_2734),
.Y(n_14855)
);

INVx2_ASAP7_75t_L g14856 ( 
.A(n_14807),
.Y(n_14856)
);

AND2x4_ASAP7_75t_L g14857 ( 
.A(n_14739),
.B(n_2735),
.Y(n_14857)
);

INVx1_ASAP7_75t_L g14858 ( 
.A(n_14804),
.Y(n_14858)
);

AOI21xp33_ASAP7_75t_L g14859 ( 
.A1(n_14701),
.A2(n_2735),
.B(n_2736),
.Y(n_14859)
);

INVx1_ASAP7_75t_L g14860 ( 
.A(n_14680),
.Y(n_14860)
);

AOI211xp5_ASAP7_75t_L g14861 ( 
.A1(n_14753),
.A2(n_2738),
.B(n_2736),
.C(n_2737),
.Y(n_14861)
);

AOI22xp5_ASAP7_75t_L g14862 ( 
.A1(n_14781),
.A2(n_2739),
.B1(n_2737),
.B2(n_2738),
.Y(n_14862)
);

A2O1A1Ixp33_ASAP7_75t_L g14863 ( 
.A1(n_14694),
.A2(n_2742),
.B(n_2740),
.C(n_2741),
.Y(n_14863)
);

AOI22x1_ASAP7_75t_L g14864 ( 
.A1(n_14802),
.A2(n_2743),
.B1(n_2740),
.B2(n_2742),
.Y(n_14864)
);

OAI21xp33_ASAP7_75t_L g14865 ( 
.A1(n_14758),
.A2(n_14784),
.B(n_14679),
.Y(n_14865)
);

INVx1_ASAP7_75t_L g14866 ( 
.A(n_14689),
.Y(n_14866)
);

INVx1_ASAP7_75t_L g14867 ( 
.A(n_14692),
.Y(n_14867)
);

INVx2_ASAP7_75t_L g14868 ( 
.A(n_14706),
.Y(n_14868)
);

INVx2_ASAP7_75t_L g14869 ( 
.A(n_14773),
.Y(n_14869)
);

INVx1_ASAP7_75t_L g14870 ( 
.A(n_14705),
.Y(n_14870)
);

INVx1_ASAP7_75t_SL g14871 ( 
.A(n_14723),
.Y(n_14871)
);

INVx2_ASAP7_75t_L g14872 ( 
.A(n_14732),
.Y(n_14872)
);

NAND2xp5_ASAP7_75t_L g14873 ( 
.A(n_14704),
.B(n_2743),
.Y(n_14873)
);

NAND2xp5_ASAP7_75t_L g14874 ( 
.A(n_14740),
.B(n_2744),
.Y(n_14874)
);

INVx1_ASAP7_75t_L g14875 ( 
.A(n_14697),
.Y(n_14875)
);

INVx1_ASAP7_75t_L g14876 ( 
.A(n_14703),
.Y(n_14876)
);

INVx1_ASAP7_75t_L g14877 ( 
.A(n_14754),
.Y(n_14877)
);

AOI22xp5_ASAP7_75t_L g14878 ( 
.A1(n_14782),
.A2(n_2747),
.B1(n_2745),
.B2(n_2746),
.Y(n_14878)
);

OAI32xp33_ASAP7_75t_L g14879 ( 
.A1(n_14763),
.A2(n_14766),
.A3(n_14806),
.B1(n_14805),
.B2(n_14808),
.Y(n_14879)
);

OAI21xp5_ASAP7_75t_L g14880 ( 
.A1(n_14726),
.A2(n_2745),
.B(n_2746),
.Y(n_14880)
);

INVx2_ASAP7_75t_L g14881 ( 
.A(n_14771),
.Y(n_14881)
);

INVx1_ASAP7_75t_L g14882 ( 
.A(n_14718),
.Y(n_14882)
);

AOI21xp5_ASAP7_75t_L g14883 ( 
.A1(n_14702),
.A2(n_2747),
.B(n_2748),
.Y(n_14883)
);

NAND2xp5_ASAP7_75t_L g14884 ( 
.A(n_14734),
.B(n_14742),
.Y(n_14884)
);

INVx1_ASAP7_75t_L g14885 ( 
.A(n_14737),
.Y(n_14885)
);

INVx1_ASAP7_75t_L g14886 ( 
.A(n_14756),
.Y(n_14886)
);

NOR2x1_ASAP7_75t_L g14887 ( 
.A(n_14787),
.B(n_2748),
.Y(n_14887)
);

NAND2xp5_ASAP7_75t_L g14888 ( 
.A(n_14716),
.B(n_2749),
.Y(n_14888)
);

INVx1_ASAP7_75t_L g14889 ( 
.A(n_14788),
.Y(n_14889)
);

INVx1_ASAP7_75t_SL g14890 ( 
.A(n_14688),
.Y(n_14890)
);

INVx2_ASAP7_75t_SL g14891 ( 
.A(n_14747),
.Y(n_14891)
);

INVx1_ASAP7_75t_L g14892 ( 
.A(n_14710),
.Y(n_14892)
);

NAND2xp5_ASAP7_75t_L g14893 ( 
.A(n_14717),
.B(n_2749),
.Y(n_14893)
);

NOR2x1_ASAP7_75t_L g14894 ( 
.A(n_14789),
.B(n_14755),
.Y(n_14894)
);

OR2x2_ASAP7_75t_L g14895 ( 
.A(n_14713),
.B(n_2750),
.Y(n_14895)
);

INVx2_ASAP7_75t_L g14896 ( 
.A(n_14765),
.Y(n_14896)
);

INVx1_ASAP7_75t_L g14897 ( 
.A(n_14709),
.Y(n_14897)
);

AOI21xp5_ASAP7_75t_L g14898 ( 
.A1(n_14746),
.A2(n_2751),
.B(n_2752),
.Y(n_14898)
);

OAI32xp33_ASAP7_75t_L g14899 ( 
.A1(n_14682),
.A2(n_2754),
.A3(n_2751),
.B1(n_2753),
.B2(n_2755),
.Y(n_14899)
);

NOR2xp33_ASAP7_75t_L g14900 ( 
.A(n_14721),
.B(n_2754),
.Y(n_14900)
);

INVxp67_ASAP7_75t_L g14901 ( 
.A(n_14775),
.Y(n_14901)
);

INVx1_ASAP7_75t_SL g14902 ( 
.A(n_14731),
.Y(n_14902)
);

OAI32xp33_ASAP7_75t_L g14903 ( 
.A1(n_14707),
.A2(n_2757),
.A3(n_2755),
.B1(n_2756),
.B2(n_2758),
.Y(n_14903)
);

INVx1_ASAP7_75t_L g14904 ( 
.A(n_14774),
.Y(n_14904)
);

INVxp67_ASAP7_75t_L g14905 ( 
.A(n_14736),
.Y(n_14905)
);

INVxp67_ASAP7_75t_L g14906 ( 
.A(n_14725),
.Y(n_14906)
);

INVx1_ASAP7_75t_L g14907 ( 
.A(n_14727),
.Y(n_14907)
);

INVx1_ASAP7_75t_SL g14908 ( 
.A(n_14793),
.Y(n_14908)
);

O2A1O1Ixp33_ASAP7_75t_L g14909 ( 
.A1(n_14720),
.A2(n_2760),
.B(n_2756),
.C(n_2759),
.Y(n_14909)
);

OAI21xp33_ASAP7_75t_L g14910 ( 
.A1(n_14674),
.A2(n_2759),
.B(n_2760),
.Y(n_14910)
);

NAND2xp5_ASAP7_75t_SL g14911 ( 
.A(n_14719),
.B(n_2761),
.Y(n_14911)
);

OAI21xp5_ASAP7_75t_L g14912 ( 
.A1(n_14745),
.A2(n_2761),
.B(n_2762),
.Y(n_14912)
);

HB1xp67_ASAP7_75t_L g14913 ( 
.A(n_14795),
.Y(n_14913)
);

INVx2_ASAP7_75t_L g14914 ( 
.A(n_14776),
.Y(n_14914)
);

HB1xp67_ASAP7_75t_L g14915 ( 
.A(n_14735),
.Y(n_14915)
);

OAI211xp5_ASAP7_75t_SL g14916 ( 
.A1(n_14801),
.A2(n_2764),
.B(n_2762),
.C(n_2763),
.Y(n_14916)
);

NAND2x1_ASAP7_75t_L g14917 ( 
.A(n_14761),
.B(n_2763),
.Y(n_14917)
);

A2O1A1Ixp33_ASAP7_75t_L g14918 ( 
.A1(n_14733),
.A2(n_2766),
.B(n_2764),
.C(n_2765),
.Y(n_14918)
);

INVx1_ASAP7_75t_L g14919 ( 
.A(n_14772),
.Y(n_14919)
);

OAI22xp5_ASAP7_75t_L g14920 ( 
.A1(n_14711),
.A2(n_2768),
.B1(n_2765),
.B2(n_2767),
.Y(n_14920)
);

INVx1_ASAP7_75t_L g14921 ( 
.A(n_14791),
.Y(n_14921)
);

NAND3xp33_ASAP7_75t_L g14922 ( 
.A(n_14685),
.B(n_2767),
.C(n_2768),
.Y(n_14922)
);

INVx2_ASAP7_75t_L g14923 ( 
.A(n_14757),
.Y(n_14923)
);

NAND2xp5_ASAP7_75t_L g14924 ( 
.A(n_14690),
.B(n_14760),
.Y(n_14924)
);

OAI33xp33_ASAP7_75t_L g14925 ( 
.A1(n_14748),
.A2(n_2771),
.A3(n_2773),
.B1(n_2769),
.B2(n_2770),
.B3(n_2772),
.Y(n_14925)
);

NAND2xp5_ASAP7_75t_L g14926 ( 
.A(n_14749),
.B(n_2769),
.Y(n_14926)
);

AOI21xp5_ASAP7_75t_SL g14927 ( 
.A1(n_14767),
.A2(n_2770),
.B(n_2772),
.Y(n_14927)
);

NAND2xp5_ASAP7_75t_L g14928 ( 
.A(n_14684),
.B(n_2773),
.Y(n_14928)
);

AND2x2_ASAP7_75t_L g14929 ( 
.A(n_14764),
.B(n_2774),
.Y(n_14929)
);

NOR3xp33_ASAP7_75t_L g14930 ( 
.A(n_14699),
.B(n_2775),
.C(n_2776),
.Y(n_14930)
);

AOI21xp5_ASAP7_75t_L g14931 ( 
.A1(n_14777),
.A2(n_2775),
.B(n_2776),
.Y(n_14931)
);

AOI21xp5_ASAP7_75t_L g14932 ( 
.A1(n_14800),
.A2(n_2777),
.B(n_2778),
.Y(n_14932)
);

AND2x2_ASAP7_75t_L g14933 ( 
.A(n_14780),
.B(n_2779),
.Y(n_14933)
);

AND2x4_ASAP7_75t_SL g14934 ( 
.A(n_14769),
.B(n_2779),
.Y(n_14934)
);

OAI22xp5_ASAP7_75t_L g14935 ( 
.A1(n_14835),
.A2(n_2782),
.B1(n_2780),
.B2(n_2781),
.Y(n_14935)
);

OAI221xp5_ASAP7_75t_L g14936 ( 
.A1(n_14818),
.A2(n_2783),
.B1(n_2780),
.B2(n_2781),
.C(n_2784),
.Y(n_14936)
);

AOI21xp5_ASAP7_75t_SL g14937 ( 
.A1(n_14865),
.A2(n_2783),
.B(n_2784),
.Y(n_14937)
);

INVx1_ASAP7_75t_L g14938 ( 
.A(n_14913),
.Y(n_14938)
);

O2A1O1Ixp33_ASAP7_75t_L g14939 ( 
.A1(n_14850),
.A2(n_2787),
.B(n_2785),
.C(n_2786),
.Y(n_14939)
);

OAI21xp33_ASAP7_75t_L g14940 ( 
.A1(n_14891),
.A2(n_2786),
.B(n_2787),
.Y(n_14940)
);

NAND2xp33_ASAP7_75t_L g14941 ( 
.A(n_14836),
.B(n_14921),
.Y(n_14941)
);

INVx1_ASAP7_75t_L g14942 ( 
.A(n_14819),
.Y(n_14942)
);

NOR2xp33_ASAP7_75t_L g14943 ( 
.A(n_14827),
.B(n_2788),
.Y(n_14943)
);

INVx2_ASAP7_75t_L g14944 ( 
.A(n_14824),
.Y(n_14944)
);

AOI21xp33_ASAP7_75t_L g14945 ( 
.A1(n_14816),
.A2(n_2788),
.B(n_2789),
.Y(n_14945)
);

INVx1_ASAP7_75t_L g14946 ( 
.A(n_14819),
.Y(n_14946)
);

OA33x2_ASAP7_75t_L g14947 ( 
.A1(n_14924),
.A2(n_2791),
.A3(n_2793),
.B1(n_2789),
.B2(n_2790),
.B3(n_2792),
.Y(n_14947)
);

INVx1_ASAP7_75t_L g14948 ( 
.A(n_14849),
.Y(n_14948)
);

OAI22xp5_ASAP7_75t_L g14949 ( 
.A1(n_14825),
.A2(n_2793),
.B1(n_2790),
.B2(n_2792),
.Y(n_14949)
);

A2O1A1Ixp33_ASAP7_75t_L g14950 ( 
.A1(n_14915),
.A2(n_2796),
.B(n_2794),
.C(n_2795),
.Y(n_14950)
);

AOI32xp33_ASAP7_75t_L g14951 ( 
.A1(n_14872),
.A2(n_2796),
.A3(n_2794),
.B1(n_2795),
.B2(n_2797),
.Y(n_14951)
);

OA21x2_ASAP7_75t_L g14952 ( 
.A1(n_14873),
.A2(n_2798),
.B(n_2799),
.Y(n_14952)
);

XOR2x2_ASAP7_75t_L g14953 ( 
.A(n_14917),
.B(n_2798),
.Y(n_14953)
);

INVx1_ASAP7_75t_L g14954 ( 
.A(n_14852),
.Y(n_14954)
);

INVx1_ASAP7_75t_SL g14955 ( 
.A(n_14934),
.Y(n_14955)
);

OAI32xp33_ASAP7_75t_L g14956 ( 
.A1(n_14860),
.A2(n_2803),
.A3(n_2799),
.B1(n_2800),
.B2(n_2804),
.Y(n_14956)
);

INVx1_ASAP7_75t_SL g14957 ( 
.A(n_14812),
.Y(n_14957)
);

OAI21xp5_ASAP7_75t_L g14958 ( 
.A1(n_14905),
.A2(n_2803),
.B(n_2805),
.Y(n_14958)
);

NAND2xp5_ASAP7_75t_L g14959 ( 
.A(n_14871),
.B(n_14822),
.Y(n_14959)
);

OAI22xp5_ASAP7_75t_L g14960 ( 
.A1(n_14906),
.A2(n_2808),
.B1(n_2806),
.B2(n_2807),
.Y(n_14960)
);

AOI211xp5_ASAP7_75t_L g14961 ( 
.A1(n_14879),
.A2(n_2811),
.B(n_2809),
.C(n_2810),
.Y(n_14961)
);

AOI22xp5_ASAP7_75t_L g14962 ( 
.A1(n_14866),
.A2(n_2812),
.B1(n_2809),
.B2(n_2810),
.Y(n_14962)
);

INVx1_ASAP7_75t_L g14963 ( 
.A(n_14919),
.Y(n_14963)
);

INVx1_ASAP7_75t_L g14964 ( 
.A(n_14857),
.Y(n_14964)
);

AOI21xp33_ASAP7_75t_L g14965 ( 
.A1(n_14890),
.A2(n_2812),
.B(n_2813),
.Y(n_14965)
);

AOI22xp5_ASAP7_75t_L g14966 ( 
.A1(n_14897),
.A2(n_2815),
.B1(n_2813),
.B2(n_2814),
.Y(n_14966)
);

OAI221xp5_ASAP7_75t_L g14967 ( 
.A1(n_14907),
.A2(n_2817),
.B1(n_2815),
.B2(n_2816),
.C(n_2818),
.Y(n_14967)
);

INVx1_ASAP7_75t_L g14968 ( 
.A(n_14857),
.Y(n_14968)
);

AOI22xp5_ASAP7_75t_L g14969 ( 
.A1(n_14892),
.A2(n_2819),
.B1(n_2816),
.B2(n_2817),
.Y(n_14969)
);

XNOR2x1_ASAP7_75t_L g14970 ( 
.A(n_14894),
.B(n_2820),
.Y(n_14970)
);

AOI22xp5_ASAP7_75t_L g14971 ( 
.A1(n_14870),
.A2(n_14875),
.B1(n_14876),
.B2(n_14851),
.Y(n_14971)
);

HB1xp67_ASAP7_75t_L g14972 ( 
.A(n_14881),
.Y(n_14972)
);

INVx2_ASAP7_75t_L g14973 ( 
.A(n_14864),
.Y(n_14973)
);

OAI211xp5_ASAP7_75t_L g14974 ( 
.A1(n_14809),
.A2(n_2822),
.B(n_2820),
.C(n_2821),
.Y(n_14974)
);

O2A1O1Ixp33_ASAP7_75t_L g14975 ( 
.A1(n_14813),
.A2(n_2824),
.B(n_2821),
.C(n_2823),
.Y(n_14975)
);

O2A1O1Ixp33_ASAP7_75t_L g14976 ( 
.A1(n_14829),
.A2(n_2825),
.B(n_2823),
.C(n_2824),
.Y(n_14976)
);

AOI21xp33_ASAP7_75t_SL g14977 ( 
.A1(n_14820),
.A2(n_2825),
.B(n_2826),
.Y(n_14977)
);

AOI22xp5_ASAP7_75t_L g14978 ( 
.A1(n_14810),
.A2(n_2828),
.B1(n_2826),
.B2(n_2827),
.Y(n_14978)
);

AND2x2_ASAP7_75t_L g14979 ( 
.A(n_14814),
.B(n_2828),
.Y(n_14979)
);

INVx1_ASAP7_75t_L g14980 ( 
.A(n_14823),
.Y(n_14980)
);

NAND3xp33_ASAP7_75t_L g14981 ( 
.A(n_14811),
.B(n_2829),
.C(n_2830),
.Y(n_14981)
);

NAND2xp5_ASAP7_75t_L g14982 ( 
.A(n_14908),
.B(n_2829),
.Y(n_14982)
);

HB1xp67_ASAP7_75t_L g14983 ( 
.A(n_14840),
.Y(n_14983)
);

INVxp67_ASAP7_75t_SL g14984 ( 
.A(n_14817),
.Y(n_14984)
);

INVx1_ASAP7_75t_L g14985 ( 
.A(n_14821),
.Y(n_14985)
);

INVx2_ASAP7_75t_L g14986 ( 
.A(n_14815),
.Y(n_14986)
);

AOI22xp5_ASAP7_75t_L g14987 ( 
.A1(n_14904),
.A2(n_2834),
.B1(n_2831),
.B2(n_2833),
.Y(n_14987)
);

AOI22xp5_ASAP7_75t_SL g14988 ( 
.A1(n_14831),
.A2(n_2835),
.B1(n_2831),
.B2(n_2833),
.Y(n_14988)
);

AOI22xp5_ASAP7_75t_L g14989 ( 
.A1(n_14911),
.A2(n_2837),
.B1(n_2835),
.B2(n_2836),
.Y(n_14989)
);

INVxp67_ASAP7_75t_L g14990 ( 
.A(n_14837),
.Y(n_14990)
);

NAND4xp25_ASAP7_75t_L g14991 ( 
.A(n_14896),
.B(n_2839),
.C(n_2836),
.D(n_2838),
.Y(n_14991)
);

NAND2xp5_ASAP7_75t_L g14992 ( 
.A(n_14848),
.B(n_2838),
.Y(n_14992)
);

INVx2_ASAP7_75t_L g14993 ( 
.A(n_14856),
.Y(n_14993)
);

OAI21xp5_ASAP7_75t_L g14994 ( 
.A1(n_14932),
.A2(n_14883),
.B(n_14898),
.Y(n_14994)
);

AOI22xp5_ASAP7_75t_L g14995 ( 
.A1(n_14902),
.A2(n_2841),
.B1(n_2839),
.B2(n_2840),
.Y(n_14995)
);

INVx2_ASAP7_75t_L g14996 ( 
.A(n_14830),
.Y(n_14996)
);

OAI22xp5_ASAP7_75t_L g14997 ( 
.A1(n_14923),
.A2(n_2843),
.B1(n_2841),
.B2(n_2842),
.Y(n_14997)
);

AOI22xp33_ASAP7_75t_L g14998 ( 
.A1(n_14885),
.A2(n_2845),
.B1(n_2843),
.B2(n_2844),
.Y(n_14998)
);

AOI22xp5_ASAP7_75t_L g14999 ( 
.A1(n_14832),
.A2(n_2847),
.B1(n_2845),
.B2(n_2846),
.Y(n_14999)
);

NAND3xp33_ASAP7_75t_L g15000 ( 
.A(n_14882),
.B(n_2846),
.C(n_2847),
.Y(n_15000)
);

O2A1O1Ixp33_ASAP7_75t_L g15001 ( 
.A1(n_14914),
.A2(n_2850),
.B(n_2848),
.C(n_2849),
.Y(n_15001)
);

NOR4xp25_ASAP7_75t_L g15002 ( 
.A(n_14868),
.B(n_14886),
.C(n_14847),
.D(n_14901),
.Y(n_15002)
);

NAND2x1_ASAP7_75t_SL g15003 ( 
.A(n_14839),
.B(n_2848),
.Y(n_15003)
);

NAND2xp5_ASAP7_75t_L g15004 ( 
.A(n_14869),
.B(n_2850),
.Y(n_15004)
);

INVxp67_ASAP7_75t_L g15005 ( 
.A(n_14841),
.Y(n_15005)
);

OAI21xp5_ASAP7_75t_L g15006 ( 
.A1(n_14863),
.A2(n_2851),
.B(n_2852),
.Y(n_15006)
);

AOI211xp5_ASAP7_75t_SL g15007 ( 
.A1(n_14927),
.A2(n_2855),
.B(n_2853),
.C(n_2854),
.Y(n_15007)
);

NAND2xp5_ASAP7_75t_L g15008 ( 
.A(n_14858),
.B(n_2853),
.Y(n_15008)
);

INVx1_ASAP7_75t_L g15009 ( 
.A(n_14884),
.Y(n_15009)
);

AOI22xp5_ASAP7_75t_L g15010 ( 
.A1(n_14867),
.A2(n_2857),
.B1(n_2854),
.B2(n_2856),
.Y(n_15010)
);

NOR2xp33_ASAP7_75t_L g15011 ( 
.A(n_14925),
.B(n_2857),
.Y(n_15011)
);

OAI22xp33_ASAP7_75t_L g15012 ( 
.A1(n_14874),
.A2(n_14893),
.B1(n_14888),
.B2(n_14895),
.Y(n_15012)
);

AOI322xp5_ASAP7_75t_L g15013 ( 
.A1(n_14887),
.A2(n_2864),
.A3(n_2863),
.B1(n_2861),
.B2(n_2858),
.C1(n_2860),
.C2(n_2862),
.Y(n_15013)
);

OAI21xp5_ASAP7_75t_L g15014 ( 
.A1(n_14931),
.A2(n_2858),
.B(n_2860),
.Y(n_15014)
);

NAND2x1_ASAP7_75t_L g15015 ( 
.A(n_14929),
.B(n_2862),
.Y(n_15015)
);

OAI22xp33_ASAP7_75t_L g15016 ( 
.A1(n_14844),
.A2(n_2865),
.B1(n_2863),
.B2(n_2864),
.Y(n_15016)
);

OAI21xp5_ASAP7_75t_L g15017 ( 
.A1(n_14922),
.A2(n_2865),
.B(n_2866),
.Y(n_15017)
);

NAND2xp5_ASAP7_75t_L g15018 ( 
.A(n_14842),
.B(n_2866),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14834),
.Y(n_15019)
);

AOI222xp33_ASAP7_75t_L g15020 ( 
.A1(n_14877),
.A2(n_2869),
.B1(n_2871),
.B2(n_2867),
.C1(n_2868),
.C2(n_2870),
.Y(n_15020)
);

OAI31xp33_ASAP7_75t_L g15021 ( 
.A1(n_14900),
.A2(n_2872),
.A3(n_2867),
.B(n_2871),
.Y(n_15021)
);

INVx1_ASAP7_75t_L g15022 ( 
.A(n_14838),
.Y(n_15022)
);

INVx1_ASAP7_75t_L g15023 ( 
.A(n_14828),
.Y(n_15023)
);

INVxp67_ASAP7_75t_L g15024 ( 
.A(n_14845),
.Y(n_15024)
);

NOR3xp33_ASAP7_75t_L g15025 ( 
.A(n_14833),
.B(n_2872),
.C(n_2873),
.Y(n_15025)
);

OAI32xp33_ASAP7_75t_L g15026 ( 
.A1(n_14930),
.A2(n_2876),
.A3(n_2874),
.B1(n_2875),
.B2(n_2877),
.Y(n_15026)
);

OAI21xp33_ASAP7_75t_L g15027 ( 
.A1(n_14910),
.A2(n_2874),
.B(n_2875),
.Y(n_15027)
);

OAI21xp5_ASAP7_75t_L g15028 ( 
.A1(n_14880),
.A2(n_2878),
.B(n_2880),
.Y(n_15028)
);

AOI322xp5_ASAP7_75t_L g15029 ( 
.A1(n_14889),
.A2(n_2885),
.A3(n_2884),
.B1(n_2882),
.B2(n_2878),
.C1(n_2881),
.C2(n_2883),
.Y(n_15029)
);

HB1xp67_ASAP7_75t_L g15030 ( 
.A(n_14843),
.Y(n_15030)
);

OAI221xp5_ASAP7_75t_L g15031 ( 
.A1(n_14855),
.A2(n_2883),
.B1(n_2881),
.B2(n_2882),
.C(n_2884),
.Y(n_15031)
);

INVxp67_ASAP7_75t_L g15032 ( 
.A(n_14926),
.Y(n_15032)
);

XOR2x2_ASAP7_75t_L g15033 ( 
.A(n_14912),
.B(n_2886),
.Y(n_15033)
);

AOI21xp5_ASAP7_75t_L g15034 ( 
.A1(n_14918),
.A2(n_14903),
.B(n_14909),
.Y(n_15034)
);

INVx1_ASAP7_75t_L g15035 ( 
.A(n_14916),
.Y(n_15035)
);

AOI21xp33_ASAP7_75t_L g15036 ( 
.A1(n_14846),
.A2(n_2886),
.B(n_2887),
.Y(n_15036)
);

NAND2xp33_ASAP7_75t_R g15037 ( 
.A(n_14928),
.B(n_2887),
.Y(n_15037)
);

INVx1_ASAP7_75t_L g15038 ( 
.A(n_14933),
.Y(n_15038)
);

AOI21xp5_ASAP7_75t_L g15039 ( 
.A1(n_14920),
.A2(n_2888),
.B(n_2889),
.Y(n_15039)
);

AOI221xp5_ASAP7_75t_L g15040 ( 
.A1(n_14853),
.A2(n_2890),
.B1(n_2888),
.B2(n_2889),
.C(n_2891),
.Y(n_15040)
);

OAI221xp5_ASAP7_75t_L g15041 ( 
.A1(n_14861),
.A2(n_2893),
.B1(n_2891),
.B2(n_2892),
.C(n_2894),
.Y(n_15041)
);

HB1xp67_ASAP7_75t_L g15042 ( 
.A(n_14862),
.Y(n_15042)
);

NOR2x1_ASAP7_75t_L g15043 ( 
.A(n_14854),
.B(n_2892),
.Y(n_15043)
);

AOI22xp5_ASAP7_75t_L g15044 ( 
.A1(n_14878),
.A2(n_2895),
.B1(n_2893),
.B2(n_2894),
.Y(n_15044)
);

OAI21xp33_ASAP7_75t_L g15045 ( 
.A1(n_14859),
.A2(n_2895),
.B(n_2896),
.Y(n_15045)
);

AOI22xp5_ASAP7_75t_L g15046 ( 
.A1(n_14826),
.A2(n_2898),
.B1(n_2896),
.B2(n_2897),
.Y(n_15046)
);

AOI22xp5_ASAP7_75t_L g15047 ( 
.A1(n_14899),
.A2(n_2900),
.B1(n_2897),
.B2(n_2899),
.Y(n_15047)
);

INVx2_ASAP7_75t_L g15048 ( 
.A(n_14824),
.Y(n_15048)
);

INVx1_ASAP7_75t_L g15049 ( 
.A(n_14913),
.Y(n_15049)
);

INVx1_ASAP7_75t_L g15050 ( 
.A(n_14913),
.Y(n_15050)
);

INVx1_ASAP7_75t_L g15051 ( 
.A(n_14913),
.Y(n_15051)
);

INVx2_ASAP7_75t_SL g15052 ( 
.A(n_14824),
.Y(n_15052)
);

OAI21xp33_ASAP7_75t_SL g15053 ( 
.A1(n_14835),
.A2(n_2900),
.B(n_2901),
.Y(n_15053)
);

OAI222xp33_ASAP7_75t_L g15054 ( 
.A1(n_14835),
.A2(n_2903),
.B1(n_2905),
.B2(n_2901),
.C1(n_2902),
.C2(n_2904),
.Y(n_15054)
);

AOI22xp5_ASAP7_75t_L g15055 ( 
.A1(n_14836),
.A2(n_2906),
.B1(n_2902),
.B2(n_2905),
.Y(n_15055)
);

AOI22xp5_ASAP7_75t_L g15056 ( 
.A1(n_14836),
.A2(n_2908),
.B1(n_2906),
.B2(n_2907),
.Y(n_15056)
);

OAI22xp5_ASAP7_75t_L g15057 ( 
.A1(n_14835),
.A2(n_2909),
.B1(n_2907),
.B2(n_2908),
.Y(n_15057)
);

AOI22xp5_ASAP7_75t_L g15058 ( 
.A1(n_14836),
.A2(n_2911),
.B1(n_2909),
.B2(n_2910),
.Y(n_15058)
);

A2O1A1Ixp33_ASAP7_75t_L g15059 ( 
.A1(n_14818),
.A2(n_2912),
.B(n_2910),
.C(n_2911),
.Y(n_15059)
);

NAND2xp5_ASAP7_75t_L g15060 ( 
.A(n_14835),
.B(n_2912),
.Y(n_15060)
);

NOR3xp33_ASAP7_75t_L g15061 ( 
.A(n_14865),
.B(n_2913),
.C(n_2914),
.Y(n_15061)
);

OAI22xp33_ASAP7_75t_SL g15062 ( 
.A1(n_14824),
.A2(n_2915),
.B1(n_2913),
.B2(n_2914),
.Y(n_15062)
);

A2O1A1Ixp33_ASAP7_75t_L g15063 ( 
.A1(n_14818),
.A2(n_2917),
.B(n_2915),
.C(n_2916),
.Y(n_15063)
);

INVx1_ASAP7_75t_L g15064 ( 
.A(n_14913),
.Y(n_15064)
);

NOR3xp33_ASAP7_75t_L g15065 ( 
.A(n_14865),
.B(n_2916),
.C(n_2917),
.Y(n_15065)
);

NAND2xp5_ASAP7_75t_L g15066 ( 
.A(n_15007),
.B(n_2918),
.Y(n_15066)
);

O2A1O1Ixp33_ASAP7_75t_L g15067 ( 
.A1(n_14941),
.A2(n_2921),
.B(n_2919),
.C(n_2920),
.Y(n_15067)
);

OAI22xp5_ASAP7_75t_L g15068 ( 
.A1(n_14938),
.A2(n_2921),
.B1(n_2919),
.B2(n_2920),
.Y(n_15068)
);

OAI21xp33_ASAP7_75t_L g15069 ( 
.A1(n_14972),
.A2(n_2922),
.B(n_2923),
.Y(n_15069)
);

AND2x2_ASAP7_75t_L g15070 ( 
.A(n_15049),
.B(n_2922),
.Y(n_15070)
);

NAND2xp5_ASAP7_75t_L g15071 ( 
.A(n_15052),
.B(n_2924),
.Y(n_15071)
);

INVx1_ASAP7_75t_L g15072 ( 
.A(n_14952),
.Y(n_15072)
);

OAI222xp33_ASAP7_75t_L g15073 ( 
.A1(n_15050),
.A2(n_2926),
.B1(n_2928),
.B2(n_2924),
.C1(n_2925),
.C2(n_2927),
.Y(n_15073)
);

AOI22xp5_ASAP7_75t_L g15074 ( 
.A1(n_15051),
.A2(n_2929),
.B1(n_2926),
.B2(n_2928),
.Y(n_15074)
);

INVx1_ASAP7_75t_L g15075 ( 
.A(n_14952),
.Y(n_15075)
);

INVx1_ASAP7_75t_SL g15076 ( 
.A(n_14979),
.Y(n_15076)
);

INVx2_ASAP7_75t_L g15077 ( 
.A(n_14953),
.Y(n_15077)
);

OAI31xp33_ASAP7_75t_L g15078 ( 
.A1(n_14948),
.A2(n_2931),
.A3(n_2929),
.B(n_2930),
.Y(n_15078)
);

INVx2_ASAP7_75t_L g15079 ( 
.A(n_14970),
.Y(n_15079)
);

AOI21xp33_ASAP7_75t_L g15080 ( 
.A1(n_14954),
.A2(n_2930),
.B(n_2931),
.Y(n_15080)
);

INVx1_ASAP7_75t_L g15081 ( 
.A(n_15030),
.Y(n_15081)
);

NAND2xp5_ASAP7_75t_L g15082 ( 
.A(n_14942),
.B(n_2932),
.Y(n_15082)
);

AOI21xp33_ASAP7_75t_SL g15083 ( 
.A1(n_15064),
.A2(n_2932),
.B(n_2933),
.Y(n_15083)
);

NOR2xp33_ASAP7_75t_L g15084 ( 
.A(n_14955),
.B(n_2934),
.Y(n_15084)
);

AOI221xp5_ASAP7_75t_L g15085 ( 
.A1(n_15024),
.A2(n_14963),
.B1(n_15011),
.B2(n_15009),
.C(n_14959),
.Y(n_15085)
);

OAI21xp5_ASAP7_75t_L g15086 ( 
.A1(n_15053),
.A2(n_2934),
.B(n_2935),
.Y(n_15086)
);

INVx1_ASAP7_75t_L g15087 ( 
.A(n_14993),
.Y(n_15087)
);

INVx2_ASAP7_75t_L g15088 ( 
.A(n_14944),
.Y(n_15088)
);

HB1xp67_ASAP7_75t_L g15089 ( 
.A(n_14946),
.Y(n_15089)
);

NAND2xp5_ASAP7_75t_L g15090 ( 
.A(n_15048),
.B(n_14977),
.Y(n_15090)
);

A2O1A1Ixp33_ASAP7_75t_L g15091 ( 
.A1(n_14939),
.A2(n_2937),
.B(n_2935),
.C(n_2936),
.Y(n_15091)
);

AOI22xp5_ASAP7_75t_L g15092 ( 
.A1(n_14984),
.A2(n_2938),
.B1(n_2936),
.B2(n_2937),
.Y(n_15092)
);

INVx1_ASAP7_75t_L g15093 ( 
.A(n_14983),
.Y(n_15093)
);

OR2x2_ASAP7_75t_L g15094 ( 
.A(n_15002),
.B(n_14991),
.Y(n_15094)
);

AOI211xp5_ASAP7_75t_L g15095 ( 
.A1(n_14937),
.A2(n_2940),
.B(n_2938),
.C(n_2939),
.Y(n_15095)
);

INVx2_ASAP7_75t_L g15096 ( 
.A(n_14964),
.Y(n_15096)
);

INVx2_ASAP7_75t_SL g15097 ( 
.A(n_15003),
.Y(n_15097)
);

NOR2x1p5_ASAP7_75t_L g15098 ( 
.A(n_14973),
.B(n_2939),
.Y(n_15098)
);

AND2x2_ASAP7_75t_L g15099 ( 
.A(n_14988),
.B(n_2940),
.Y(n_15099)
);

NOR2xp67_ASAP7_75t_L g15100 ( 
.A(n_14974),
.B(n_2941),
.Y(n_15100)
);

INVxp67_ASAP7_75t_SL g15101 ( 
.A(n_14961),
.Y(n_15101)
);

INVxp67_ASAP7_75t_L g15102 ( 
.A(n_14947),
.Y(n_15102)
);

INVx1_ASAP7_75t_L g15103 ( 
.A(n_14968),
.Y(n_15103)
);

INVx1_ASAP7_75t_L g15104 ( 
.A(n_14996),
.Y(n_15104)
);

INVx1_ASAP7_75t_L g15105 ( 
.A(n_15060),
.Y(n_15105)
);

AND2x2_ASAP7_75t_L g15106 ( 
.A(n_15043),
.B(n_2941),
.Y(n_15106)
);

NAND2xp5_ASAP7_75t_L g15107 ( 
.A(n_14957),
.B(n_2942),
.Y(n_15107)
);

AOI22xp5_ASAP7_75t_L g15108 ( 
.A1(n_14971),
.A2(n_2944),
.B1(n_2942),
.B2(n_2943),
.Y(n_15108)
);

NOR2xp67_ASAP7_75t_L g15109 ( 
.A(n_14995),
.B(n_2943),
.Y(n_15109)
);

AOI22xp5_ASAP7_75t_L g15110 ( 
.A1(n_15023),
.A2(n_2947),
.B1(n_2945),
.B2(n_2946),
.Y(n_15110)
);

NAND2xp5_ASAP7_75t_L g15111 ( 
.A(n_14986),
.B(n_2945),
.Y(n_15111)
);

INVx1_ASAP7_75t_L g15112 ( 
.A(n_15015),
.Y(n_15112)
);

AOI322xp5_ASAP7_75t_L g15113 ( 
.A1(n_15035),
.A2(n_2951),
.A3(n_2950),
.B1(n_2948),
.B2(n_2946),
.C1(n_2947),
.C2(n_2949),
.Y(n_15113)
);

NAND2xp5_ASAP7_75t_L g15114 ( 
.A(n_14985),
.B(n_2948),
.Y(n_15114)
);

AND2x2_ASAP7_75t_L g15115 ( 
.A(n_15061),
.B(n_2949),
.Y(n_15115)
);

INVxp67_ASAP7_75t_L g15116 ( 
.A(n_15037),
.Y(n_15116)
);

NAND2xp5_ASAP7_75t_L g15117 ( 
.A(n_15012),
.B(n_2950),
.Y(n_15117)
);

OAI21xp5_ASAP7_75t_SL g15118 ( 
.A1(n_14989),
.A2(n_2951),
.B(n_2952),
.Y(n_15118)
);

NAND2xp5_ASAP7_75t_L g15119 ( 
.A(n_14980),
.B(n_2952),
.Y(n_15119)
);

AOI22xp33_ASAP7_75t_L g15120 ( 
.A1(n_15019),
.A2(n_2956),
.B1(n_2954),
.B2(n_2955),
.Y(n_15120)
);

INVx2_ASAP7_75t_L g15121 ( 
.A(n_15033),
.Y(n_15121)
);

AND2x2_ASAP7_75t_L g15122 ( 
.A(n_15065),
.B(n_2954),
.Y(n_15122)
);

OAI21xp5_ASAP7_75t_L g15123 ( 
.A1(n_15034),
.A2(n_14990),
.B(n_15039),
.Y(n_15123)
);

INVx1_ASAP7_75t_L g15124 ( 
.A(n_15062),
.Y(n_15124)
);

OAI32xp33_ASAP7_75t_SL g15125 ( 
.A1(n_15000),
.A2(n_2958),
.A3(n_2956),
.B1(n_2957),
.B2(n_2959),
.Y(n_15125)
);

AND2x2_ASAP7_75t_L g15126 ( 
.A(n_14994),
.B(n_14943),
.Y(n_15126)
);

INVx2_ASAP7_75t_L g15127 ( 
.A(n_15038),
.Y(n_15127)
);

AND2x2_ASAP7_75t_L g15128 ( 
.A(n_14958),
.B(n_2957),
.Y(n_15128)
);

NOR2xp33_ASAP7_75t_L g15129 ( 
.A(n_15032),
.B(n_2958),
.Y(n_15129)
);

NOR2xp33_ASAP7_75t_L g15130 ( 
.A(n_15054),
.B(n_2959),
.Y(n_15130)
);

NOR2xp33_ASAP7_75t_L g15131 ( 
.A(n_14981),
.B(n_2960),
.Y(n_15131)
);

OAI22xp5_ASAP7_75t_SL g15132 ( 
.A1(n_15031),
.A2(n_2962),
.B1(n_2960),
.B2(n_2961),
.Y(n_15132)
);

AOI321xp33_ASAP7_75t_L g15133 ( 
.A1(n_15022),
.A2(n_2963),
.A3(n_2965),
.B1(n_2961),
.B2(n_2962),
.C(n_2964),
.Y(n_15133)
);

NAND3x2_ASAP7_75t_L g15134 ( 
.A(n_14975),
.B(n_2963),
.C(n_2964),
.Y(n_15134)
);

INVx1_ASAP7_75t_L g15135 ( 
.A(n_14982),
.Y(n_15135)
);

OAI21xp5_ASAP7_75t_L g15136 ( 
.A1(n_15005),
.A2(n_2965),
.B(n_2966),
.Y(n_15136)
);

AOI21xp33_ASAP7_75t_SL g15137 ( 
.A1(n_14945),
.A2(n_2966),
.B(n_2967),
.Y(n_15137)
);

INVx1_ASAP7_75t_L g15138 ( 
.A(n_15004),
.Y(n_15138)
);

INVx1_ASAP7_75t_L g15139 ( 
.A(n_14992),
.Y(n_15139)
);

INVx2_ASAP7_75t_L g15140 ( 
.A(n_15008),
.Y(n_15140)
);

INVx1_ASAP7_75t_L g15141 ( 
.A(n_15018),
.Y(n_15141)
);

INVx1_ASAP7_75t_L g15142 ( 
.A(n_15042),
.Y(n_15142)
);

NOR2xp33_ASAP7_75t_SL g15143 ( 
.A(n_15021),
.B(n_2967),
.Y(n_15143)
);

AOI21xp5_ASAP7_75t_L g15144 ( 
.A1(n_15059),
.A2(n_2968),
.B(n_2969),
.Y(n_15144)
);

AOI221xp5_ASAP7_75t_L g15145 ( 
.A1(n_15027),
.A2(n_2970),
.B1(n_2968),
.B2(n_2969),
.C(n_2971),
.Y(n_15145)
);

INVx1_ASAP7_75t_L g15146 ( 
.A(n_15001),
.Y(n_15146)
);

AOI21xp5_ASAP7_75t_L g15147 ( 
.A1(n_15063),
.A2(n_15057),
.B(n_14935),
.Y(n_15147)
);

OAI221xp5_ASAP7_75t_L g15148 ( 
.A1(n_14940),
.A2(n_2973),
.B1(n_2971),
.B2(n_2972),
.C(n_2975),
.Y(n_15148)
);

INVx1_ASAP7_75t_SL g15149 ( 
.A(n_14965),
.Y(n_15149)
);

NAND2xp5_ASAP7_75t_L g15150 ( 
.A(n_15013),
.B(n_2972),
.Y(n_15150)
);

AOI221xp5_ASAP7_75t_L g15151 ( 
.A1(n_15017),
.A2(n_2976),
.B1(n_2973),
.B2(n_2975),
.C(n_2977),
.Y(n_15151)
);

NAND2xp5_ASAP7_75t_L g15152 ( 
.A(n_15020),
.B(n_2976),
.Y(n_15152)
);

INVx2_ASAP7_75t_L g15153 ( 
.A(n_15047),
.Y(n_15153)
);

INVx1_ASAP7_75t_L g15154 ( 
.A(n_14950),
.Y(n_15154)
);

AOI21xp33_ASAP7_75t_SL g15155 ( 
.A1(n_15025),
.A2(n_2977),
.B(n_2978),
.Y(n_15155)
);

INVx2_ASAP7_75t_L g15156 ( 
.A(n_15041),
.Y(n_15156)
);

NAND2xp5_ASAP7_75t_L g15157 ( 
.A(n_14951),
.B(n_2978),
.Y(n_15157)
);

AND2x4_ASAP7_75t_L g15158 ( 
.A(n_15028),
.B(n_2979),
.Y(n_15158)
);

OAI22xp33_ASAP7_75t_L g15159 ( 
.A1(n_15044),
.A2(n_2981),
.B1(n_2979),
.B2(n_2980),
.Y(n_15159)
);

A2O1A1Ixp33_ASAP7_75t_L g15160 ( 
.A1(n_14976),
.A2(n_2982),
.B(n_2980),
.C(n_2981),
.Y(n_15160)
);

NOR2xp67_ASAP7_75t_L g15161 ( 
.A(n_14936),
.B(n_2982),
.Y(n_15161)
);

AND2x4_ASAP7_75t_L g15162 ( 
.A(n_15014),
.B(n_2983),
.Y(n_15162)
);

INVx1_ASAP7_75t_L g15163 ( 
.A(n_14997),
.Y(n_15163)
);

OR2x2_ASAP7_75t_L g15164 ( 
.A(n_15006),
.B(n_2984),
.Y(n_15164)
);

OAI221xp5_ASAP7_75t_L g15165 ( 
.A1(n_15046),
.A2(n_2988),
.B1(n_2985),
.B2(n_2987),
.C(n_2989),
.Y(n_15165)
);

NAND2xp5_ASAP7_75t_L g15166 ( 
.A(n_15045),
.B(n_2987),
.Y(n_15166)
);

XOR2xp5_ASAP7_75t_L g15167 ( 
.A(n_15055),
.B(n_15056),
.Y(n_15167)
);

OR2x2_ASAP7_75t_L g15168 ( 
.A(n_14949),
.B(n_14960),
.Y(n_15168)
);

INVx1_ASAP7_75t_L g15169 ( 
.A(n_14999),
.Y(n_15169)
);

NAND2xp5_ASAP7_75t_L g15170 ( 
.A(n_14998),
.B(n_2988),
.Y(n_15170)
);

INVx2_ASAP7_75t_L g15171 ( 
.A(n_14967),
.Y(n_15171)
);

AOI22xp5_ASAP7_75t_L g15172 ( 
.A1(n_15016),
.A2(n_2991),
.B1(n_2989),
.B2(n_2990),
.Y(n_15172)
);

INVx2_ASAP7_75t_SL g15173 ( 
.A(n_14978),
.Y(n_15173)
);

INVx1_ASAP7_75t_L g15174 ( 
.A(n_14987),
.Y(n_15174)
);

INVx1_ASAP7_75t_L g15175 ( 
.A(n_14962),
.Y(n_15175)
);

OAI222xp33_ASAP7_75t_L g15176 ( 
.A1(n_14966),
.A2(n_2993),
.B1(n_2995),
.B2(n_2991),
.C1(n_2992),
.C2(n_2994),
.Y(n_15176)
);

AND2x2_ASAP7_75t_L g15177 ( 
.A(n_15036),
.B(n_15058),
.Y(n_15177)
);

INVx1_ASAP7_75t_L g15178 ( 
.A(n_14969),
.Y(n_15178)
);

OAI21xp5_ASAP7_75t_L g15179 ( 
.A1(n_15026),
.A2(n_2992),
.B(n_2993),
.Y(n_15179)
);

AOI22xp5_ASAP7_75t_L g15180 ( 
.A1(n_15081),
.A2(n_15010),
.B1(n_15040),
.B2(n_14956),
.Y(n_15180)
);

AOI221xp5_ASAP7_75t_L g15181 ( 
.A1(n_15085),
.A2(n_15029),
.B1(n_2997),
.B2(n_2994),
.C(n_2996),
.Y(n_15181)
);

AOI21xp5_ASAP7_75t_SL g15182 ( 
.A1(n_15067),
.A2(n_2996),
.B(n_2997),
.Y(n_15182)
);

AOI21xp5_ASAP7_75t_SL g15183 ( 
.A1(n_15094),
.A2(n_2998),
.B(n_2999),
.Y(n_15183)
);

INVx1_ASAP7_75t_L g15184 ( 
.A(n_15072),
.Y(n_15184)
);

NAND4xp25_ASAP7_75t_L g15185 ( 
.A(n_15093),
.B(n_15104),
.C(n_15090),
.D(n_15095),
.Y(n_15185)
);

INVx1_ASAP7_75t_L g15186 ( 
.A(n_15075),
.Y(n_15186)
);

OAI22xp5_ASAP7_75t_L g15187 ( 
.A1(n_15108),
.A2(n_3002),
.B1(n_3000),
.B2(n_3001),
.Y(n_15187)
);

NOR4xp25_ASAP7_75t_L g15188 ( 
.A(n_15087),
.B(n_15116),
.C(n_15097),
.D(n_15123),
.Y(n_15188)
);

INVx1_ASAP7_75t_L g15189 ( 
.A(n_15089),
.Y(n_15189)
);

AOI221xp5_ASAP7_75t_L g15190 ( 
.A1(n_15125),
.A2(n_3002),
.B1(n_3000),
.B2(n_3001),
.C(n_3003),
.Y(n_15190)
);

AND2x2_ASAP7_75t_L g15191 ( 
.A(n_15102),
.B(n_3003),
.Y(n_15191)
);

OAI211xp5_ASAP7_75t_L g15192 ( 
.A1(n_15078),
.A2(n_3006),
.B(n_3004),
.C(n_3005),
.Y(n_15192)
);

AOI211xp5_ASAP7_75t_L g15193 ( 
.A1(n_15118),
.A2(n_3008),
.B(n_3006),
.C(n_3007),
.Y(n_15193)
);

OAI221xp5_ASAP7_75t_L g15194 ( 
.A1(n_15091),
.A2(n_3009),
.B1(n_3007),
.B2(n_3008),
.C(n_3010),
.Y(n_15194)
);

OA21x2_ASAP7_75t_L g15195 ( 
.A1(n_15071),
.A2(n_15114),
.B(n_15119),
.Y(n_15195)
);

NAND3xp33_ASAP7_75t_SL g15196 ( 
.A(n_15076),
.B(n_3009),
.C(n_3010),
.Y(n_15196)
);

OA22x2_ASAP7_75t_L g15197 ( 
.A1(n_15172),
.A2(n_3013),
.B1(n_3011),
.B2(n_3012),
.Y(n_15197)
);

O2A1O1Ixp33_ASAP7_75t_L g15198 ( 
.A1(n_15117),
.A2(n_3014),
.B(n_3012),
.C(n_3013),
.Y(n_15198)
);

AOI211xp5_ASAP7_75t_SL g15199 ( 
.A1(n_15101),
.A2(n_3017),
.B(n_3015),
.C(n_3016),
.Y(n_15199)
);

AOI322xp5_ASAP7_75t_L g15200 ( 
.A1(n_15106),
.A2(n_3020),
.A3(n_3019),
.B1(n_3017),
.B2(n_3015),
.C1(n_3016),
.C2(n_3018),
.Y(n_15200)
);

XOR2x2_ASAP7_75t_L g15201 ( 
.A(n_15134),
.B(n_3018),
.Y(n_15201)
);

OAI22xp5_ASAP7_75t_L g15202 ( 
.A1(n_15148),
.A2(n_3021),
.B1(n_3019),
.B2(n_3020),
.Y(n_15202)
);

NOR2x1_ASAP7_75t_L g15203 ( 
.A(n_15082),
.B(n_3021),
.Y(n_15203)
);

INVx1_ASAP7_75t_L g15204 ( 
.A(n_15142),
.Y(n_15204)
);

AOI22xp5_ASAP7_75t_L g15205 ( 
.A1(n_15130),
.A2(n_3024),
.B1(n_3022),
.B2(n_3023),
.Y(n_15205)
);

INVx1_ASAP7_75t_L g15206 ( 
.A(n_15099),
.Y(n_15206)
);

OAI21xp33_ASAP7_75t_L g15207 ( 
.A1(n_15126),
.A2(n_15143),
.B(n_15088),
.Y(n_15207)
);

AOI221xp5_ASAP7_75t_L g15208 ( 
.A1(n_15155),
.A2(n_3025),
.B1(n_3023),
.B2(n_3024),
.C(n_3026),
.Y(n_15208)
);

AOI21xp5_ASAP7_75t_L g15209 ( 
.A1(n_15150),
.A2(n_3025),
.B(n_3026),
.Y(n_15209)
);

OAI221xp5_ASAP7_75t_L g15210 ( 
.A1(n_15069),
.A2(n_3029),
.B1(n_3027),
.B2(n_3028),
.C(n_3030),
.Y(n_15210)
);

OAI211xp5_ASAP7_75t_L g15211 ( 
.A1(n_15080),
.A2(n_3032),
.B(n_3027),
.C(n_3029),
.Y(n_15211)
);

AOI322xp5_ASAP7_75t_L g15212 ( 
.A1(n_15124),
.A2(n_3038),
.A3(n_3037),
.B1(n_3035),
.B2(n_3033),
.C1(n_3034),
.C2(n_3036),
.Y(n_15212)
);

OAI21xp5_ASAP7_75t_L g15213 ( 
.A1(n_15100),
.A2(n_3033),
.B(n_3034),
.Y(n_15213)
);

OAI31xp33_ASAP7_75t_L g15214 ( 
.A1(n_15098),
.A2(n_3037),
.A3(n_3035),
.B(n_3036),
.Y(n_15214)
);

AO22x1_ASAP7_75t_L g15215 ( 
.A1(n_15136),
.A2(n_3040),
.B1(n_3038),
.B2(n_3039),
.Y(n_15215)
);

AOI22xp5_ASAP7_75t_L g15216 ( 
.A1(n_15079),
.A2(n_3041),
.B1(n_3039),
.B2(n_3040),
.Y(n_15216)
);

NAND2xp5_ASAP7_75t_SL g15217 ( 
.A(n_15133),
.B(n_3041),
.Y(n_15217)
);

OAI21xp5_ASAP7_75t_L g15218 ( 
.A1(n_15086),
.A2(n_3042),
.B(n_3043),
.Y(n_15218)
);

NAND4xp25_ASAP7_75t_SL g15219 ( 
.A(n_15145),
.B(n_15151),
.C(n_15147),
.D(n_15157),
.Y(n_15219)
);

AOI21xp33_ASAP7_75t_L g15220 ( 
.A1(n_15096),
.A2(n_3043),
.B(n_3044),
.Y(n_15220)
);

AOI21xp5_ASAP7_75t_L g15221 ( 
.A1(n_15066),
.A2(n_3044),
.B(n_3045),
.Y(n_15221)
);

AOI221xp5_ASAP7_75t_L g15222 ( 
.A1(n_15137),
.A2(n_3047),
.B1(n_3045),
.B2(n_3046),
.C(n_3048),
.Y(n_15222)
);

AOI211xp5_ASAP7_75t_SL g15223 ( 
.A1(n_15084),
.A2(n_3048),
.B(n_3046),
.C(n_3047),
.Y(n_15223)
);

NAND4xp25_ASAP7_75t_SL g15224 ( 
.A(n_15144),
.B(n_3051),
.C(n_3049),
.D(n_3050),
.Y(n_15224)
);

NOR2xp33_ASAP7_75t_SL g15225 ( 
.A(n_15073),
.B(n_15127),
.Y(n_15225)
);

AOI22xp5_ASAP7_75t_L g15226 ( 
.A1(n_15109),
.A2(n_3052),
.B1(n_3049),
.B2(n_3050),
.Y(n_15226)
);

AOI22xp5_ASAP7_75t_L g15227 ( 
.A1(n_15077),
.A2(n_3055),
.B1(n_3052),
.B2(n_3053),
.Y(n_15227)
);

AOI31xp33_ASAP7_75t_L g15228 ( 
.A1(n_15112),
.A2(n_3058),
.A3(n_3053),
.B(n_3056),
.Y(n_15228)
);

OAI221xp5_ASAP7_75t_L g15229 ( 
.A1(n_15179),
.A2(n_3059),
.B1(n_3056),
.B2(n_3058),
.C(n_3060),
.Y(n_15229)
);

INVx1_ASAP7_75t_L g15230 ( 
.A(n_15070),
.Y(n_15230)
);

INVx2_ASAP7_75t_L g15231 ( 
.A(n_15164),
.Y(n_15231)
);

NOR2xp33_ASAP7_75t_L g15232 ( 
.A(n_15083),
.B(n_3060),
.Y(n_15232)
);

AOI22xp5_ASAP7_75t_L g15233 ( 
.A1(n_15177),
.A2(n_3063),
.B1(n_3061),
.B2(n_3062),
.Y(n_15233)
);

OAI21xp33_ASAP7_75t_SL g15234 ( 
.A1(n_15152),
.A2(n_3061),
.B(n_3062),
.Y(n_15234)
);

AOI211xp5_ASAP7_75t_L g15235 ( 
.A1(n_15132),
.A2(n_3065),
.B(n_3063),
.C(n_3064),
.Y(n_15235)
);

XNOR2xp5_ASAP7_75t_L g15236 ( 
.A(n_15167),
.B(n_3065),
.Y(n_15236)
);

AOI211xp5_ASAP7_75t_L g15237 ( 
.A1(n_15159),
.A2(n_15165),
.B(n_15176),
.C(n_15131),
.Y(n_15237)
);

AOI221xp5_ASAP7_75t_L g15238 ( 
.A1(n_15103),
.A2(n_3068),
.B1(n_3066),
.B2(n_3067),
.C(n_3069),
.Y(n_15238)
);

NAND2x1_ASAP7_75t_L g15239 ( 
.A(n_15162),
.B(n_3066),
.Y(n_15239)
);

AOI221xp5_ASAP7_75t_L g15240 ( 
.A1(n_15154),
.A2(n_3069),
.B1(n_3067),
.B2(n_3068),
.C(n_3071),
.Y(n_15240)
);

AOI22xp5_ASAP7_75t_L g15241 ( 
.A1(n_15146),
.A2(n_3073),
.B1(n_3071),
.B2(n_3072),
.Y(n_15241)
);

NAND3xp33_ASAP7_75t_SL g15242 ( 
.A(n_15149),
.B(n_15107),
.C(n_15121),
.Y(n_15242)
);

AOI211xp5_ASAP7_75t_L g15243 ( 
.A1(n_15161),
.A2(n_3075),
.B(n_3072),
.C(n_3074),
.Y(n_15243)
);

O2A1O1Ixp33_ASAP7_75t_L g15244 ( 
.A1(n_15171),
.A2(n_3076),
.B(n_3074),
.C(n_3075),
.Y(n_15244)
);

AOI22xp33_ASAP7_75t_L g15245 ( 
.A1(n_15140),
.A2(n_3078),
.B1(n_3076),
.B2(n_3077),
.Y(n_15245)
);

OR2x2_ASAP7_75t_L g15246 ( 
.A(n_15111),
.B(n_3077),
.Y(n_15246)
);

AOI22xp5_ASAP7_75t_L g15247 ( 
.A1(n_15128),
.A2(n_3081),
.B1(n_3079),
.B2(n_3080),
.Y(n_15247)
);

AOI221x1_ASAP7_75t_L g15248 ( 
.A1(n_15163),
.A2(n_3082),
.B1(n_3079),
.B2(n_3081),
.C(n_3083),
.Y(n_15248)
);

OAI22xp5_ASAP7_75t_L g15249 ( 
.A1(n_15092),
.A2(n_3085),
.B1(n_3083),
.B2(n_3084),
.Y(n_15249)
);

AOI211xp5_ASAP7_75t_L g15250 ( 
.A1(n_15115),
.A2(n_3086),
.B(n_3084),
.C(n_3085),
.Y(n_15250)
);

XNOR2xp5_ASAP7_75t_L g15251 ( 
.A(n_15162),
.B(n_3086),
.Y(n_15251)
);

INVx1_ASAP7_75t_L g15252 ( 
.A(n_15122),
.Y(n_15252)
);

INVx1_ASAP7_75t_L g15253 ( 
.A(n_15158),
.Y(n_15253)
);

AND4x1_ASAP7_75t_L g15254 ( 
.A(n_15129),
.B(n_3089),
.C(n_3087),
.D(n_3088),
.Y(n_15254)
);

AOI322xp5_ASAP7_75t_L g15255 ( 
.A1(n_15173),
.A2(n_15105),
.A3(n_15141),
.B1(n_15139),
.B2(n_15135),
.C1(n_15158),
.C2(n_15138),
.Y(n_15255)
);

AOI21xp5_ASAP7_75t_L g15256 ( 
.A1(n_15068),
.A2(n_3087),
.B(n_3089),
.Y(n_15256)
);

INVx1_ASAP7_75t_L g15257 ( 
.A(n_15166),
.Y(n_15257)
);

AOI322xp5_ASAP7_75t_L g15258 ( 
.A1(n_15174),
.A2(n_3095),
.A3(n_3094),
.B1(n_3092),
.B2(n_3090),
.C1(n_3091),
.C2(n_3093),
.Y(n_15258)
);

INVx1_ASAP7_75t_L g15259 ( 
.A(n_15170),
.Y(n_15259)
);

OAI211xp5_ASAP7_75t_SL g15260 ( 
.A1(n_15169),
.A2(n_3094),
.B(n_3090),
.C(n_3093),
.Y(n_15260)
);

OAI211xp5_ASAP7_75t_SL g15261 ( 
.A1(n_15175),
.A2(n_3097),
.B(n_3095),
.C(n_3096),
.Y(n_15261)
);

NOR2xp33_ASAP7_75t_SL g15262 ( 
.A(n_15153),
.B(n_3096),
.Y(n_15262)
);

O2A1O1Ixp33_ASAP7_75t_L g15263 ( 
.A1(n_15160),
.A2(n_3100),
.B(n_3098),
.C(n_3099),
.Y(n_15263)
);

INVx1_ASAP7_75t_L g15264 ( 
.A(n_15168),
.Y(n_15264)
);

OAI221xp5_ASAP7_75t_L g15265 ( 
.A1(n_15120),
.A2(n_3102),
.B1(n_3098),
.B2(n_3101),
.C(n_3103),
.Y(n_15265)
);

AOI22xp5_ASAP7_75t_L g15266 ( 
.A1(n_15178),
.A2(n_3104),
.B1(n_3101),
.B2(n_3102),
.Y(n_15266)
);

AOI221xp5_ASAP7_75t_L g15267 ( 
.A1(n_15156),
.A2(n_3106),
.B1(n_3104),
.B2(n_3105),
.C(n_3107),
.Y(n_15267)
);

NAND2xp5_ASAP7_75t_SL g15268 ( 
.A(n_15074),
.B(n_3105),
.Y(n_15268)
);

OAI22xp5_ASAP7_75t_L g15269 ( 
.A1(n_15110),
.A2(n_3110),
.B1(n_3107),
.B2(n_3109),
.Y(n_15269)
);

AOI22xp5_ASAP7_75t_L g15270 ( 
.A1(n_15113),
.A2(n_3111),
.B1(n_3109),
.B2(n_3110),
.Y(n_15270)
);

OAI321xp33_ASAP7_75t_L g15271 ( 
.A1(n_15116),
.A2(n_3113),
.A3(n_3115),
.B1(n_3111),
.B2(n_3112),
.C(n_3114),
.Y(n_15271)
);

NOR3xp33_ASAP7_75t_L g15272 ( 
.A(n_15081),
.B(n_3112),
.C(n_3113),
.Y(n_15272)
);

NAND3xp33_ASAP7_75t_L g15273 ( 
.A(n_15085),
.B(n_3115),
.C(n_3116),
.Y(n_15273)
);

AOI211xp5_ASAP7_75t_L g15274 ( 
.A1(n_15081),
.A2(n_3119),
.B(n_3120),
.C(n_3118),
.Y(n_15274)
);

INVx1_ASAP7_75t_L g15275 ( 
.A(n_15072),
.Y(n_15275)
);

OAI21xp33_ASAP7_75t_L g15276 ( 
.A1(n_15087),
.A2(n_3117),
.B(n_3118),
.Y(n_15276)
);

AOI21xp5_ASAP7_75t_L g15277 ( 
.A1(n_15081),
.A2(n_3117),
.B(n_3120),
.Y(n_15277)
);

AOI21xp5_ASAP7_75t_L g15278 ( 
.A1(n_15081),
.A2(n_3121),
.B(n_3122),
.Y(n_15278)
);

NOR2x1_ASAP7_75t_L g15279 ( 
.A(n_15081),
.B(n_3121),
.Y(n_15279)
);

NOR4xp25_ASAP7_75t_L g15280 ( 
.A(n_15081),
.B(n_3124),
.C(n_3122),
.D(n_3123),
.Y(n_15280)
);

OAI211xp5_ASAP7_75t_L g15281 ( 
.A1(n_15081),
.A2(n_3125),
.B(n_3123),
.C(n_3124),
.Y(n_15281)
);

AOI211xp5_ASAP7_75t_SL g15282 ( 
.A1(n_15264),
.A2(n_3128),
.B(n_3126),
.C(n_3127),
.Y(n_15282)
);

NAND4xp75_ASAP7_75t_L g15283 ( 
.A(n_15189),
.B(n_3129),
.C(n_3126),
.D(n_3127),
.Y(n_15283)
);

NAND3xp33_ASAP7_75t_L g15284 ( 
.A(n_15184),
.B(n_4119),
.C(n_4118),
.Y(n_15284)
);

AOI222xp33_ASAP7_75t_L g15285 ( 
.A1(n_15186),
.A2(n_3132),
.B1(n_3134),
.B2(n_3130),
.C1(n_3131),
.C2(n_3133),
.Y(n_15285)
);

OAI221xp5_ASAP7_75t_L g15286 ( 
.A1(n_15188),
.A2(n_3134),
.B1(n_3130),
.B2(n_3132),
.C(n_3135),
.Y(n_15286)
);

NOR2xp67_ASAP7_75t_L g15287 ( 
.A(n_15271),
.B(n_3135),
.Y(n_15287)
);

OAI211xp5_ASAP7_75t_L g15288 ( 
.A1(n_15185),
.A2(n_3138),
.B(n_3136),
.C(n_3137),
.Y(n_15288)
);

AOI221xp5_ASAP7_75t_L g15289 ( 
.A1(n_15275),
.A2(n_3141),
.B1(n_3137),
.B2(n_3140),
.C(n_3142),
.Y(n_15289)
);

NAND3xp33_ASAP7_75t_SL g15290 ( 
.A(n_15204),
.B(n_3142),
.C(n_3141),
.Y(n_15290)
);

AOI21xp5_ASAP7_75t_L g15291 ( 
.A1(n_15183),
.A2(n_3140),
.B(n_3143),
.Y(n_15291)
);

OAI21xp33_ASAP7_75t_L g15292 ( 
.A1(n_15225),
.A2(n_3144),
.B(n_3145),
.Y(n_15292)
);

NAND2xp5_ASAP7_75t_L g15293 ( 
.A(n_15279),
.B(n_3145),
.Y(n_15293)
);

AOI211xp5_ASAP7_75t_L g15294 ( 
.A1(n_15229),
.A2(n_3148),
.B(n_3146),
.C(n_3147),
.Y(n_15294)
);

OR2x2_ASAP7_75t_L g15295 ( 
.A(n_15239),
.B(n_3148),
.Y(n_15295)
);

OAI21xp33_ASAP7_75t_L g15296 ( 
.A1(n_15207),
.A2(n_3147),
.B(n_3149),
.Y(n_15296)
);

NAND2xp5_ASAP7_75t_L g15297 ( 
.A(n_15203),
.B(n_3149),
.Y(n_15297)
);

AOI22x1_ASAP7_75t_L g15298 ( 
.A1(n_15251),
.A2(n_3153),
.B1(n_3151),
.B2(n_3152),
.Y(n_15298)
);

AOI211xp5_ASAP7_75t_L g15299 ( 
.A1(n_15280),
.A2(n_15219),
.B(n_15249),
.C(n_15187),
.Y(n_15299)
);

NAND2xp5_ASAP7_75t_L g15300 ( 
.A(n_15206),
.B(n_3152),
.Y(n_15300)
);

AOI21xp33_ASAP7_75t_L g15301 ( 
.A1(n_15230),
.A2(n_3155),
.B(n_3154),
.Y(n_15301)
);

AOI22xp33_ASAP7_75t_L g15302 ( 
.A1(n_15242),
.A2(n_3155),
.B1(n_3153),
.B2(n_3154),
.Y(n_15302)
);

OAI21xp5_ASAP7_75t_SL g15303 ( 
.A1(n_15199),
.A2(n_15223),
.B(n_15205),
.Y(n_15303)
);

NOR2xp33_ASAP7_75t_L g15304 ( 
.A(n_15234),
.B(n_3156),
.Y(n_15304)
);

NOR2xp67_ASAP7_75t_L g15305 ( 
.A(n_15281),
.B(n_3156),
.Y(n_15305)
);

NAND3xp33_ASAP7_75t_L g15306 ( 
.A(n_15255),
.B(n_4112),
.C(n_4111),
.Y(n_15306)
);

INVx1_ASAP7_75t_L g15307 ( 
.A(n_15236),
.Y(n_15307)
);

NAND2xp5_ASAP7_75t_L g15308 ( 
.A(n_15253),
.B(n_3157),
.Y(n_15308)
);

OAI32xp33_ASAP7_75t_L g15309 ( 
.A1(n_15232),
.A2(n_4113),
.A3(n_4114),
.B1(n_4112),
.B2(n_4111),
.Y(n_15309)
);

NAND2xp5_ASAP7_75t_L g15310 ( 
.A(n_15215),
.B(n_3157),
.Y(n_15310)
);

AOI221xp5_ASAP7_75t_L g15311 ( 
.A1(n_15182),
.A2(n_3160),
.B1(n_3158),
.B2(n_3159),
.C(n_3161),
.Y(n_15311)
);

NAND4xp25_ASAP7_75t_L g15312 ( 
.A(n_15243),
.B(n_15235),
.C(n_15193),
.D(n_15181),
.Y(n_15312)
);

INVx1_ASAP7_75t_L g15313 ( 
.A(n_15228),
.Y(n_15313)
);

AOI22xp5_ASAP7_75t_L g15314 ( 
.A1(n_15191),
.A2(n_3160),
.B1(n_3158),
.B2(n_3159),
.Y(n_15314)
);

AOI21xp5_ASAP7_75t_L g15315 ( 
.A1(n_15217),
.A2(n_3163),
.B(n_3164),
.Y(n_15315)
);

NOR3xp33_ASAP7_75t_L g15316 ( 
.A(n_15252),
.B(n_3163),
.C(n_3164),
.Y(n_15316)
);

AOI22x1_ASAP7_75t_L g15317 ( 
.A1(n_15277),
.A2(n_3167),
.B1(n_3165),
.B2(n_3166),
.Y(n_15317)
);

NAND2xp5_ASAP7_75t_L g15318 ( 
.A(n_15254),
.B(n_3165),
.Y(n_15318)
);

AOI22xp5_ASAP7_75t_L g15319 ( 
.A1(n_15180),
.A2(n_3168),
.B1(n_3166),
.B2(n_3167),
.Y(n_15319)
);

AND2x2_ASAP7_75t_L g15320 ( 
.A(n_15195),
.B(n_3168),
.Y(n_15320)
);

NOR2x1_ASAP7_75t_L g15321 ( 
.A(n_15273),
.B(n_15196),
.Y(n_15321)
);

AOI22xp5_ASAP7_75t_L g15322 ( 
.A1(n_15190),
.A2(n_15268),
.B1(n_15270),
.B2(n_15202),
.Y(n_15322)
);

OAI211xp5_ASAP7_75t_L g15323 ( 
.A1(n_15241),
.A2(n_3171),
.B(n_3169),
.C(n_3170),
.Y(n_15323)
);

OAI221xp5_ASAP7_75t_L g15324 ( 
.A1(n_15276),
.A2(n_3172),
.B1(n_3169),
.B2(n_3171),
.C(n_3173),
.Y(n_15324)
);

OAI22xp5_ASAP7_75t_L g15325 ( 
.A1(n_15227),
.A2(n_3175),
.B1(n_3173),
.B2(n_3174),
.Y(n_15325)
);

INVx1_ASAP7_75t_L g15326 ( 
.A(n_15201),
.Y(n_15326)
);

NAND3xp33_ASAP7_75t_SL g15327 ( 
.A(n_15213),
.B(n_3177),
.C(n_3176),
.Y(n_15327)
);

AOI222xp33_ASAP7_75t_L g15328 ( 
.A1(n_15259),
.A2(n_3178),
.B1(n_3180),
.B2(n_3175),
.C1(n_3177),
.C2(n_3179),
.Y(n_15328)
);

NOR3xp33_ASAP7_75t_L g15329 ( 
.A(n_15231),
.B(n_3179),
.C(n_3180),
.Y(n_15329)
);

NOR2xp33_ASAP7_75t_SL g15330 ( 
.A(n_15214),
.B(n_3181),
.Y(n_15330)
);

OAI211xp5_ASAP7_75t_SL g15331 ( 
.A1(n_15209),
.A2(n_3183),
.B(n_3181),
.C(n_3182),
.Y(n_15331)
);

OAI21xp5_ASAP7_75t_SL g15332 ( 
.A1(n_15192),
.A2(n_3184),
.B(n_3183),
.Y(n_15332)
);

AOI311xp33_ASAP7_75t_L g15333 ( 
.A1(n_15237),
.A2(n_3186),
.A3(n_3182),
.B(n_3185),
.C(n_3187),
.Y(n_15333)
);

NAND4xp25_ASAP7_75t_L g15334 ( 
.A(n_15262),
.B(n_3187),
.C(n_3185),
.D(n_3186),
.Y(n_15334)
);

AOI22xp5_ASAP7_75t_L g15335 ( 
.A1(n_15269),
.A2(n_3190),
.B1(n_3188),
.B2(n_3189),
.Y(n_15335)
);

NOR4xp25_ASAP7_75t_L g15336 ( 
.A(n_15257),
.B(n_3193),
.C(n_3191),
.D(n_3192),
.Y(n_15336)
);

OAI221xp5_ASAP7_75t_L g15337 ( 
.A1(n_15210),
.A2(n_3193),
.B1(n_3191),
.B2(n_3192),
.C(n_3194),
.Y(n_15337)
);

NAND2xp5_ASAP7_75t_L g15338 ( 
.A(n_15195),
.B(n_3194),
.Y(n_15338)
);

NAND2xp5_ASAP7_75t_L g15339 ( 
.A(n_15200),
.B(n_3195),
.Y(n_15339)
);

NAND2xp5_ASAP7_75t_SL g15340 ( 
.A(n_15208),
.B(n_3195),
.Y(n_15340)
);

AOI211x1_ASAP7_75t_L g15341 ( 
.A1(n_15218),
.A2(n_3198),
.B(n_3196),
.C(n_3197),
.Y(n_15341)
);

OAI21xp5_ASAP7_75t_L g15342 ( 
.A1(n_15221),
.A2(n_3196),
.B(n_3197),
.Y(n_15342)
);

AOI221xp5_ASAP7_75t_L g15343 ( 
.A1(n_15244),
.A2(n_3200),
.B1(n_3198),
.B2(n_3199),
.C(n_3201),
.Y(n_15343)
);

AOI21xp5_ASAP7_75t_L g15344 ( 
.A1(n_15278),
.A2(n_3199),
.B(n_3200),
.Y(n_15344)
);

AOI211xp5_ASAP7_75t_L g15345 ( 
.A1(n_15194),
.A2(n_3203),
.B(n_3201),
.C(n_3202),
.Y(n_15345)
);

NAND3xp33_ASAP7_75t_L g15346 ( 
.A(n_15272),
.B(n_4108),
.C(n_4107),
.Y(n_15346)
);

AND2x2_ASAP7_75t_L g15347 ( 
.A(n_15197),
.B(n_3202),
.Y(n_15347)
);

NAND2xp5_ASAP7_75t_L g15348 ( 
.A(n_15226),
.B(n_3203),
.Y(n_15348)
);

NAND3xp33_ASAP7_75t_L g15349 ( 
.A(n_15248),
.B(n_4110),
.C(n_4109),
.Y(n_15349)
);

NOR4xp25_ASAP7_75t_L g15350 ( 
.A(n_15198),
.B(n_3206),
.C(n_3204),
.D(n_3205),
.Y(n_15350)
);

AOI21xp5_ASAP7_75t_L g15351 ( 
.A1(n_15220),
.A2(n_3206),
.B(n_3207),
.Y(n_15351)
);

OAI21xp5_ASAP7_75t_SL g15352 ( 
.A1(n_15260),
.A2(n_3209),
.B(n_3208),
.Y(n_15352)
);

A2O1A1Ixp33_ASAP7_75t_L g15353 ( 
.A1(n_15263),
.A2(n_15256),
.B(n_15247),
.C(n_15222),
.Y(n_15353)
);

AOI221xp5_ASAP7_75t_L g15354 ( 
.A1(n_15224),
.A2(n_3210),
.B1(n_3207),
.B2(n_3208),
.C(n_3211),
.Y(n_15354)
);

OAI21xp33_ASAP7_75t_SL g15355 ( 
.A1(n_15246),
.A2(n_3211),
.B(n_3213),
.Y(n_15355)
);

AOI221xp5_ASAP7_75t_L g15356 ( 
.A1(n_15265),
.A2(n_3215),
.B1(n_3213),
.B2(n_3214),
.C(n_3216),
.Y(n_15356)
);

OAI21xp5_ASAP7_75t_L g15357 ( 
.A1(n_15211),
.A2(n_3216),
.B(n_3217),
.Y(n_15357)
);

NAND2xp5_ASAP7_75t_L g15358 ( 
.A(n_15250),
.B(n_15274),
.Y(n_15358)
);

AOI211xp5_ASAP7_75t_L g15359 ( 
.A1(n_15261),
.A2(n_3219),
.B(n_3217),
.C(n_3218),
.Y(n_15359)
);

NOR4xp25_ASAP7_75t_L g15360 ( 
.A(n_15267),
.B(n_15240),
.C(n_15245),
.D(n_15238),
.Y(n_15360)
);

OAI211xp5_ASAP7_75t_L g15361 ( 
.A1(n_15266),
.A2(n_3220),
.B(n_3218),
.C(n_3219),
.Y(n_15361)
);

AOI222xp33_ASAP7_75t_L g15362 ( 
.A1(n_15212),
.A2(n_3222),
.B1(n_3224),
.B2(n_3220),
.C1(n_3221),
.C2(n_3223),
.Y(n_15362)
);

A2O1A1Ixp33_ASAP7_75t_SL g15363 ( 
.A1(n_15216),
.A2(n_3225),
.B(n_3221),
.C(n_3224),
.Y(n_15363)
);

AOI21xp33_ASAP7_75t_SL g15364 ( 
.A1(n_15233),
.A2(n_3234),
.B(n_3225),
.Y(n_15364)
);

NAND2xp5_ASAP7_75t_SL g15365 ( 
.A(n_15258),
.B(n_3226),
.Y(n_15365)
);

XNOR2x2_ASAP7_75t_L g15366 ( 
.A(n_15185),
.B(n_4118),
.Y(n_15366)
);

NAND2xp5_ASAP7_75t_L g15367 ( 
.A(n_15189),
.B(n_3226),
.Y(n_15367)
);

AOI21xp5_ASAP7_75t_L g15368 ( 
.A1(n_15188),
.A2(n_3227),
.B(n_3228),
.Y(n_15368)
);

O2A1O1Ixp33_ASAP7_75t_L g15369 ( 
.A1(n_15189),
.A2(n_3230),
.B(n_3227),
.C(n_3229),
.Y(n_15369)
);

AOI211xp5_ASAP7_75t_L g15370 ( 
.A1(n_15188),
.A2(n_3233),
.B(n_3229),
.C(n_3232),
.Y(n_15370)
);

AOI211xp5_ASAP7_75t_SL g15371 ( 
.A1(n_15264),
.A2(n_3234),
.B(n_3232),
.C(n_3233),
.Y(n_15371)
);

AOI322xp5_ASAP7_75t_L g15372 ( 
.A1(n_15189),
.A2(n_3259),
.A3(n_3243),
.B1(n_3267),
.B2(n_3275),
.C1(n_3251),
.C2(n_3235),
.Y(n_15372)
);

OAI21xp5_ASAP7_75t_L g15373 ( 
.A1(n_15189),
.A2(n_3235),
.B(n_3236),
.Y(n_15373)
);

AOI221xp5_ASAP7_75t_L g15374 ( 
.A1(n_15188),
.A2(n_3238),
.B1(n_3236),
.B2(n_3237),
.C(n_3239),
.Y(n_15374)
);

AOI221xp5_ASAP7_75t_SL g15375 ( 
.A1(n_15264),
.A2(n_3239),
.B1(n_3237),
.B2(n_3238),
.C(n_3240),
.Y(n_15375)
);

OAI21xp5_ASAP7_75t_SL g15376 ( 
.A1(n_15189),
.A2(n_3243),
.B(n_3242),
.Y(n_15376)
);

NAND2xp5_ASAP7_75t_SL g15377 ( 
.A(n_15189),
.B(n_3241),
.Y(n_15377)
);

AOI22xp5_ASAP7_75t_L g15378 ( 
.A1(n_15189),
.A2(n_3244),
.B1(n_3241),
.B2(n_3242),
.Y(n_15378)
);

INVx1_ASAP7_75t_L g15379 ( 
.A(n_15320),
.Y(n_15379)
);

INVx1_ASAP7_75t_L g15380 ( 
.A(n_15295),
.Y(n_15380)
);

INVx1_ASAP7_75t_L g15381 ( 
.A(n_15338),
.Y(n_15381)
);

NAND3xp33_ASAP7_75t_L g15382 ( 
.A(n_15370),
.B(n_15368),
.C(n_15306),
.Y(n_15382)
);

NAND2xp5_ASAP7_75t_L g15383 ( 
.A(n_15304),
.B(n_3245),
.Y(n_15383)
);

AO21x1_ASAP7_75t_L g15384 ( 
.A1(n_15377),
.A2(n_3246),
.B(n_3247),
.Y(n_15384)
);

NAND4xp25_ASAP7_75t_SL g15385 ( 
.A(n_15374),
.B(n_3249),
.C(n_3246),
.D(n_3248),
.Y(n_15385)
);

NAND2xp5_ASAP7_75t_L g15386 ( 
.A(n_15313),
.B(n_3248),
.Y(n_15386)
);

NAND4xp25_ASAP7_75t_SL g15387 ( 
.A(n_15375),
.B(n_3253),
.C(n_3250),
.D(n_3252),
.Y(n_15387)
);

INVx1_ASAP7_75t_L g15388 ( 
.A(n_15366),
.Y(n_15388)
);

XNOR2xp5_ASAP7_75t_L g15389 ( 
.A(n_15307),
.B(n_4108),
.Y(n_15389)
);

AND2x2_ASAP7_75t_L g15390 ( 
.A(n_15347),
.B(n_3250),
.Y(n_15390)
);

INVx1_ASAP7_75t_L g15391 ( 
.A(n_15293),
.Y(n_15391)
);

OAI211xp5_ASAP7_75t_L g15392 ( 
.A1(n_15292),
.A2(n_3255),
.B(n_3253),
.C(n_3254),
.Y(n_15392)
);

OAI22xp33_ASAP7_75t_SL g15393 ( 
.A1(n_15297),
.A2(n_3256),
.B1(n_3254),
.B2(n_3255),
.Y(n_15393)
);

NOR2xp33_ASAP7_75t_L g15394 ( 
.A(n_15355),
.B(n_3257),
.Y(n_15394)
);

INVx1_ASAP7_75t_L g15395 ( 
.A(n_15318),
.Y(n_15395)
);

AOI322xp5_ASAP7_75t_L g15396 ( 
.A1(n_15327),
.A2(n_3263),
.A3(n_3262),
.B1(n_3260),
.B2(n_3258),
.C1(n_3259),
.C2(n_3261),
.Y(n_15396)
);

NOR3xp33_ASAP7_75t_L g15397 ( 
.A(n_15326),
.B(n_3258),
.C(n_3260),
.Y(n_15397)
);

NAND4xp25_ASAP7_75t_L g15398 ( 
.A(n_15333),
.B(n_3265),
.C(n_3263),
.D(n_3264),
.Y(n_15398)
);

NOR2xp33_ASAP7_75t_L g15399 ( 
.A(n_15303),
.B(n_3264),
.Y(n_15399)
);

INVx1_ASAP7_75t_L g15400 ( 
.A(n_15349),
.Y(n_15400)
);

AOI211xp5_ASAP7_75t_L g15401 ( 
.A1(n_15286),
.A2(n_3267),
.B(n_3265),
.C(n_3266),
.Y(n_15401)
);

AOI221xp5_ASAP7_75t_L g15402 ( 
.A1(n_15350),
.A2(n_3269),
.B1(n_3266),
.B2(n_3268),
.C(n_3270),
.Y(n_15402)
);

OAI211xp5_ASAP7_75t_L g15403 ( 
.A1(n_15302),
.A2(n_3271),
.B(n_3268),
.C(n_3269),
.Y(n_15403)
);

AOI221xp5_ASAP7_75t_L g15404 ( 
.A1(n_15364),
.A2(n_3274),
.B1(n_3272),
.B2(n_3273),
.C(n_3275),
.Y(n_15404)
);

NAND2xp5_ASAP7_75t_SL g15405 ( 
.A(n_15336),
.B(n_3273),
.Y(n_15405)
);

OAI22xp5_ASAP7_75t_L g15406 ( 
.A1(n_15319),
.A2(n_3277),
.B1(n_3274),
.B2(n_3276),
.Y(n_15406)
);

INVx1_ASAP7_75t_SL g15407 ( 
.A(n_15283),
.Y(n_15407)
);

NOR2xp33_ASAP7_75t_L g15408 ( 
.A(n_15300),
.B(n_3276),
.Y(n_15408)
);

NAND2xp5_ASAP7_75t_L g15409 ( 
.A(n_15291),
.B(n_3277),
.Y(n_15409)
);

INVx1_ASAP7_75t_L g15410 ( 
.A(n_15298),
.Y(n_15410)
);

XOR2xp5_ASAP7_75t_L g15411 ( 
.A(n_15312),
.B(n_3278),
.Y(n_15411)
);

INVxp67_ASAP7_75t_SL g15412 ( 
.A(n_15308),
.Y(n_15412)
);

INVx1_ASAP7_75t_L g15413 ( 
.A(n_15310),
.Y(n_15413)
);

NOR2xp33_ASAP7_75t_SL g15414 ( 
.A(n_15287),
.B(n_3278),
.Y(n_15414)
);

INVx1_ASAP7_75t_SL g15415 ( 
.A(n_15367),
.Y(n_15415)
);

NOR2xp33_ASAP7_75t_L g15416 ( 
.A(n_15334),
.B(n_3279),
.Y(n_15416)
);

NOR2xp33_ASAP7_75t_SL g15417 ( 
.A(n_15296),
.B(n_3279),
.Y(n_15417)
);

INVx1_ASAP7_75t_L g15418 ( 
.A(n_15305),
.Y(n_15418)
);

INVx1_ASAP7_75t_L g15419 ( 
.A(n_15341),
.Y(n_15419)
);

INVx1_ASAP7_75t_L g15420 ( 
.A(n_15317),
.Y(n_15420)
);

NAND2xp5_ASAP7_75t_SL g15421 ( 
.A(n_15311),
.B(n_3280),
.Y(n_15421)
);

NAND4xp25_ASAP7_75t_L g15422 ( 
.A(n_15299),
.B(n_3282),
.C(n_3280),
.D(n_3281),
.Y(n_15422)
);

INVx2_ASAP7_75t_L g15423 ( 
.A(n_15321),
.Y(n_15423)
);

NOR2xp33_ASAP7_75t_L g15424 ( 
.A(n_15376),
.B(n_3281),
.Y(n_15424)
);

INVx1_ASAP7_75t_L g15425 ( 
.A(n_15290),
.Y(n_15425)
);

NOR2x1_ASAP7_75t_L g15426 ( 
.A(n_15284),
.B(n_3282),
.Y(n_15426)
);

NOR3x1_ASAP7_75t_L g15427 ( 
.A(n_15288),
.B(n_3285),
.C(n_3284),
.Y(n_15427)
);

OAI322xp33_ASAP7_75t_L g15428 ( 
.A1(n_15330),
.A2(n_3288),
.A3(n_3287),
.B1(n_3285),
.B2(n_3283),
.C1(n_3284),
.C2(n_3286),
.Y(n_15428)
);

INVx1_ASAP7_75t_L g15429 ( 
.A(n_15339),
.Y(n_15429)
);

AOI211xp5_ASAP7_75t_L g15430 ( 
.A1(n_15309),
.A2(n_3289),
.B(n_3283),
.C(n_3287),
.Y(n_15430)
);

INVx1_ASAP7_75t_L g15431 ( 
.A(n_15357),
.Y(n_15431)
);

NAND3xp33_ASAP7_75t_L g15432 ( 
.A(n_15282),
.B(n_3290),
.C(n_3291),
.Y(n_15432)
);

NAND4xp25_ASAP7_75t_L g15433 ( 
.A(n_15315),
.B(n_3292),
.C(n_3290),
.D(n_3291),
.Y(n_15433)
);

NAND4xp25_ASAP7_75t_L g15434 ( 
.A(n_15371),
.B(n_3294),
.C(n_3292),
.D(n_3293),
.Y(n_15434)
);

AOI221xp5_ASAP7_75t_L g15435 ( 
.A1(n_15332),
.A2(n_3295),
.B1(n_3293),
.B2(n_3294),
.C(n_3296),
.Y(n_15435)
);

NAND2xp33_ASAP7_75t_L g15436 ( 
.A(n_15316),
.B(n_3295),
.Y(n_15436)
);

INVx1_ASAP7_75t_L g15437 ( 
.A(n_15348),
.Y(n_15437)
);

NAND4xp25_ASAP7_75t_L g15438 ( 
.A(n_15362),
.B(n_3298),
.C(n_3296),
.D(n_3297),
.Y(n_15438)
);

NAND3xp33_ASAP7_75t_L g15439 ( 
.A(n_15329),
.B(n_3297),
.C(n_3298),
.Y(n_15439)
);

NOR3xp33_ASAP7_75t_L g15440 ( 
.A(n_15301),
.B(n_3299),
.C(n_3300),
.Y(n_15440)
);

INVx1_ASAP7_75t_L g15441 ( 
.A(n_15358),
.Y(n_15441)
);

NAND2xp5_ASAP7_75t_L g15442 ( 
.A(n_15352),
.B(n_3300),
.Y(n_15442)
);

NAND2xp5_ASAP7_75t_L g15443 ( 
.A(n_15359),
.B(n_3301),
.Y(n_15443)
);

NAND2xp5_ASAP7_75t_L g15444 ( 
.A(n_15344),
.B(n_3302),
.Y(n_15444)
);

AOI21xp5_ASAP7_75t_L g15445 ( 
.A1(n_15365),
.A2(n_3303),
.B(n_3304),
.Y(n_15445)
);

NAND2xp5_ASAP7_75t_L g15446 ( 
.A(n_15351),
.B(n_15363),
.Y(n_15446)
);

OA22x2_ASAP7_75t_L g15447 ( 
.A1(n_15335),
.A2(n_3305),
.B1(n_3303),
.B2(n_3304),
.Y(n_15447)
);

XNOR2x1_ASAP7_75t_L g15448 ( 
.A(n_15342),
.B(n_4117),
.Y(n_15448)
);

AOI221xp5_ASAP7_75t_L g15449 ( 
.A1(n_15360),
.A2(n_15331),
.B1(n_15343),
.B2(n_15346),
.C(n_15325),
.Y(n_15449)
);

NAND2xp5_ASAP7_75t_SL g15450 ( 
.A(n_15354),
.B(n_3305),
.Y(n_15450)
);

A2O1A1Ixp33_ASAP7_75t_L g15451 ( 
.A1(n_15369),
.A2(n_3308),
.B(n_3306),
.C(n_3307),
.Y(n_15451)
);

NOR2xp33_ASAP7_75t_L g15452 ( 
.A(n_15323),
.B(n_3306),
.Y(n_15452)
);

NAND2xp5_ASAP7_75t_L g15453 ( 
.A(n_15314),
.B(n_3307),
.Y(n_15453)
);

NAND2xp5_ASAP7_75t_L g15454 ( 
.A(n_15353),
.B(n_3308),
.Y(n_15454)
);

O2A1O1Ixp5_ASAP7_75t_L g15455 ( 
.A1(n_15340),
.A2(n_15361),
.B(n_15373),
.C(n_15294),
.Y(n_15455)
);

NOR3xp33_ASAP7_75t_L g15456 ( 
.A(n_15324),
.B(n_3309),
.C(n_3310),
.Y(n_15456)
);

AOI211xp5_ASAP7_75t_SL g15457 ( 
.A1(n_15337),
.A2(n_3312),
.B(n_3310),
.C(n_3311),
.Y(n_15457)
);

NOR2x1_ASAP7_75t_L g15458 ( 
.A(n_15285),
.B(n_3311),
.Y(n_15458)
);

NOR4xp25_ASAP7_75t_L g15459 ( 
.A(n_15356),
.B(n_15289),
.C(n_15322),
.D(n_15345),
.Y(n_15459)
);

INVx1_ASAP7_75t_L g15460 ( 
.A(n_15378),
.Y(n_15460)
);

NOR2x1_ASAP7_75t_L g15461 ( 
.A(n_15328),
.B(n_3313),
.Y(n_15461)
);

NAND5xp2_ASAP7_75t_L g15462 ( 
.A(n_15372),
.B(n_3315),
.C(n_3313),
.D(n_3314),
.E(n_3316),
.Y(n_15462)
);

INVx2_ASAP7_75t_L g15463 ( 
.A(n_15295),
.Y(n_15463)
);

AOI221xp5_ASAP7_75t_L g15464 ( 
.A1(n_15350),
.A2(n_3316),
.B1(n_3314),
.B2(n_3315),
.C(n_3317),
.Y(n_15464)
);

NOR2xp33_ASAP7_75t_L g15465 ( 
.A(n_15320),
.B(n_3318),
.Y(n_15465)
);

OAI322xp33_ASAP7_75t_L g15466 ( 
.A1(n_15366),
.A2(n_3325),
.A3(n_3324),
.B1(n_3322),
.B2(n_3319),
.C1(n_3320),
.C2(n_3323),
.Y(n_15466)
);

AOI21xp5_ASAP7_75t_L g15467 ( 
.A1(n_15368),
.A2(n_3319),
.B(n_3320),
.Y(n_15467)
);

INVx1_ASAP7_75t_L g15468 ( 
.A(n_15320),
.Y(n_15468)
);

INVx1_ASAP7_75t_L g15469 ( 
.A(n_15320),
.Y(n_15469)
);

INVx2_ASAP7_75t_L g15470 ( 
.A(n_15295),
.Y(n_15470)
);

NOR2xp33_ASAP7_75t_SL g15471 ( 
.A(n_15292),
.B(n_3322),
.Y(n_15471)
);

NOR3xp33_ASAP7_75t_L g15472 ( 
.A(n_15307),
.B(n_3323),
.C(n_3324),
.Y(n_15472)
);

OR2x2_ASAP7_75t_L g15473 ( 
.A(n_15295),
.B(n_3325),
.Y(n_15473)
);

NAND2xp5_ASAP7_75t_SL g15474 ( 
.A(n_15336),
.B(n_3326),
.Y(n_15474)
);

AOI22xp5_ASAP7_75t_L g15475 ( 
.A1(n_15326),
.A2(n_3328),
.B1(n_3326),
.B2(n_3327),
.Y(n_15475)
);

NOR3xp33_ASAP7_75t_L g15476 ( 
.A(n_15307),
.B(n_3327),
.C(n_3328),
.Y(n_15476)
);

NOR3xp33_ASAP7_75t_L g15477 ( 
.A(n_15379),
.B(n_3329),
.C(n_3330),
.Y(n_15477)
);

AOI21xp5_ASAP7_75t_L g15478 ( 
.A1(n_15454),
.A2(n_15411),
.B(n_15389),
.Y(n_15478)
);

INVxp67_ASAP7_75t_L g15479 ( 
.A(n_15394),
.Y(n_15479)
);

O2A1O1Ixp33_ASAP7_75t_L g15480 ( 
.A1(n_15388),
.A2(n_3331),
.B(n_3329),
.C(n_3330),
.Y(n_15480)
);

OAI21xp33_ASAP7_75t_L g15481 ( 
.A1(n_15462),
.A2(n_4107),
.B(n_4106),
.Y(n_15481)
);

NOR4xp75_ASAP7_75t_L g15482 ( 
.A(n_15384),
.B(n_3333),
.C(n_3331),
.D(n_3332),
.Y(n_15482)
);

INVx1_ASAP7_75t_L g15483 ( 
.A(n_15390),
.Y(n_15483)
);

NOR2xp33_ASAP7_75t_L g15484 ( 
.A(n_15468),
.B(n_3332),
.Y(n_15484)
);

HB1xp67_ASAP7_75t_L g15485 ( 
.A(n_15469),
.Y(n_15485)
);

HB1xp67_ASAP7_75t_L g15486 ( 
.A(n_15473),
.Y(n_15486)
);

INVx1_ASAP7_75t_L g15487 ( 
.A(n_15463),
.Y(n_15487)
);

INVx1_ASAP7_75t_L g15488 ( 
.A(n_15470),
.Y(n_15488)
);

INVx2_ASAP7_75t_L g15489 ( 
.A(n_15427),
.Y(n_15489)
);

NOR3xp33_ASAP7_75t_L g15490 ( 
.A(n_15381),
.B(n_3333),
.C(n_3334),
.Y(n_15490)
);

INVx2_ASAP7_75t_L g15491 ( 
.A(n_15380),
.Y(n_15491)
);

AOI221xp5_ASAP7_75t_L g15492 ( 
.A1(n_15466),
.A2(n_3337),
.B1(n_3335),
.B2(n_3336),
.C(n_3338),
.Y(n_15492)
);

AOI21xp33_ASAP7_75t_SL g15493 ( 
.A1(n_15465),
.A2(n_3335),
.B(n_3336),
.Y(n_15493)
);

NOR2x1_ASAP7_75t_L g15494 ( 
.A(n_15423),
.B(n_3338),
.Y(n_15494)
);

AND3x1_ASAP7_75t_L g15495 ( 
.A(n_15414),
.B(n_3339),
.C(n_3340),
.Y(n_15495)
);

INVxp67_ASAP7_75t_SL g15496 ( 
.A(n_15386),
.Y(n_15496)
);

AOI211xp5_ASAP7_75t_L g15497 ( 
.A1(n_15399),
.A2(n_3341),
.B(n_3339),
.C(n_3340),
.Y(n_15497)
);

NAND2xp5_ASAP7_75t_L g15498 ( 
.A(n_15418),
.B(n_15412),
.Y(n_15498)
);

NAND4xp75_ASAP7_75t_L g15499 ( 
.A(n_15441),
.B(n_3344),
.C(n_3342),
.D(n_3343),
.Y(n_15499)
);

NAND4xp75_ASAP7_75t_L g15500 ( 
.A(n_15400),
.B(n_3345),
.C(n_3342),
.D(n_3344),
.Y(n_15500)
);

O2A1O1Ixp33_ASAP7_75t_SL g15501 ( 
.A1(n_15451),
.A2(n_3353),
.B(n_3363),
.C(n_3345),
.Y(n_15501)
);

AOI211xp5_ASAP7_75t_SL g15502 ( 
.A1(n_15420),
.A2(n_3354),
.B(n_3365),
.C(n_3346),
.Y(n_15502)
);

AOI21xp5_ASAP7_75t_L g15503 ( 
.A1(n_15383),
.A2(n_3346),
.B(n_3347),
.Y(n_15503)
);

AND2x2_ASAP7_75t_L g15504 ( 
.A(n_15419),
.B(n_3348),
.Y(n_15504)
);

AOI222xp33_ASAP7_75t_L g15505 ( 
.A1(n_15405),
.A2(n_3350),
.B1(n_3352),
.B2(n_3348),
.C1(n_3349),
.C2(n_3351),
.Y(n_15505)
);

NOR2xp33_ASAP7_75t_L g15506 ( 
.A(n_15415),
.B(n_3349),
.Y(n_15506)
);

INVx1_ASAP7_75t_L g15507 ( 
.A(n_15474),
.Y(n_15507)
);

AND4x1_ASAP7_75t_L g15508 ( 
.A(n_15413),
.B(n_3354),
.C(n_3351),
.D(n_3353),
.Y(n_15508)
);

NAND4xp25_ASAP7_75t_SL g15509 ( 
.A(n_15435),
.B(n_3357),
.C(n_3355),
.D(n_3356),
.Y(n_15509)
);

NAND4xp25_ASAP7_75t_L g15510 ( 
.A(n_15449),
.B(n_3358),
.C(n_3355),
.D(n_3357),
.Y(n_15510)
);

NAND3xp33_ASAP7_75t_SL g15511 ( 
.A(n_15407),
.B(n_3358),
.C(n_3359),
.Y(n_15511)
);

AND2x2_ASAP7_75t_L g15512 ( 
.A(n_15458),
.B(n_15461),
.Y(n_15512)
);

INVx1_ASAP7_75t_SL g15513 ( 
.A(n_15448),
.Y(n_15513)
);

HB1xp67_ASAP7_75t_L g15514 ( 
.A(n_15387),
.Y(n_15514)
);

INVx1_ASAP7_75t_L g15515 ( 
.A(n_15446),
.Y(n_15515)
);

NAND2xp5_ASAP7_75t_L g15516 ( 
.A(n_15391),
.B(n_3359),
.Y(n_15516)
);

NAND2xp5_ASAP7_75t_L g15517 ( 
.A(n_15395),
.B(n_3360),
.Y(n_15517)
);

NAND4xp25_ASAP7_75t_L g15518 ( 
.A(n_15455),
.B(n_3367),
.C(n_3363),
.D(n_3366),
.Y(n_15518)
);

AOI21xp33_ASAP7_75t_SL g15519 ( 
.A1(n_15397),
.A2(n_3367),
.B(n_3368),
.Y(n_15519)
);

NAND2xp5_ASAP7_75t_SL g15520 ( 
.A(n_15393),
.B(n_3368),
.Y(n_15520)
);

NAND4xp75_ASAP7_75t_L g15521 ( 
.A(n_15429),
.B(n_3371),
.C(n_3369),
.D(n_3370),
.Y(n_15521)
);

INVx2_ASAP7_75t_SL g15522 ( 
.A(n_15426),
.Y(n_15522)
);

NAND4xp25_ASAP7_75t_L g15523 ( 
.A(n_15416),
.B(n_3373),
.C(n_3371),
.D(n_3372),
.Y(n_15523)
);

INVx1_ASAP7_75t_L g15524 ( 
.A(n_15409),
.Y(n_15524)
);

INVxp67_ASAP7_75t_L g15525 ( 
.A(n_15408),
.Y(n_15525)
);

AOI221xp5_ASAP7_75t_L g15526 ( 
.A1(n_15398),
.A2(n_3374),
.B1(n_3372),
.B2(n_3373),
.C(n_3375),
.Y(n_15526)
);

NAND3xp33_ASAP7_75t_SL g15527 ( 
.A(n_15425),
.B(n_3374),
.C(n_3375),
.Y(n_15527)
);

NOR3xp33_ASAP7_75t_L g15528 ( 
.A(n_15437),
.B(n_3376),
.C(n_3377),
.Y(n_15528)
);

INVx1_ASAP7_75t_L g15529 ( 
.A(n_15432),
.Y(n_15529)
);

AOI22xp33_ASAP7_75t_L g15530 ( 
.A1(n_15440),
.A2(n_3378),
.B1(n_3376),
.B2(n_3377),
.Y(n_15530)
);

INVx1_ASAP7_75t_L g15531 ( 
.A(n_15442),
.Y(n_15531)
);

NAND4xp75_ASAP7_75t_L g15532 ( 
.A(n_15445),
.B(n_3380),
.C(n_3378),
.D(n_3379),
.Y(n_15532)
);

AOI21xp5_ASAP7_75t_L g15533 ( 
.A1(n_15443),
.A2(n_3379),
.B(n_3380),
.Y(n_15533)
);

OAI221xp5_ASAP7_75t_L g15534 ( 
.A1(n_15422),
.A2(n_3383),
.B1(n_3381),
.B2(n_3382),
.C(n_3384),
.Y(n_15534)
);

INVxp67_ASAP7_75t_L g15535 ( 
.A(n_15424),
.Y(n_15535)
);

AND2x2_ASAP7_75t_L g15536 ( 
.A(n_15410),
.B(n_3381),
.Y(n_15536)
);

OAI211xp5_ASAP7_75t_L g15537 ( 
.A1(n_15396),
.A2(n_3385),
.B(n_3382),
.C(n_3383),
.Y(n_15537)
);

NAND4xp25_ASAP7_75t_L g15538 ( 
.A(n_15382),
.B(n_3387),
.C(n_3385),
.D(n_3386),
.Y(n_15538)
);

NOR2xp33_ASAP7_75t_L g15539 ( 
.A(n_15434),
.B(n_3386),
.Y(n_15539)
);

NAND2xp5_ASAP7_75t_L g15540 ( 
.A(n_15431),
.B(n_3388),
.Y(n_15540)
);

OR2x2_ASAP7_75t_L g15541 ( 
.A(n_15444),
.B(n_3388),
.Y(n_15541)
);

AOI21xp33_ASAP7_75t_L g15542 ( 
.A1(n_15460),
.A2(n_3389),
.B(n_3391),
.Y(n_15542)
);

NAND4xp25_ASAP7_75t_SL g15543 ( 
.A(n_15401),
.B(n_3392),
.C(n_3389),
.D(n_3391),
.Y(n_15543)
);

BUFx2_ASAP7_75t_L g15544 ( 
.A(n_15447),
.Y(n_15544)
);

INVx1_ASAP7_75t_L g15545 ( 
.A(n_15436),
.Y(n_15545)
);

NOR3xp33_ASAP7_75t_L g15546 ( 
.A(n_15428),
.B(n_3392),
.C(n_3393),
.Y(n_15546)
);

AO21x1_ASAP7_75t_L g15547 ( 
.A1(n_15452),
.A2(n_3393),
.B(n_3394),
.Y(n_15547)
);

AOI21xp33_ASAP7_75t_SL g15548 ( 
.A1(n_15472),
.A2(n_3394),
.B(n_3395),
.Y(n_15548)
);

NAND2xp5_ASAP7_75t_L g15549 ( 
.A(n_15467),
.B(n_3395),
.Y(n_15549)
);

NAND4xp25_ASAP7_75t_L g15550 ( 
.A(n_15402),
.B(n_3399),
.C(n_3397),
.D(n_3398),
.Y(n_15550)
);

NAND2xp5_ASAP7_75t_SL g15551 ( 
.A(n_15464),
.B(n_3397),
.Y(n_15551)
);

NAND2xp5_ASAP7_75t_L g15552 ( 
.A(n_15459),
.B(n_3398),
.Y(n_15552)
);

NAND3xp33_ASAP7_75t_SL g15553 ( 
.A(n_15476),
.B(n_3399),
.C(n_3400),
.Y(n_15553)
);

NAND2xp5_ASAP7_75t_L g15554 ( 
.A(n_15457),
.B(n_3400),
.Y(n_15554)
);

NOR4xp25_ASAP7_75t_L g15555 ( 
.A(n_15438),
.B(n_3403),
.C(n_3401),
.D(n_3402),
.Y(n_15555)
);

NOR2x1_ASAP7_75t_L g15556 ( 
.A(n_15433),
.B(n_3401),
.Y(n_15556)
);

NAND4xp25_ASAP7_75t_L g15557 ( 
.A(n_15430),
.B(n_15471),
.C(n_15404),
.D(n_15417),
.Y(n_15557)
);

XNOR2xp5_ASAP7_75t_L g15558 ( 
.A(n_15439),
.B(n_3402),
.Y(n_15558)
);

OAI21xp5_ASAP7_75t_SL g15559 ( 
.A1(n_15392),
.A2(n_3403),
.B(n_3404),
.Y(n_15559)
);

AOI211xp5_ASAP7_75t_L g15560 ( 
.A1(n_15385),
.A2(n_3406),
.B(n_3404),
.C(n_3405),
.Y(n_15560)
);

NAND5xp2_ASAP7_75t_L g15561 ( 
.A(n_15456),
.B(n_3408),
.C(n_3406),
.D(n_3407),
.E(n_3409),
.Y(n_15561)
);

NAND4xp75_ASAP7_75t_L g15562 ( 
.A(n_15487),
.B(n_15453),
.C(n_15450),
.D(n_15421),
.Y(n_15562)
);

OAI322xp33_ASAP7_75t_L g15563 ( 
.A1(n_15488),
.A2(n_15406),
.A3(n_15475),
.B1(n_15403),
.B2(n_3410),
.C1(n_3413),
.C2(n_3412),
.Y(n_15563)
);

NAND5xp2_ASAP7_75t_L g15564 ( 
.A(n_15512),
.B(n_3425),
.C(n_3433),
.D(n_3417),
.E(n_3408),
.Y(n_15564)
);

NAND4xp75_ASAP7_75t_L g15565 ( 
.A(n_15494),
.B(n_3411),
.C(n_3409),
.D(n_3410),
.Y(n_15565)
);

NOR2xp67_ASAP7_75t_L g15566 ( 
.A(n_15511),
.B(n_3413),
.Y(n_15566)
);

O2A1O1Ixp33_ASAP7_75t_L g15567 ( 
.A1(n_15485),
.A2(n_3415),
.B(n_3411),
.C(n_3414),
.Y(n_15567)
);

NOR3x1_ASAP7_75t_L g15568 ( 
.A(n_15521),
.B(n_3414),
.C(n_3415),
.Y(n_15568)
);

NOR3x1_ASAP7_75t_L g15569 ( 
.A(n_15552),
.B(n_3416),
.C(n_3417),
.Y(n_15569)
);

AO22x2_ASAP7_75t_L g15570 ( 
.A1(n_15483),
.A2(n_15522),
.B1(n_15491),
.B2(n_15507),
.Y(n_15570)
);

NOR3xp33_ASAP7_75t_SL g15571 ( 
.A(n_15498),
.B(n_3418),
.C(n_3419),
.Y(n_15571)
);

NOR3xp33_ASAP7_75t_SL g15572 ( 
.A(n_15515),
.B(n_3418),
.C(n_3419),
.Y(n_15572)
);

NAND2xp5_ASAP7_75t_L g15573 ( 
.A(n_15486),
.B(n_4117),
.Y(n_15573)
);

NAND3xp33_ASAP7_75t_L g15574 ( 
.A(n_15479),
.B(n_3420),
.C(n_3421),
.Y(n_15574)
);

NOR2x1_ASAP7_75t_L g15575 ( 
.A(n_15545),
.B(n_3421),
.Y(n_15575)
);

NOR2x1_ASAP7_75t_L g15576 ( 
.A(n_15489),
.B(n_3422),
.Y(n_15576)
);

AND2x2_ASAP7_75t_L g15577 ( 
.A(n_15544),
.B(n_3422),
.Y(n_15577)
);

AND2x2_ASAP7_75t_SL g15578 ( 
.A(n_15495),
.B(n_3423),
.Y(n_15578)
);

NAND2xp5_ASAP7_75t_L g15579 ( 
.A(n_15496),
.B(n_15513),
.Y(n_15579)
);

INVx1_ASAP7_75t_L g15580 ( 
.A(n_15504),
.Y(n_15580)
);

NAND2xp5_ASAP7_75t_L g15581 ( 
.A(n_15478),
.B(n_4121),
.Y(n_15581)
);

AND2x4_ASAP7_75t_L g15582 ( 
.A(n_15482),
.B(n_3423),
.Y(n_15582)
);

OAI21xp33_ASAP7_75t_SL g15583 ( 
.A1(n_15505),
.A2(n_3424),
.B(n_3426),
.Y(n_15583)
);

NAND4xp25_ASAP7_75t_L g15584 ( 
.A(n_15561),
.B(n_4122),
.C(n_3427),
.D(n_3424),
.Y(n_15584)
);

NOR2xp33_ASAP7_75t_L g15585 ( 
.A(n_15525),
.B(n_3426),
.Y(n_15585)
);

NOR3xp33_ASAP7_75t_L g15586 ( 
.A(n_15524),
.B(n_3427),
.C(n_3428),
.Y(n_15586)
);

AND5x1_ASAP7_75t_L g15587 ( 
.A(n_15546),
.B(n_3430),
.C(n_3428),
.D(n_3429),
.E(n_3431),
.Y(n_15587)
);

INVx1_ASAP7_75t_L g15588 ( 
.A(n_15536),
.Y(n_15588)
);

AND2x4_ASAP7_75t_L g15589 ( 
.A(n_15529),
.B(n_3429),
.Y(n_15589)
);

INVx1_ASAP7_75t_L g15590 ( 
.A(n_15547),
.Y(n_15590)
);

NOR2xp33_ASAP7_75t_L g15591 ( 
.A(n_15535),
.B(n_3430),
.Y(n_15591)
);

AOI31xp33_ASAP7_75t_L g15592 ( 
.A1(n_15514),
.A2(n_3434),
.A3(n_3435),
.B(n_3432),
.Y(n_15592)
);

INVx1_ASAP7_75t_L g15593 ( 
.A(n_15540),
.Y(n_15593)
);

NAND2x1_ASAP7_75t_SL g15594 ( 
.A(n_15506),
.B(n_3431),
.Y(n_15594)
);

NOR3xp33_ASAP7_75t_L g15595 ( 
.A(n_15531),
.B(n_3432),
.C(n_3434),
.Y(n_15595)
);

OAI22xp5_ASAP7_75t_L g15596 ( 
.A1(n_15530),
.A2(n_3437),
.B1(n_3435),
.B2(n_3436),
.Y(n_15596)
);

INVx1_ASAP7_75t_L g15597 ( 
.A(n_15541),
.Y(n_15597)
);

NAND2xp5_ASAP7_75t_L g15598 ( 
.A(n_15481),
.B(n_4116),
.Y(n_15598)
);

NAND2xp5_ASAP7_75t_L g15599 ( 
.A(n_15484),
.B(n_4116),
.Y(n_15599)
);

NAND2xp5_ASAP7_75t_L g15600 ( 
.A(n_15493),
.B(n_4119),
.Y(n_15600)
);

INVx1_ASAP7_75t_L g15601 ( 
.A(n_15554),
.Y(n_15601)
);

NOR2x1_ASAP7_75t_L g15602 ( 
.A(n_15527),
.B(n_3437),
.Y(n_15602)
);

NOR2x1p5_ASAP7_75t_L g15603 ( 
.A(n_15532),
.B(n_3438),
.Y(n_15603)
);

NOR2x1p5_ASAP7_75t_SL g15604 ( 
.A(n_15499),
.B(n_3438),
.Y(n_15604)
);

AOI211x1_ASAP7_75t_L g15605 ( 
.A1(n_15537),
.A2(n_3441),
.B(n_3439),
.C(n_3440),
.Y(n_15605)
);

NAND2xp5_ASAP7_75t_L g15606 ( 
.A(n_15556),
.B(n_4122),
.Y(n_15606)
);

OAI211xp5_ASAP7_75t_SL g15607 ( 
.A1(n_15520),
.A2(n_3442),
.B(n_3439),
.C(n_3440),
.Y(n_15607)
);

NOR2x1_ASAP7_75t_L g15608 ( 
.A(n_15500),
.B(n_3443),
.Y(n_15608)
);

NAND5xp2_ASAP7_75t_L g15609 ( 
.A(n_15559),
.B(n_3460),
.C(n_3468),
.D(n_3452),
.E(n_3444),
.Y(n_15609)
);

OAI21xp5_ASAP7_75t_L g15610 ( 
.A1(n_15533),
.A2(n_3445),
.B(n_3446),
.Y(n_15610)
);

NAND3xp33_ASAP7_75t_L g15611 ( 
.A(n_15477),
.B(n_3445),
.C(n_3446),
.Y(n_15611)
);

AND2x2_ASAP7_75t_L g15612 ( 
.A(n_15555),
.B(n_3447),
.Y(n_15612)
);

NAND2x1p5_ASAP7_75t_L g15613 ( 
.A(n_15508),
.B(n_3447),
.Y(n_15613)
);

AND2x2_ASAP7_75t_L g15614 ( 
.A(n_15502),
.B(n_3448),
.Y(n_15614)
);

NAND2xp5_ASAP7_75t_L g15615 ( 
.A(n_15503),
.B(n_4106),
.Y(n_15615)
);

NOR2x1_ASAP7_75t_L g15616 ( 
.A(n_15523),
.B(n_3448),
.Y(n_15616)
);

NOR2x1_ASAP7_75t_L g15617 ( 
.A(n_15518),
.B(n_3449),
.Y(n_15617)
);

NOR3xp33_ASAP7_75t_L g15618 ( 
.A(n_15553),
.B(n_3450),
.C(n_3451),
.Y(n_15618)
);

INVx1_ASAP7_75t_L g15619 ( 
.A(n_15516),
.Y(n_15619)
);

NOR3xp33_ASAP7_75t_L g15620 ( 
.A(n_15517),
.B(n_3450),
.C(n_3451),
.Y(n_15620)
);

NAND2xp5_ASAP7_75t_L g15621 ( 
.A(n_15539),
.B(n_15519),
.Y(n_15621)
);

AND2x4_ASAP7_75t_L g15622 ( 
.A(n_15549),
.B(n_3452),
.Y(n_15622)
);

NAND4xp25_ASAP7_75t_L g15623 ( 
.A(n_15526),
.B(n_4121),
.C(n_3455),
.D(n_3453),
.Y(n_15623)
);

NAND5xp2_ASAP7_75t_L g15624 ( 
.A(n_15560),
.B(n_3471),
.C(n_3479),
.D(n_3462),
.E(n_3454),
.Y(n_15624)
);

NOR2xp33_ASAP7_75t_L g15625 ( 
.A(n_15510),
.B(n_3454),
.Y(n_15625)
);

INVx1_ASAP7_75t_L g15626 ( 
.A(n_15558),
.Y(n_15626)
);

NOR3x1_ASAP7_75t_L g15627 ( 
.A(n_15538),
.B(n_3455),
.C(n_3456),
.Y(n_15627)
);

NOR2xp33_ASAP7_75t_L g15628 ( 
.A(n_15548),
.B(n_3457),
.Y(n_15628)
);

INVx1_ASAP7_75t_L g15629 ( 
.A(n_15501),
.Y(n_15629)
);

O2A1O1Ixp33_ASAP7_75t_L g15630 ( 
.A1(n_15480),
.A2(n_3460),
.B(n_3458),
.C(n_3459),
.Y(n_15630)
);

AOI21xp5_ASAP7_75t_L g15631 ( 
.A1(n_15542),
.A2(n_3461),
.B(n_3462),
.Y(n_15631)
);

NOR3xp33_ASAP7_75t_L g15632 ( 
.A(n_15490),
.B(n_3461),
.C(n_3463),
.Y(n_15632)
);

NOR3xp33_ASAP7_75t_L g15633 ( 
.A(n_15557),
.B(n_3463),
.C(n_3464),
.Y(n_15633)
);

NAND4xp25_ASAP7_75t_L g15634 ( 
.A(n_15497),
.B(n_15492),
.C(n_15528),
.D(n_15550),
.Y(n_15634)
);

INVx1_ASAP7_75t_L g15635 ( 
.A(n_15534),
.Y(n_15635)
);

NAND3xp33_ASAP7_75t_L g15636 ( 
.A(n_15551),
.B(n_3465),
.C(n_3466),
.Y(n_15636)
);

NAND3xp33_ASAP7_75t_L g15637 ( 
.A(n_15543),
.B(n_3465),
.C(n_3467),
.Y(n_15637)
);

INVx2_ASAP7_75t_SL g15638 ( 
.A(n_15509),
.Y(n_15638)
);

NOR2xp67_ASAP7_75t_L g15639 ( 
.A(n_15511),
.B(n_3469),
.Y(n_15639)
);

INVx1_ASAP7_75t_SL g15640 ( 
.A(n_15512),
.Y(n_15640)
);

NOR3xp33_ASAP7_75t_L g15641 ( 
.A(n_15485),
.B(n_3467),
.C(n_3469),
.Y(n_15641)
);

INVx2_ASAP7_75t_SL g15642 ( 
.A(n_15485),
.Y(n_15642)
);

OAI211xp5_ASAP7_75t_SL g15643 ( 
.A1(n_15487),
.A2(n_3472),
.B(n_3470),
.C(n_3471),
.Y(n_15643)
);

INVx1_ASAP7_75t_L g15644 ( 
.A(n_15486),
.Y(n_15644)
);

INVx2_ASAP7_75t_SL g15645 ( 
.A(n_15485),
.Y(n_15645)
);

INVx1_ASAP7_75t_L g15646 ( 
.A(n_15486),
.Y(n_15646)
);

CKINVDCx20_ASAP7_75t_R g15647 ( 
.A(n_15486),
.Y(n_15647)
);

INVx1_ASAP7_75t_L g15648 ( 
.A(n_15486),
.Y(n_15648)
);

OAI22xp5_ASAP7_75t_L g15649 ( 
.A1(n_15515),
.A2(n_3473),
.B1(n_3470),
.B2(n_3472),
.Y(n_15649)
);

INVxp33_ASAP7_75t_L g15650 ( 
.A(n_15485),
.Y(n_15650)
);

INVx1_ASAP7_75t_L g15651 ( 
.A(n_15486),
.Y(n_15651)
);

INVx2_ASAP7_75t_SL g15652 ( 
.A(n_15642),
.Y(n_15652)
);

NAND4xp25_ASAP7_75t_L g15653 ( 
.A(n_15644),
.B(n_15646),
.C(n_15651),
.D(n_15648),
.Y(n_15653)
);

NOR2x1_ASAP7_75t_L g15654 ( 
.A(n_15647),
.B(n_3473),
.Y(n_15654)
);

NAND2xp5_ASAP7_75t_L g15655 ( 
.A(n_15645),
.B(n_3474),
.Y(n_15655)
);

NOR4xp75_ASAP7_75t_L g15656 ( 
.A(n_15579),
.B(n_3476),
.C(n_3474),
.D(n_3475),
.Y(n_15656)
);

NOR3xp33_ASAP7_75t_L g15657 ( 
.A(n_15640),
.B(n_3476),
.C(n_3477),
.Y(n_15657)
);

OAI211xp5_ASAP7_75t_L g15658 ( 
.A1(n_15590),
.A2(n_3480),
.B(n_3481),
.C(n_3478),
.Y(n_15658)
);

NOR3xp33_ASAP7_75t_L g15659 ( 
.A(n_15597),
.B(n_15588),
.C(n_15580),
.Y(n_15659)
);

NAND3xp33_ASAP7_75t_L g15660 ( 
.A(n_15650),
.B(n_3477),
.C(n_3478),
.Y(n_15660)
);

NAND2xp5_ASAP7_75t_L g15661 ( 
.A(n_15570),
.B(n_3482),
.Y(n_15661)
);

NAND2xp5_ASAP7_75t_L g15662 ( 
.A(n_15570),
.B(n_3482),
.Y(n_15662)
);

NAND3xp33_ASAP7_75t_L g15663 ( 
.A(n_15601),
.B(n_15593),
.C(n_15619),
.Y(n_15663)
);

AND2x2_ASAP7_75t_L g15664 ( 
.A(n_15577),
.B(n_15578),
.Y(n_15664)
);

NOR3xp33_ASAP7_75t_L g15665 ( 
.A(n_15626),
.B(n_3483),
.C(n_3484),
.Y(n_15665)
);

NAND3xp33_ASAP7_75t_L g15666 ( 
.A(n_15581),
.B(n_3483),
.C(n_3484),
.Y(n_15666)
);

HB1xp67_ASAP7_75t_L g15667 ( 
.A(n_15566),
.Y(n_15667)
);

NOR3xp33_ASAP7_75t_L g15668 ( 
.A(n_15562),
.B(n_3485),
.C(n_3486),
.Y(n_15668)
);

NAND4xp75_ASAP7_75t_L g15669 ( 
.A(n_15576),
.B(n_3487),
.C(n_3485),
.D(n_3486),
.Y(n_15669)
);

NAND2xp5_ASAP7_75t_L g15670 ( 
.A(n_15594),
.B(n_3487),
.Y(n_15670)
);

INVx1_ASAP7_75t_L g15671 ( 
.A(n_15613),
.Y(n_15671)
);

NAND3xp33_ASAP7_75t_SL g15672 ( 
.A(n_15621),
.B(n_15606),
.C(n_15620),
.Y(n_15672)
);

NOR4xp25_ASAP7_75t_L g15673 ( 
.A(n_15629),
.B(n_3490),
.C(n_3488),
.D(n_3489),
.Y(n_15673)
);

NAND2xp5_ASAP7_75t_L g15674 ( 
.A(n_15639),
.B(n_3488),
.Y(n_15674)
);

OAI21xp33_ASAP7_75t_L g15675 ( 
.A1(n_15609),
.A2(n_3489),
.B(n_3490),
.Y(n_15675)
);

NAND4xp25_ASAP7_75t_L g15676 ( 
.A(n_15569),
.B(n_3493),
.C(n_3491),
.D(n_3492),
.Y(n_15676)
);

NOR4xp25_ASAP7_75t_L g15677 ( 
.A(n_15635),
.B(n_15638),
.C(n_15563),
.D(n_15583),
.Y(n_15677)
);

INVx2_ASAP7_75t_SL g15678 ( 
.A(n_15575),
.Y(n_15678)
);

NAND3xp33_ASAP7_75t_L g15679 ( 
.A(n_15572),
.B(n_3491),
.C(n_3492),
.Y(n_15679)
);

INVxp33_ASAP7_75t_L g15680 ( 
.A(n_15573),
.Y(n_15680)
);

OAI21xp33_ASAP7_75t_SL g15681 ( 
.A1(n_15584),
.A2(n_3495),
.B(n_3494),
.Y(n_15681)
);

NOR3xp33_ASAP7_75t_L g15682 ( 
.A(n_15599),
.B(n_3493),
.C(n_3494),
.Y(n_15682)
);

NOR2x1_ASAP7_75t_L g15683 ( 
.A(n_15565),
.B(n_3495),
.Y(n_15683)
);

OAI211xp5_ASAP7_75t_L g15684 ( 
.A1(n_15612),
.A2(n_3498),
.B(n_3499),
.C(n_3497),
.Y(n_15684)
);

NOR3xp33_ASAP7_75t_L g15685 ( 
.A(n_15615),
.B(n_3496),
.C(n_3497),
.Y(n_15685)
);

NAND3xp33_ASAP7_75t_L g15686 ( 
.A(n_15622),
.B(n_15641),
.C(n_15571),
.Y(n_15686)
);

NOR2xp33_ASAP7_75t_L g15687 ( 
.A(n_15564),
.B(n_3496),
.Y(n_15687)
);

NAND2xp5_ASAP7_75t_L g15688 ( 
.A(n_15582),
.B(n_3498),
.Y(n_15688)
);

NAND2xp5_ASAP7_75t_SL g15689 ( 
.A(n_15582),
.B(n_3499),
.Y(n_15689)
);

NOR2xp67_ASAP7_75t_L g15690 ( 
.A(n_15574),
.B(n_3500),
.Y(n_15690)
);

NAND3xp33_ASAP7_75t_L g15691 ( 
.A(n_15622),
.B(n_3500),
.C(n_3501),
.Y(n_15691)
);

AND2x2_ASAP7_75t_L g15692 ( 
.A(n_15614),
.B(n_3501),
.Y(n_15692)
);

AOI211x1_ASAP7_75t_L g15693 ( 
.A1(n_15610),
.A2(n_3504),
.B(n_3502),
.C(n_3503),
.Y(n_15693)
);

AND2x2_ASAP7_75t_L g15694 ( 
.A(n_15602),
.B(n_15617),
.Y(n_15694)
);

INVx1_ASAP7_75t_L g15695 ( 
.A(n_15604),
.Y(n_15695)
);

NOR3x1_ASAP7_75t_L g15696 ( 
.A(n_15636),
.B(n_3502),
.C(n_3503),
.Y(n_15696)
);

NOR3x1_ASAP7_75t_L g15697 ( 
.A(n_15637),
.B(n_3504),
.C(n_3505),
.Y(n_15697)
);

OAI211xp5_ASAP7_75t_L g15698 ( 
.A1(n_15598),
.A2(n_3508),
.B(n_3509),
.C(n_3507),
.Y(n_15698)
);

INVxp67_ASAP7_75t_SL g15699 ( 
.A(n_15591),
.Y(n_15699)
);

NOR2x1_ASAP7_75t_L g15700 ( 
.A(n_15603),
.B(n_15608),
.Y(n_15700)
);

NAND3xp33_ASAP7_75t_L g15701 ( 
.A(n_15628),
.B(n_3506),
.C(n_3507),
.Y(n_15701)
);

NOR4xp25_ASAP7_75t_L g15702 ( 
.A(n_15634),
.B(n_3509),
.C(n_3506),
.D(n_3508),
.Y(n_15702)
);

NOR2x1_ASAP7_75t_L g15703 ( 
.A(n_15607),
.B(n_3510),
.Y(n_15703)
);

NOR2x1_ASAP7_75t_L g15704 ( 
.A(n_15611),
.B(n_3510),
.Y(n_15704)
);

NAND3xp33_ASAP7_75t_L g15705 ( 
.A(n_15595),
.B(n_3511),
.C(n_3512),
.Y(n_15705)
);

CKINVDCx5p33_ASAP7_75t_R g15706 ( 
.A(n_15625),
.Y(n_15706)
);

NAND2xp5_ASAP7_75t_L g15707 ( 
.A(n_15616),
.B(n_3511),
.Y(n_15707)
);

NAND4xp25_ASAP7_75t_L g15708 ( 
.A(n_15568),
.B(n_3514),
.C(n_3512),
.D(n_3513),
.Y(n_15708)
);

NOR3xp33_ASAP7_75t_L g15709 ( 
.A(n_15600),
.B(n_15643),
.C(n_15586),
.Y(n_15709)
);

NAND2x1p5_ASAP7_75t_L g15710 ( 
.A(n_15587),
.B(n_15627),
.Y(n_15710)
);

NOR2x1_ASAP7_75t_L g15711 ( 
.A(n_15592),
.B(n_3515),
.Y(n_15711)
);

NOR2xp33_ASAP7_75t_L g15712 ( 
.A(n_15624),
.B(n_3515),
.Y(n_15712)
);

INVx1_ASAP7_75t_L g15713 ( 
.A(n_15589),
.Y(n_15713)
);

NOR3xp33_ASAP7_75t_L g15714 ( 
.A(n_15585),
.B(n_3516),
.C(n_3517),
.Y(n_15714)
);

AOI211xp5_ASAP7_75t_L g15715 ( 
.A1(n_15567),
.A2(n_3518),
.B(n_3516),
.C(n_3517),
.Y(n_15715)
);

NOR2xp33_ASAP7_75t_L g15716 ( 
.A(n_15623),
.B(n_3518),
.Y(n_15716)
);

NOR2x1_ASAP7_75t_L g15717 ( 
.A(n_15649),
.B(n_15630),
.Y(n_15717)
);

NOR4xp25_ASAP7_75t_L g15718 ( 
.A(n_15596),
.B(n_15605),
.C(n_15618),
.D(n_15631),
.Y(n_15718)
);

NAND3xp33_ASAP7_75t_L g15719 ( 
.A(n_15633),
.B(n_3519),
.C(n_3520),
.Y(n_15719)
);

NOR2xp67_ASAP7_75t_L g15720 ( 
.A(n_15589),
.B(n_3519),
.Y(n_15720)
);

INVx1_ASAP7_75t_L g15721 ( 
.A(n_15632),
.Y(n_15721)
);

NOR4xp25_ASAP7_75t_L g15722 ( 
.A(n_15642),
.B(n_3523),
.C(n_3521),
.D(n_3522),
.Y(n_15722)
);

NOR3xp33_ASAP7_75t_L g15723 ( 
.A(n_15642),
.B(n_3521),
.C(n_3522),
.Y(n_15723)
);

INVxp33_ASAP7_75t_SL g15724 ( 
.A(n_15640),
.Y(n_15724)
);

OAI211xp5_ASAP7_75t_SL g15725 ( 
.A1(n_15644),
.A2(n_4103),
.B(n_4104),
.C(n_4102),
.Y(n_15725)
);

INVx1_ASAP7_75t_L g15726 ( 
.A(n_15647),
.Y(n_15726)
);

AOI211xp5_ASAP7_75t_L g15727 ( 
.A1(n_15650),
.A2(n_3525),
.B(n_3523),
.C(n_3524),
.Y(n_15727)
);

INVx1_ASAP7_75t_L g15728 ( 
.A(n_15647),
.Y(n_15728)
);

NOR3x1_ASAP7_75t_L g15729 ( 
.A(n_15642),
.B(n_3525),
.C(n_3526),
.Y(n_15729)
);

NAND3xp33_ASAP7_75t_SL g15730 ( 
.A(n_15647),
.B(n_3534),
.C(n_3526),
.Y(n_15730)
);

NAND3xp33_ASAP7_75t_L g15731 ( 
.A(n_15642),
.B(n_3527),
.C(n_3528),
.Y(n_15731)
);

NAND4xp25_ASAP7_75t_SL g15732 ( 
.A(n_15640),
.B(n_3529),
.C(n_3527),
.D(n_3528),
.Y(n_15732)
);

NAND2xp5_ASAP7_75t_L g15733 ( 
.A(n_15642),
.B(n_3529),
.Y(n_15733)
);

NOR3xp33_ASAP7_75t_L g15734 ( 
.A(n_15642),
.B(n_3530),
.C(n_3531),
.Y(n_15734)
);

NOR3xp33_ASAP7_75t_L g15735 ( 
.A(n_15642),
.B(n_3531),
.C(n_3532),
.Y(n_15735)
);

NOR3xp33_ASAP7_75t_L g15736 ( 
.A(n_15642),
.B(n_3532),
.C(n_3533),
.Y(n_15736)
);

OAI21xp33_ASAP7_75t_L g15737 ( 
.A1(n_15650),
.A2(n_3533),
.B(n_3534),
.Y(n_15737)
);

NAND3x1_ASAP7_75t_L g15738 ( 
.A(n_15644),
.B(n_3535),
.C(n_3536),
.Y(n_15738)
);

NAND2xp33_ASAP7_75t_SL g15739 ( 
.A(n_15650),
.B(n_4099),
.Y(n_15739)
);

NAND4xp25_ASAP7_75t_L g15740 ( 
.A(n_15644),
.B(n_3538),
.C(n_3535),
.D(n_3537),
.Y(n_15740)
);

NOR2x1_ASAP7_75t_L g15741 ( 
.A(n_15647),
.B(n_3537),
.Y(n_15741)
);

NAND2xp5_ASAP7_75t_L g15742 ( 
.A(n_15642),
.B(n_3538),
.Y(n_15742)
);

NAND4xp25_ASAP7_75t_L g15743 ( 
.A(n_15644),
.B(n_3541),
.C(n_3539),
.D(n_3540),
.Y(n_15743)
);

NAND3xp33_ASAP7_75t_L g15744 ( 
.A(n_15642),
.B(n_3539),
.C(n_3540),
.Y(n_15744)
);

NOR3xp33_ASAP7_75t_L g15745 ( 
.A(n_15642),
.B(n_3541),
.C(n_3542),
.Y(n_15745)
);

AND2x2_ASAP7_75t_L g15746 ( 
.A(n_15650),
.B(n_3543),
.Y(n_15746)
);

NOR2xp33_ASAP7_75t_L g15747 ( 
.A(n_15650),
.B(n_3543),
.Y(n_15747)
);

OAI211xp5_ASAP7_75t_SL g15748 ( 
.A1(n_15644),
.A2(n_4113),
.B(n_4114),
.C(n_4105),
.Y(n_15748)
);

NOR3xp33_ASAP7_75t_L g15749 ( 
.A(n_15642),
.B(n_3545),
.C(n_3546),
.Y(n_15749)
);

NOR3xp33_ASAP7_75t_L g15750 ( 
.A(n_15642),
.B(n_3545),
.C(n_3546),
.Y(n_15750)
);

INVx1_ASAP7_75t_L g15751 ( 
.A(n_15647),
.Y(n_15751)
);

NOR3xp33_ASAP7_75t_L g15752 ( 
.A(n_15642),
.B(n_3547),
.C(n_3548),
.Y(n_15752)
);

INVxp33_ASAP7_75t_SL g15753 ( 
.A(n_15640),
.Y(n_15753)
);

NAND2xp5_ASAP7_75t_L g15754 ( 
.A(n_15642),
.B(n_3547),
.Y(n_15754)
);

NOR2x1_ASAP7_75t_L g15755 ( 
.A(n_15647),
.B(n_3549),
.Y(n_15755)
);

NOR2x1_ASAP7_75t_L g15756 ( 
.A(n_15647),
.B(n_3549),
.Y(n_15756)
);

NOR2x1_ASAP7_75t_L g15757 ( 
.A(n_15647),
.B(n_3550),
.Y(n_15757)
);

NOR2xp33_ASAP7_75t_L g15758 ( 
.A(n_15650),
.B(n_3550),
.Y(n_15758)
);

BUFx6f_ASAP7_75t_L g15759 ( 
.A(n_15652),
.Y(n_15759)
);

OAI211xp5_ASAP7_75t_L g15760 ( 
.A1(n_15726),
.A2(n_3553),
.B(n_3551),
.C(n_3552),
.Y(n_15760)
);

NOR4xp25_ASAP7_75t_L g15761 ( 
.A(n_15653),
.B(n_3554),
.C(n_3551),
.D(n_3553),
.Y(n_15761)
);

INVxp67_ASAP7_75t_L g15762 ( 
.A(n_15728),
.Y(n_15762)
);

INVx1_ASAP7_75t_L g15763 ( 
.A(n_15751),
.Y(n_15763)
);

AOI221xp5_ASAP7_75t_L g15764 ( 
.A1(n_15724),
.A2(n_3556),
.B1(n_3554),
.B2(n_3555),
.C(n_3558),
.Y(n_15764)
);

AOI221xp5_ASAP7_75t_L g15765 ( 
.A1(n_15753),
.A2(n_3558),
.B1(n_3555),
.B2(n_3556),
.C(n_3559),
.Y(n_15765)
);

AOI221xp5_ASAP7_75t_L g15766 ( 
.A1(n_15677),
.A2(n_3561),
.B1(n_3559),
.B2(n_3560),
.C(n_3562),
.Y(n_15766)
);

AOI221xp5_ASAP7_75t_L g15767 ( 
.A1(n_15695),
.A2(n_3563),
.B1(n_3560),
.B2(n_3561),
.C(n_3564),
.Y(n_15767)
);

OAI321xp33_ASAP7_75t_L g15768 ( 
.A1(n_15710),
.A2(n_3565),
.A3(n_3567),
.B1(n_3563),
.B2(n_3564),
.C(n_3566),
.Y(n_15768)
);

INVx1_ASAP7_75t_L g15769 ( 
.A(n_15661),
.Y(n_15769)
);

NAND2xp5_ASAP7_75t_SL g15770 ( 
.A(n_15720),
.B(n_3565),
.Y(n_15770)
);

AOI221xp5_ASAP7_75t_L g15771 ( 
.A1(n_15659),
.A2(n_3568),
.B1(n_3566),
.B2(n_3567),
.C(n_3569),
.Y(n_15771)
);

OAI211xp5_ASAP7_75t_SL g15772 ( 
.A1(n_15662),
.A2(n_3571),
.B(n_3572),
.C(n_3570),
.Y(n_15772)
);

OAI22xp5_ASAP7_75t_L g15773 ( 
.A1(n_15663),
.A2(n_3579),
.B1(n_3587),
.B2(n_3568),
.Y(n_15773)
);

OAI211xp5_ASAP7_75t_SL g15774 ( 
.A1(n_15713),
.A2(n_3573),
.B(n_3574),
.C(n_3571),
.Y(n_15774)
);

AOI22xp5_ASAP7_75t_L g15775 ( 
.A1(n_15664),
.A2(n_15687),
.B1(n_15671),
.B2(n_15692),
.Y(n_15775)
);

NAND2xp5_ASAP7_75t_L g15776 ( 
.A(n_15667),
.B(n_3570),
.Y(n_15776)
);

HB1xp67_ASAP7_75t_L g15777 ( 
.A(n_15678),
.Y(n_15777)
);

INVx1_ASAP7_75t_L g15778 ( 
.A(n_15694),
.Y(n_15778)
);

OAI221xp5_ASAP7_75t_L g15779 ( 
.A1(n_15673),
.A2(n_3576),
.B1(n_3573),
.B2(n_3575),
.C(n_3578),
.Y(n_15779)
);

AOI21xp5_ASAP7_75t_L g15780 ( 
.A1(n_15689),
.A2(n_15688),
.B(n_15674),
.Y(n_15780)
);

INVx2_ASAP7_75t_SL g15781 ( 
.A(n_15700),
.Y(n_15781)
);

INVx1_ASAP7_75t_L g15782 ( 
.A(n_15654),
.Y(n_15782)
);

NAND2xp5_ASAP7_75t_L g15783 ( 
.A(n_15699),
.B(n_3575),
.Y(n_15783)
);

AOI221xp5_ASAP7_75t_L g15784 ( 
.A1(n_15739),
.A2(n_3580),
.B1(n_3578),
.B2(n_3579),
.C(n_3581),
.Y(n_15784)
);

AOI221xp5_ASAP7_75t_L g15785 ( 
.A1(n_15712),
.A2(n_3583),
.B1(n_3580),
.B2(n_3582),
.C(n_3584),
.Y(n_15785)
);

AOI211xp5_ASAP7_75t_L g15786 ( 
.A1(n_15680),
.A2(n_3586),
.B(n_3584),
.C(n_3585),
.Y(n_15786)
);

NAND4xp25_ASAP7_75t_SL g15787 ( 
.A(n_15715),
.B(n_3587),
.C(n_3585),
.D(n_3586),
.Y(n_15787)
);

AOI22xp5_ASAP7_75t_L g15788 ( 
.A1(n_15668),
.A2(n_3590),
.B1(n_3588),
.B2(n_3589),
.Y(n_15788)
);

AND4x1_ASAP7_75t_L g15789 ( 
.A(n_15686),
.B(n_3592),
.C(n_3588),
.D(n_3591),
.Y(n_15789)
);

AOI221xp5_ASAP7_75t_L g15790 ( 
.A1(n_15702),
.A2(n_3594),
.B1(n_3591),
.B2(n_3593),
.C(n_3595),
.Y(n_15790)
);

AOI221xp5_ASAP7_75t_L g15791 ( 
.A1(n_15718),
.A2(n_3596),
.B1(n_3594),
.B2(n_3595),
.C(n_3597),
.Y(n_15791)
);

AOI211xp5_ASAP7_75t_SL g15792 ( 
.A1(n_15707),
.A2(n_3598),
.B(n_3596),
.C(n_3597),
.Y(n_15792)
);

NOR2xp33_ASAP7_75t_R g15793 ( 
.A(n_15672),
.B(n_3598),
.Y(n_15793)
);

CKINVDCx11_ASAP7_75t_R g15794 ( 
.A(n_15721),
.Y(n_15794)
);

NAND2xp5_ASAP7_75t_SL g15795 ( 
.A(n_15670),
.B(n_3599),
.Y(n_15795)
);

BUFx2_ASAP7_75t_L g15796 ( 
.A(n_15741),
.Y(n_15796)
);

OAI211xp5_ASAP7_75t_L g15797 ( 
.A1(n_15684),
.A2(n_3601),
.B(n_3599),
.C(n_3600),
.Y(n_15797)
);

AOI31xp33_ASAP7_75t_L g15798 ( 
.A1(n_15706),
.A2(n_3602),
.A3(n_3600),
.B(n_3601),
.Y(n_15798)
);

OAI211xp5_ASAP7_75t_SL g15799 ( 
.A1(n_15681),
.A2(n_3605),
.B(n_3606),
.C(n_3604),
.Y(n_15799)
);

AOI221xp5_ASAP7_75t_SL g15800 ( 
.A1(n_15708),
.A2(n_3620),
.B1(n_3628),
.B2(n_3611),
.C(n_3603),
.Y(n_15800)
);

AOI211xp5_ASAP7_75t_SL g15801 ( 
.A1(n_15698),
.A2(n_3605),
.B(n_3603),
.C(n_3604),
.Y(n_15801)
);

NOR3xp33_ASAP7_75t_L g15802 ( 
.A(n_15755),
.B(n_3606),
.C(n_3607),
.Y(n_15802)
);

AOI222xp33_ASAP7_75t_L g15803 ( 
.A1(n_15675),
.A2(n_3610),
.B1(n_3612),
.B2(n_3608),
.C1(n_3609),
.C2(n_3611),
.Y(n_15803)
);

AOI211x1_ASAP7_75t_SL g15804 ( 
.A1(n_15690),
.A2(n_3612),
.B(n_3609),
.C(n_3610),
.Y(n_15804)
);

NAND3xp33_ASAP7_75t_L g15805 ( 
.A(n_15756),
.B(n_3613),
.C(n_3614),
.Y(n_15805)
);

OAI211xp5_ASAP7_75t_L g15806 ( 
.A1(n_15757),
.A2(n_3615),
.B(n_3613),
.C(n_3614),
.Y(n_15806)
);

AOI211xp5_ASAP7_75t_L g15807 ( 
.A1(n_15676),
.A2(n_3618),
.B(n_3615),
.C(n_3617),
.Y(n_15807)
);

NAND3xp33_ASAP7_75t_L g15808 ( 
.A(n_15709),
.B(n_3617),
.C(n_3619),
.Y(n_15808)
);

OAI211xp5_ASAP7_75t_L g15809 ( 
.A1(n_15722),
.A2(n_3621),
.B(n_3619),
.C(n_3620),
.Y(n_15809)
);

NOR2xp33_ASAP7_75t_L g15810 ( 
.A(n_15711),
.B(n_3621),
.Y(n_15810)
);

AND2x2_ASAP7_75t_L g15811 ( 
.A(n_15729),
.B(n_3622),
.Y(n_15811)
);

NAND2xp5_ASAP7_75t_L g15812 ( 
.A(n_15746),
.B(n_3622),
.Y(n_15812)
);

NOR2x1_ASAP7_75t_L g15813 ( 
.A(n_15669),
.B(n_3623),
.Y(n_15813)
);

AOI221xp5_ASAP7_75t_L g15814 ( 
.A1(n_15679),
.A2(n_3625),
.B1(n_3623),
.B2(n_3624),
.C(n_3626),
.Y(n_15814)
);

INVx1_ASAP7_75t_SL g15815 ( 
.A(n_15655),
.Y(n_15815)
);

NAND4xp25_ASAP7_75t_L g15816 ( 
.A(n_15697),
.B(n_3633),
.C(n_3641),
.D(n_3624),
.Y(n_15816)
);

OAI211xp5_ASAP7_75t_SL g15817 ( 
.A1(n_15717),
.A2(n_15683),
.B(n_15704),
.C(n_15703),
.Y(n_15817)
);

OAI211xp5_ASAP7_75t_L g15818 ( 
.A1(n_15658),
.A2(n_3628),
.B(n_3625),
.C(n_3627),
.Y(n_15818)
);

AOI22xp5_ASAP7_75t_L g15819 ( 
.A1(n_15716),
.A2(n_15657),
.B1(n_15732),
.B2(n_15723),
.Y(n_15819)
);

NOR2xp33_ASAP7_75t_R g15820 ( 
.A(n_15730),
.B(n_3629),
.Y(n_15820)
);

AOI22x1_ASAP7_75t_L g15821 ( 
.A1(n_15738),
.A2(n_15656),
.B1(n_15685),
.B2(n_15693),
.Y(n_15821)
);

AOI221xp5_ASAP7_75t_L g15822 ( 
.A1(n_15701),
.A2(n_3631),
.B1(n_3629),
.B2(n_3630),
.C(n_3632),
.Y(n_15822)
);

AOI21xp5_ASAP7_75t_L g15823 ( 
.A1(n_15747),
.A2(n_3630),
.B(n_3631),
.Y(n_15823)
);

NOR3xp33_ASAP7_75t_L g15824 ( 
.A(n_15691),
.B(n_3632),
.C(n_3634),
.Y(n_15824)
);

O2A1O1Ixp33_ASAP7_75t_L g15825 ( 
.A1(n_15682),
.A2(n_3636),
.B(n_3634),
.C(n_3635),
.Y(n_15825)
);

OAI211xp5_ASAP7_75t_SL g15826 ( 
.A1(n_15719),
.A2(n_3638),
.B(n_3639),
.C(n_3637),
.Y(n_15826)
);

OAI311xp33_ASAP7_75t_L g15827 ( 
.A1(n_15705),
.A2(n_3638),
.A3(n_3635),
.B1(n_3637),
.C1(n_3639),
.Y(n_15827)
);

AOI21xp33_ASAP7_75t_L g15828 ( 
.A1(n_15666),
.A2(n_4104),
.B(n_4103),
.Y(n_15828)
);

INVx1_ASAP7_75t_L g15829 ( 
.A(n_15733),
.Y(n_15829)
);

INVx2_ASAP7_75t_L g15830 ( 
.A(n_15696),
.Y(n_15830)
);

INVxp67_ASAP7_75t_SL g15831 ( 
.A(n_15742),
.Y(n_15831)
);

OAI211xp5_ASAP7_75t_L g15832 ( 
.A1(n_15737),
.A2(n_3642),
.B(n_3640),
.C(n_3641),
.Y(n_15832)
);

NOR3xp33_ASAP7_75t_SL g15833 ( 
.A(n_15725),
.B(n_3642),
.C(n_3643),
.Y(n_15833)
);

AOI22xp5_ASAP7_75t_L g15834 ( 
.A1(n_15734),
.A2(n_3645),
.B1(n_3643),
.B2(n_3644),
.Y(n_15834)
);

AOI322xp5_ASAP7_75t_L g15835 ( 
.A1(n_15714),
.A2(n_3650),
.A3(n_3649),
.B1(n_3647),
.B2(n_3644),
.C1(n_3646),
.C2(n_3648),
.Y(n_15835)
);

OAI221xp5_ASAP7_75t_SL g15836 ( 
.A1(n_15735),
.A2(n_3651),
.B1(n_3647),
.B2(n_3649),
.C(n_3652),
.Y(n_15836)
);

NOR2x1_ASAP7_75t_L g15837 ( 
.A(n_15763),
.B(n_15731),
.Y(n_15837)
);

INVx1_ASAP7_75t_L g15838 ( 
.A(n_15759),
.Y(n_15838)
);

INVx1_ASAP7_75t_L g15839 ( 
.A(n_15759),
.Y(n_15839)
);

NOR2x1_ASAP7_75t_L g15840 ( 
.A(n_15778),
.B(n_15744),
.Y(n_15840)
);

NOR3xp33_ASAP7_75t_L g15841 ( 
.A(n_15762),
.B(n_15758),
.C(n_15748),
.Y(n_15841)
);

NOR3xp33_ASAP7_75t_L g15842 ( 
.A(n_15781),
.B(n_15660),
.C(n_15754),
.Y(n_15842)
);

INVx1_ASAP7_75t_L g15843 ( 
.A(n_15759),
.Y(n_15843)
);

AND2x2_ASAP7_75t_L g15844 ( 
.A(n_15796),
.B(n_15736),
.Y(n_15844)
);

INVx1_ASAP7_75t_L g15845 ( 
.A(n_15777),
.Y(n_15845)
);

NOR3x2_ASAP7_75t_L g15846 ( 
.A(n_15794),
.B(n_15817),
.C(n_15775),
.Y(n_15846)
);

NAND3xp33_ASAP7_75t_L g15847 ( 
.A(n_15782),
.B(n_15665),
.C(n_15745),
.Y(n_15847)
);

NOR3xp33_ASAP7_75t_L g15848 ( 
.A(n_15769),
.B(n_15750),
.C(n_15749),
.Y(n_15848)
);

NOR2x1_ASAP7_75t_L g15849 ( 
.A(n_15829),
.B(n_15740),
.Y(n_15849)
);

INVx3_ASAP7_75t_SL g15850 ( 
.A(n_15815),
.Y(n_15850)
);

NOR2xp67_ASAP7_75t_L g15851 ( 
.A(n_15780),
.B(n_15743),
.Y(n_15851)
);

NOR2xp33_ASAP7_75t_L g15852 ( 
.A(n_15831),
.B(n_15752),
.Y(n_15852)
);

NOR2x1p5_ASAP7_75t_L g15853 ( 
.A(n_15812),
.B(n_15727),
.Y(n_15853)
);

NOR3xp33_ASAP7_75t_L g15854 ( 
.A(n_15770),
.B(n_3651),
.C(n_3652),
.Y(n_15854)
);

INVx1_ASAP7_75t_SL g15855 ( 
.A(n_15793),
.Y(n_15855)
);

AND3x4_ASAP7_75t_L g15856 ( 
.A(n_15802),
.B(n_3661),
.C(n_3653),
.Y(n_15856)
);

NOR4xp25_ASAP7_75t_L g15857 ( 
.A(n_15830),
.B(n_3655),
.C(n_3653),
.D(n_3654),
.Y(n_15857)
);

NAND2x2_ASAP7_75t_L g15858 ( 
.A(n_15783),
.B(n_4102),
.Y(n_15858)
);

NOR3x2_ASAP7_75t_L g15859 ( 
.A(n_15810),
.B(n_3655),
.C(n_3656),
.Y(n_15859)
);

NOR3xp33_ASAP7_75t_L g15860 ( 
.A(n_15795),
.B(n_3656),
.C(n_3657),
.Y(n_15860)
);

NOR3xp33_ASAP7_75t_L g15861 ( 
.A(n_15799),
.B(n_3657),
.C(n_3658),
.Y(n_15861)
);

NOR3xp33_ASAP7_75t_L g15862 ( 
.A(n_15772),
.B(n_3658),
.C(n_3659),
.Y(n_15862)
);

OR2x2_ASAP7_75t_L g15863 ( 
.A(n_15761),
.B(n_3659),
.Y(n_15863)
);

AOI21x1_ASAP7_75t_L g15864 ( 
.A1(n_15811),
.A2(n_3660),
.B(n_3661),
.Y(n_15864)
);

NAND4xp75_ASAP7_75t_L g15865 ( 
.A(n_15813),
.B(n_3663),
.C(n_3660),
.D(n_3662),
.Y(n_15865)
);

INVx1_ASAP7_75t_L g15866 ( 
.A(n_15821),
.Y(n_15866)
);

INVx1_ASAP7_75t_L g15867 ( 
.A(n_15805),
.Y(n_15867)
);

AND2x2_ASAP7_75t_L g15868 ( 
.A(n_15792),
.B(n_15833),
.Y(n_15868)
);

NOR3xp33_ASAP7_75t_L g15869 ( 
.A(n_15806),
.B(n_3662),
.C(n_3663),
.Y(n_15869)
);

INVx1_ASAP7_75t_L g15870 ( 
.A(n_15819),
.Y(n_15870)
);

NOR2x1_ASAP7_75t_L g15871 ( 
.A(n_15816),
.B(n_3664),
.Y(n_15871)
);

AND2x2_ASAP7_75t_L g15872 ( 
.A(n_15801),
.B(n_3664),
.Y(n_15872)
);

NAND3xp33_ASAP7_75t_L g15873 ( 
.A(n_15785),
.B(n_3665),
.C(n_3666),
.Y(n_15873)
);

NAND2xp5_ASAP7_75t_L g15874 ( 
.A(n_15804),
.B(n_3665),
.Y(n_15874)
);

NAND4xp75_ASAP7_75t_L g15875 ( 
.A(n_15800),
.B(n_3669),
.C(n_3667),
.D(n_3668),
.Y(n_15875)
);

NAND3xp33_ASAP7_75t_SL g15876 ( 
.A(n_15820),
.B(n_3667),
.C(n_3668),
.Y(n_15876)
);

NAND2xp5_ASAP7_75t_L g15877 ( 
.A(n_15807),
.B(n_3669),
.Y(n_15877)
);

XOR2x1_ASAP7_75t_L g15878 ( 
.A(n_15773),
.B(n_3670),
.Y(n_15878)
);

NOR3xp33_ASAP7_75t_L g15879 ( 
.A(n_15809),
.B(n_3670),
.C(n_3671),
.Y(n_15879)
);

NAND2xp5_ASAP7_75t_L g15880 ( 
.A(n_15789),
.B(n_3671),
.Y(n_15880)
);

NOR2xp33_ASAP7_75t_L g15881 ( 
.A(n_15779),
.B(n_3672),
.Y(n_15881)
);

NOR2x1_ASAP7_75t_L g15882 ( 
.A(n_15808),
.B(n_3672),
.Y(n_15882)
);

OAI21xp33_ASAP7_75t_L g15883 ( 
.A1(n_15774),
.A2(n_3673),
.B(n_3674),
.Y(n_15883)
);

NAND2xp5_ASAP7_75t_SL g15884 ( 
.A(n_15766),
.B(n_3673),
.Y(n_15884)
);

AND3x4_ASAP7_75t_L g15885 ( 
.A(n_15824),
.B(n_3682),
.C(n_3674),
.Y(n_15885)
);

NOR2x1_ASAP7_75t_L g15886 ( 
.A(n_15797),
.B(n_3675),
.Y(n_15886)
);

INVx1_ASAP7_75t_L g15887 ( 
.A(n_15776),
.Y(n_15887)
);

OR2x2_ASAP7_75t_L g15888 ( 
.A(n_15798),
.B(n_15787),
.Y(n_15888)
);

NOR2x1_ASAP7_75t_L g15889 ( 
.A(n_15818),
.B(n_3675),
.Y(n_15889)
);

NOR2x1p5_ASAP7_75t_L g15890 ( 
.A(n_15827),
.B(n_4120),
.Y(n_15890)
);

NOR2x1_ASAP7_75t_L g15891 ( 
.A(n_15826),
.B(n_15832),
.Y(n_15891)
);

AND3x1_ASAP7_75t_L g15892 ( 
.A(n_15784),
.B(n_3676),
.C(n_3677),
.Y(n_15892)
);

NOR2x1_ASAP7_75t_L g15893 ( 
.A(n_15760),
.B(n_3677),
.Y(n_15893)
);

NAND2xp5_ASAP7_75t_L g15894 ( 
.A(n_15823),
.B(n_3678),
.Y(n_15894)
);

NOR2x1_ASAP7_75t_L g15895 ( 
.A(n_15825),
.B(n_3678),
.Y(n_15895)
);

INVx1_ASAP7_75t_L g15896 ( 
.A(n_15834),
.Y(n_15896)
);

INVxp67_ASAP7_75t_L g15897 ( 
.A(n_15803),
.Y(n_15897)
);

NOR2x1_ASAP7_75t_L g15898 ( 
.A(n_15828),
.B(n_3679),
.Y(n_15898)
);

INVx1_ASAP7_75t_L g15899 ( 
.A(n_15788),
.Y(n_15899)
);

INVx1_ASAP7_75t_L g15900 ( 
.A(n_15845),
.Y(n_15900)
);

INVx1_ASAP7_75t_L g15901 ( 
.A(n_15846),
.Y(n_15901)
);

INVx1_ASAP7_75t_L g15902 ( 
.A(n_15838),
.Y(n_15902)
);

XNOR2xp5_ASAP7_75t_SL g15903 ( 
.A(n_15839),
.B(n_15790),
.Y(n_15903)
);

INVx1_ASAP7_75t_L g15904 ( 
.A(n_15843),
.Y(n_15904)
);

AOI22xp5_ASAP7_75t_L g15905 ( 
.A1(n_15850),
.A2(n_15866),
.B1(n_15856),
.B2(n_15870),
.Y(n_15905)
);

NAND2xp5_ASAP7_75t_L g15906 ( 
.A(n_15855),
.B(n_15814),
.Y(n_15906)
);

INVx1_ASAP7_75t_L g15907 ( 
.A(n_15837),
.Y(n_15907)
);

OR2x2_ASAP7_75t_L g15908 ( 
.A(n_15887),
.B(n_15888),
.Y(n_15908)
);

AOI22xp5_ASAP7_75t_L g15909 ( 
.A1(n_15890),
.A2(n_15791),
.B1(n_15822),
.B2(n_15786),
.Y(n_15909)
);

INVx1_ASAP7_75t_L g15910 ( 
.A(n_15840),
.Y(n_15910)
);

NOR3xp33_ASAP7_75t_L g15911 ( 
.A(n_15852),
.B(n_15836),
.C(n_15768),
.Y(n_15911)
);

HB1xp67_ASAP7_75t_L g15912 ( 
.A(n_15851),
.Y(n_15912)
);

INVx2_ASAP7_75t_L g15913 ( 
.A(n_15868),
.Y(n_15913)
);

XNOR2xp5_ASAP7_75t_L g15914 ( 
.A(n_15853),
.B(n_15771),
.Y(n_15914)
);

BUFx3_ASAP7_75t_L g15915 ( 
.A(n_15844),
.Y(n_15915)
);

NOR3xp33_ASAP7_75t_L g15916 ( 
.A(n_15849),
.B(n_15765),
.C(n_15764),
.Y(n_15916)
);

NAND4xp75_ASAP7_75t_L g15917 ( 
.A(n_15898),
.B(n_15767),
.C(n_15835),
.D(n_3682),
.Y(n_15917)
);

OAI221xp5_ASAP7_75t_L g15918 ( 
.A1(n_15858),
.A2(n_15874),
.B1(n_15863),
.B2(n_15854),
.C(n_15857),
.Y(n_15918)
);

NOR2x1_ASAP7_75t_L g15919 ( 
.A(n_15847),
.B(n_3680),
.Y(n_15919)
);

NAND2xp5_ASAP7_75t_L g15920 ( 
.A(n_15842),
.B(n_4096),
.Y(n_15920)
);

INVx2_ASAP7_75t_L g15921 ( 
.A(n_15864),
.Y(n_15921)
);

NOR2xp33_ASAP7_75t_L g15922 ( 
.A(n_15897),
.B(n_15876),
.Y(n_15922)
);

NOR2x1_ASAP7_75t_L g15923 ( 
.A(n_15867),
.B(n_3680),
.Y(n_15923)
);

NAND2xp5_ASAP7_75t_L g15924 ( 
.A(n_15841),
.B(n_4097),
.Y(n_15924)
);

INVx1_ASAP7_75t_L g15925 ( 
.A(n_15872),
.Y(n_15925)
);

INVx2_ASAP7_75t_L g15926 ( 
.A(n_15859),
.Y(n_15926)
);

XOR2xp5_ASAP7_75t_L g15927 ( 
.A(n_15878),
.B(n_3681),
.Y(n_15927)
);

OR2x2_ASAP7_75t_L g15928 ( 
.A(n_15880),
.B(n_3681),
.Y(n_15928)
);

INVx2_ASAP7_75t_L g15929 ( 
.A(n_15891),
.Y(n_15929)
);

XNOR2x1_ASAP7_75t_L g15930 ( 
.A(n_15885),
.B(n_3684),
.Y(n_15930)
);

HB1xp67_ASAP7_75t_L g15931 ( 
.A(n_15848),
.Y(n_15931)
);

INVx1_ASAP7_75t_L g15932 ( 
.A(n_15871),
.Y(n_15932)
);

AO22x2_ASAP7_75t_L g15933 ( 
.A1(n_15899),
.A2(n_3686),
.B1(n_3684),
.B2(n_3685),
.Y(n_15933)
);

AND2x2_ASAP7_75t_L g15934 ( 
.A(n_15886),
.B(n_3685),
.Y(n_15934)
);

NOR2x1_ASAP7_75t_L g15935 ( 
.A(n_15865),
.B(n_3686),
.Y(n_15935)
);

AOI22xp5_ASAP7_75t_L g15936 ( 
.A1(n_15862),
.A2(n_3689),
.B1(n_3687),
.B2(n_3688),
.Y(n_15936)
);

OAI21xp5_ASAP7_75t_L g15937 ( 
.A1(n_15889),
.A2(n_15882),
.B(n_15877),
.Y(n_15937)
);

NOR2x1_ASAP7_75t_L g15938 ( 
.A(n_15896),
.B(n_3687),
.Y(n_15938)
);

INVx1_ASAP7_75t_L g15939 ( 
.A(n_15893),
.Y(n_15939)
);

INVx1_ASAP7_75t_L g15940 ( 
.A(n_15894),
.Y(n_15940)
);

AND2x2_ASAP7_75t_L g15941 ( 
.A(n_15895),
.B(n_3689),
.Y(n_15941)
);

AOI22xp33_ASAP7_75t_SL g15942 ( 
.A1(n_15881),
.A2(n_3692),
.B1(n_3690),
.B2(n_3691),
.Y(n_15942)
);

INVx2_ASAP7_75t_SL g15943 ( 
.A(n_15884),
.Y(n_15943)
);

XOR2xp5_ASAP7_75t_L g15944 ( 
.A(n_15875),
.B(n_3690),
.Y(n_15944)
);

INVxp67_ASAP7_75t_L g15945 ( 
.A(n_15892),
.Y(n_15945)
);

AOI211xp5_ASAP7_75t_L g15946 ( 
.A1(n_15860),
.A2(n_3694),
.B(n_3691),
.C(n_3693),
.Y(n_15946)
);

NAND4xp75_ASAP7_75t_L g15947 ( 
.A(n_15879),
.B(n_3695),
.C(n_3693),
.D(n_3694),
.Y(n_15947)
);

INVxp33_ASAP7_75t_SL g15948 ( 
.A(n_15861),
.Y(n_15948)
);

XNOR2xp5_ASAP7_75t_L g15949 ( 
.A(n_15873),
.B(n_3696),
.Y(n_15949)
);

HB1xp67_ASAP7_75t_L g15950 ( 
.A(n_15869),
.Y(n_15950)
);

XNOR2x1_ASAP7_75t_L g15951 ( 
.A(n_15883),
.B(n_3695),
.Y(n_15951)
);

AOI22xp5_ASAP7_75t_L g15952 ( 
.A1(n_15845),
.A2(n_3698),
.B1(n_3696),
.B2(n_3697),
.Y(n_15952)
);

NAND2xp5_ASAP7_75t_L g15953 ( 
.A(n_15845),
.B(n_4096),
.Y(n_15953)
);

INVx1_ASAP7_75t_L g15954 ( 
.A(n_15845),
.Y(n_15954)
);

INVxp33_ASAP7_75t_L g15955 ( 
.A(n_15845),
.Y(n_15955)
);

AND2x4_ASAP7_75t_L g15956 ( 
.A(n_15845),
.B(n_3698),
.Y(n_15956)
);

AND2x2_ASAP7_75t_L g15957 ( 
.A(n_15955),
.B(n_3699),
.Y(n_15957)
);

NAND4xp75_ASAP7_75t_L g15958 ( 
.A(n_15910),
.B(n_3703),
.C(n_3701),
.D(n_3702),
.Y(n_15958)
);

INVx1_ASAP7_75t_L g15959 ( 
.A(n_15907),
.Y(n_15959)
);

XOR2xp5_ASAP7_75t_L g15960 ( 
.A(n_15931),
.B(n_3701),
.Y(n_15960)
);

NAND2xp5_ASAP7_75t_L g15961 ( 
.A(n_15900),
.B(n_3702),
.Y(n_15961)
);

NAND3xp33_ASAP7_75t_L g15962 ( 
.A(n_15954),
.B(n_3703),
.C(n_3704),
.Y(n_15962)
);

AND3x1_ASAP7_75t_L g15963 ( 
.A(n_15921),
.B(n_3704),
.C(n_3705),
.Y(n_15963)
);

INVx1_ASAP7_75t_L g15964 ( 
.A(n_15912),
.Y(n_15964)
);

INVx1_ASAP7_75t_L g15965 ( 
.A(n_15915),
.Y(n_15965)
);

AND2x4_ASAP7_75t_L g15966 ( 
.A(n_15901),
.B(n_3705),
.Y(n_15966)
);

INVx1_ASAP7_75t_L g15967 ( 
.A(n_15929),
.Y(n_15967)
);

NOR2x1_ASAP7_75t_L g15968 ( 
.A(n_15908),
.B(n_3706),
.Y(n_15968)
);

XOR2x1_ASAP7_75t_L g15969 ( 
.A(n_15902),
.B(n_15904),
.Y(n_15969)
);

NAND2xp5_ASAP7_75t_L g15970 ( 
.A(n_15905),
.B(n_3706),
.Y(n_15970)
);

INVx3_ASAP7_75t_L g15971 ( 
.A(n_15913),
.Y(n_15971)
);

INVx2_ASAP7_75t_L g15972 ( 
.A(n_15939),
.Y(n_15972)
);

NAND2xp5_ASAP7_75t_SL g15973 ( 
.A(n_15932),
.B(n_3707),
.Y(n_15973)
);

INVx2_ASAP7_75t_L g15974 ( 
.A(n_15930),
.Y(n_15974)
);

NAND2xp5_ASAP7_75t_L g15975 ( 
.A(n_15925),
.B(n_3707),
.Y(n_15975)
);

XNOR2x1_ASAP7_75t_L g15976 ( 
.A(n_15914),
.B(n_3709),
.Y(n_15976)
);

INVx2_ASAP7_75t_L g15977 ( 
.A(n_15926),
.Y(n_15977)
);

INVx1_ASAP7_75t_L g15978 ( 
.A(n_15927),
.Y(n_15978)
);

INVx2_ASAP7_75t_SL g15979 ( 
.A(n_15940),
.Y(n_15979)
);

XNOR2xp5_ASAP7_75t_L g15980 ( 
.A(n_15918),
.B(n_3709),
.Y(n_15980)
);

NOR2x1_ASAP7_75t_L g15981 ( 
.A(n_15922),
.B(n_3710),
.Y(n_15981)
);

XOR2xp5_ASAP7_75t_L g15982 ( 
.A(n_15903),
.B(n_3711),
.Y(n_15982)
);

NOR2xp67_ASAP7_75t_L g15983 ( 
.A(n_15945),
.B(n_3712),
.Y(n_15983)
);

XNOR2xp5_ASAP7_75t_L g15984 ( 
.A(n_15948),
.B(n_3711),
.Y(n_15984)
);

XNOR2xp5_ASAP7_75t_L g15985 ( 
.A(n_15944),
.B(n_3713),
.Y(n_15985)
);

NAND2xp5_ASAP7_75t_L g15986 ( 
.A(n_15937),
.B(n_3713),
.Y(n_15986)
);

INVx1_ASAP7_75t_L g15987 ( 
.A(n_15934),
.Y(n_15987)
);

INVx1_ASAP7_75t_L g15988 ( 
.A(n_15941),
.Y(n_15988)
);

NOR2x1_ASAP7_75t_L g15989 ( 
.A(n_15906),
.B(n_3714),
.Y(n_15989)
);

INVx2_ASAP7_75t_L g15990 ( 
.A(n_15928),
.Y(n_15990)
);

AND2x2_ASAP7_75t_L g15991 ( 
.A(n_15950),
.B(n_3714),
.Y(n_15991)
);

AND2x2_ASAP7_75t_L g15992 ( 
.A(n_15938),
.B(n_3715),
.Y(n_15992)
);

INVx2_ASAP7_75t_L g15993 ( 
.A(n_15943),
.Y(n_15993)
);

NAND2xp5_ASAP7_75t_L g15994 ( 
.A(n_15911),
.B(n_3715),
.Y(n_15994)
);

INVx1_ASAP7_75t_L g15995 ( 
.A(n_15923),
.Y(n_15995)
);

INVx2_ASAP7_75t_SL g15996 ( 
.A(n_15919),
.Y(n_15996)
);

OAI22xp5_ASAP7_75t_L g15997 ( 
.A1(n_15936),
.A2(n_3718),
.B1(n_3716),
.B2(n_3717),
.Y(n_15997)
);

INVx1_ASAP7_75t_L g15998 ( 
.A(n_15924),
.Y(n_15998)
);

NAND3xp33_ASAP7_75t_L g15999 ( 
.A(n_15916),
.B(n_3717),
.C(n_3719),
.Y(n_15999)
);

INVx1_ASAP7_75t_L g16000 ( 
.A(n_15920),
.Y(n_16000)
);

XNOR2xp5_ASAP7_75t_L g16001 ( 
.A(n_15909),
.B(n_3719),
.Y(n_16001)
);

NAND2xp5_ASAP7_75t_L g16002 ( 
.A(n_15935),
.B(n_3720),
.Y(n_16002)
);

NOR4xp75_ASAP7_75t_L g16003 ( 
.A(n_15917),
.B(n_3722),
.C(n_3720),
.D(n_3721),
.Y(n_16003)
);

NOR2x1_ASAP7_75t_L g16004 ( 
.A(n_15947),
.B(n_3721),
.Y(n_16004)
);

AOI22xp5_ASAP7_75t_L g16005 ( 
.A1(n_15942),
.A2(n_15949),
.B1(n_15951),
.B2(n_15946),
.Y(n_16005)
);

NAND4xp75_ASAP7_75t_L g16006 ( 
.A(n_15953),
.B(n_3725),
.C(n_3723),
.D(n_3724),
.Y(n_16006)
);

AND2x4_ASAP7_75t_L g16007 ( 
.A(n_15956),
.B(n_3723),
.Y(n_16007)
);

NAND4xp75_ASAP7_75t_L g16008 ( 
.A(n_15952),
.B(n_3727),
.C(n_3725),
.D(n_3726),
.Y(n_16008)
);

XNOR2x1_ASAP7_75t_L g16009 ( 
.A(n_15933),
.B(n_3727),
.Y(n_16009)
);

INVx1_ASAP7_75t_L g16010 ( 
.A(n_15956),
.Y(n_16010)
);

NOR2xp67_ASAP7_75t_L g16011 ( 
.A(n_15933),
.B(n_3729),
.Y(n_16011)
);

INVx1_ASAP7_75t_L g16012 ( 
.A(n_15910),
.Y(n_16012)
);

INVx1_ASAP7_75t_L g16013 ( 
.A(n_15910),
.Y(n_16013)
);

AND2x4_ASAP7_75t_L g16014 ( 
.A(n_15910),
.B(n_3728),
.Y(n_16014)
);

HB1xp67_ASAP7_75t_L g16015 ( 
.A(n_15910),
.Y(n_16015)
);

XNOR2xp5_ASAP7_75t_L g16016 ( 
.A(n_15955),
.B(n_3728),
.Y(n_16016)
);

INVx2_ASAP7_75t_L g16017 ( 
.A(n_15921),
.Y(n_16017)
);

NOR3xp33_ASAP7_75t_L g16018 ( 
.A(n_15971),
.B(n_16015),
.C(n_15964),
.Y(n_16018)
);

XNOR2xp5_ASAP7_75t_L g16019 ( 
.A(n_15969),
.B(n_3729),
.Y(n_16019)
);

NAND2xp5_ASAP7_75t_L g16020 ( 
.A(n_15965),
.B(n_15959),
.Y(n_16020)
);

NAND3x1_ASAP7_75t_L g16021 ( 
.A(n_16012),
.B(n_16013),
.C(n_15967),
.Y(n_16021)
);

NOR3xp33_ASAP7_75t_L g16022 ( 
.A(n_15979),
.B(n_3730),
.C(n_3731),
.Y(n_16022)
);

INVx1_ASAP7_75t_L g16023 ( 
.A(n_16017),
.Y(n_16023)
);

NOR3xp33_ASAP7_75t_SL g16024 ( 
.A(n_15987),
.B(n_3731),
.C(n_3732),
.Y(n_16024)
);

AND2x2_ASAP7_75t_L g16025 ( 
.A(n_15972),
.B(n_3733),
.Y(n_16025)
);

AOI21xp33_ASAP7_75t_SL g16026 ( 
.A1(n_15993),
.A2(n_3734),
.B(n_3735),
.Y(n_16026)
);

NAND2xp5_ASAP7_75t_L g16027 ( 
.A(n_15988),
.B(n_3734),
.Y(n_16027)
);

INVx1_ASAP7_75t_L g16028 ( 
.A(n_15995),
.Y(n_16028)
);

OAI211xp5_ASAP7_75t_L g16029 ( 
.A1(n_15977),
.A2(n_3737),
.B(n_3735),
.C(n_3736),
.Y(n_16029)
);

NOR2x1_ASAP7_75t_L g16030 ( 
.A(n_16010),
.B(n_3737),
.Y(n_16030)
);

XOR2xp5_ASAP7_75t_L g16031 ( 
.A(n_15978),
.B(n_15990),
.Y(n_16031)
);

NOR2xp33_ASAP7_75t_L g16032 ( 
.A(n_15996),
.B(n_3738),
.Y(n_16032)
);

NAND4xp25_ASAP7_75t_SL g16033 ( 
.A(n_15968),
.B(n_3747),
.C(n_3755),
.D(n_3739),
.Y(n_16033)
);

NAND2x1_ASAP7_75t_L g16034 ( 
.A(n_15992),
.B(n_3739),
.Y(n_16034)
);

NOR2x1p5_ASAP7_75t_L g16035 ( 
.A(n_15974),
.B(n_3740),
.Y(n_16035)
);

AOI221xp5_ASAP7_75t_L g16036 ( 
.A1(n_15963),
.A2(n_16002),
.B1(n_15980),
.B2(n_15998),
.C(n_16000),
.Y(n_16036)
);

INVx1_ASAP7_75t_L g16037 ( 
.A(n_16009),
.Y(n_16037)
);

INVx1_ASAP7_75t_L g16038 ( 
.A(n_16011),
.Y(n_16038)
);

AO22x2_ASAP7_75t_L g16039 ( 
.A1(n_15982),
.A2(n_3742),
.B1(n_3740),
.B2(n_3741),
.Y(n_16039)
);

NAND3xp33_ASAP7_75t_SL g16040 ( 
.A(n_16005),
.B(n_3741),
.C(n_3742),
.Y(n_16040)
);

AND5x1_ASAP7_75t_L g16041 ( 
.A(n_15985),
.B(n_3745),
.C(n_3743),
.D(n_3744),
.E(n_3746),
.Y(n_16041)
);

AOI21xp5_ASAP7_75t_L g16042 ( 
.A1(n_15994),
.A2(n_3744),
.B(n_3746),
.Y(n_16042)
);

NAND3xp33_ASAP7_75t_SL g16043 ( 
.A(n_16003),
.B(n_15970),
.C(n_15986),
.Y(n_16043)
);

OR2x2_ASAP7_75t_L g16044 ( 
.A(n_16007),
.B(n_3747),
.Y(n_16044)
);

AOI21xp5_ASAP7_75t_L g16045 ( 
.A1(n_15989),
.A2(n_3748),
.B(n_3749),
.Y(n_16045)
);

AOI22xp5_ASAP7_75t_L g16046 ( 
.A1(n_15983),
.A2(n_15981),
.B1(n_15991),
.B2(n_15976),
.Y(n_16046)
);

NAND3xp33_ASAP7_75t_SL g16047 ( 
.A(n_15973),
.B(n_3749),
.C(n_3750),
.Y(n_16047)
);

AND2x2_ASAP7_75t_L g16048 ( 
.A(n_15957),
.B(n_3750),
.Y(n_16048)
);

NOR2xp67_ASAP7_75t_L g16049 ( 
.A(n_15975),
.B(n_3751),
.Y(n_16049)
);

INVx1_ASAP7_75t_L g16050 ( 
.A(n_16001),
.Y(n_16050)
);

A2O1A1Ixp33_ASAP7_75t_L g16051 ( 
.A1(n_16004),
.A2(n_3754),
.B(n_3752),
.C(n_3753),
.Y(n_16051)
);

HB1xp67_ASAP7_75t_L g16052 ( 
.A(n_15966),
.Y(n_16052)
);

HB1xp67_ASAP7_75t_L g16053 ( 
.A(n_15960),
.Y(n_16053)
);

NOR4xp75_ASAP7_75t_L g16054 ( 
.A(n_16008),
.B(n_3754),
.C(n_3752),
.D(n_3753),
.Y(n_16054)
);

AO22x2_ASAP7_75t_L g16055 ( 
.A1(n_16006),
.A2(n_3758),
.B1(n_3755),
.B2(n_3756),
.Y(n_16055)
);

AOI22xp5_ASAP7_75t_L g16056 ( 
.A1(n_16016),
.A2(n_3759),
.B1(n_3756),
.B2(n_3758),
.Y(n_16056)
);

INVx1_ASAP7_75t_L g16057 ( 
.A(n_15984),
.Y(n_16057)
);

NOR3xp33_ASAP7_75t_L g16058 ( 
.A(n_15999),
.B(n_3760),
.C(n_3761),
.Y(n_16058)
);

INVx1_ASAP7_75t_L g16059 ( 
.A(n_15961),
.Y(n_16059)
);

AOI221xp5_ASAP7_75t_SL g16060 ( 
.A1(n_15997),
.A2(n_3762),
.B1(n_3760),
.B2(n_3761),
.C(n_3763),
.Y(n_16060)
);

NOR3xp33_ASAP7_75t_L g16061 ( 
.A(n_15962),
.B(n_3762),
.C(n_3763),
.Y(n_16061)
);

INVx3_ASAP7_75t_L g16062 ( 
.A(n_16014),
.Y(n_16062)
);

AOI21xp5_ASAP7_75t_L g16063 ( 
.A1(n_15958),
.A2(n_3764),
.B(n_3765),
.Y(n_16063)
);

AND2x4_ASAP7_75t_L g16064 ( 
.A(n_15971),
.B(n_3765),
.Y(n_16064)
);

AOI211xp5_ASAP7_75t_L g16065 ( 
.A1(n_16015),
.A2(n_3767),
.B(n_3764),
.C(n_3766),
.Y(n_16065)
);

AND2x4_ASAP7_75t_L g16066 ( 
.A(n_15971),
.B(n_3767),
.Y(n_16066)
);

INVx1_ASAP7_75t_L g16067 ( 
.A(n_16015),
.Y(n_16067)
);

AOI221xp5_ASAP7_75t_L g16068 ( 
.A1(n_16015),
.A2(n_3770),
.B1(n_3766),
.B2(n_3768),
.C(n_3771),
.Y(n_16068)
);

AOI22xp5_ASAP7_75t_L g16069 ( 
.A1(n_16015),
.A2(n_3771),
.B1(n_3768),
.B2(n_3770),
.Y(n_16069)
);

OAI22xp5_ASAP7_75t_L g16070 ( 
.A1(n_16015),
.A2(n_3774),
.B1(n_3772),
.B2(n_3773),
.Y(n_16070)
);

HB1xp67_ASAP7_75t_L g16071 ( 
.A(n_16015),
.Y(n_16071)
);

AOI31xp33_ASAP7_75t_L g16072 ( 
.A1(n_16015),
.A2(n_3774),
.A3(n_3772),
.B(n_3773),
.Y(n_16072)
);

AOI22xp5_ASAP7_75t_L g16073 ( 
.A1(n_16015),
.A2(n_3777),
.B1(n_3775),
.B2(n_3776),
.Y(n_16073)
);

AND2x4_ASAP7_75t_L g16074 ( 
.A(n_15971),
.B(n_3776),
.Y(n_16074)
);

AO22x2_ASAP7_75t_L g16075 ( 
.A1(n_15965),
.A2(n_3778),
.B1(n_3775),
.B2(n_3777),
.Y(n_16075)
);

AOI22xp5_ASAP7_75t_L g16076 ( 
.A1(n_16015),
.A2(n_3780),
.B1(n_3778),
.B2(n_3779),
.Y(n_16076)
);

CKINVDCx20_ASAP7_75t_R g16077 ( 
.A(n_16015),
.Y(n_16077)
);

NOR2x2_ASAP7_75t_L g16078 ( 
.A(n_16017),
.B(n_3780),
.Y(n_16078)
);

NAND2xp5_ASAP7_75t_L g16079 ( 
.A(n_16015),
.B(n_3781),
.Y(n_16079)
);

OAI211xp5_ASAP7_75t_SL g16080 ( 
.A1(n_15964),
.A2(n_3783),
.B(n_3781),
.C(n_3782),
.Y(n_16080)
);

AND2x4_ASAP7_75t_L g16081 ( 
.A(n_15971),
.B(n_3783),
.Y(n_16081)
);

NOR2xp67_ASAP7_75t_L g16082 ( 
.A(n_16015),
.B(n_3782),
.Y(n_16082)
);

INVx1_ASAP7_75t_L g16083 ( 
.A(n_16015),
.Y(n_16083)
);

NAND4xp25_ASAP7_75t_L g16084 ( 
.A(n_15964),
.B(n_3786),
.C(n_3784),
.D(n_3785),
.Y(n_16084)
);

NOR4xp25_ASAP7_75t_L g16085 ( 
.A(n_15964),
.B(n_3786),
.C(n_3784),
.D(n_3785),
.Y(n_16085)
);

OAI221xp5_ASAP7_75t_L g16086 ( 
.A1(n_16015),
.A2(n_3789),
.B1(n_3787),
.B2(n_3788),
.C(n_3791),
.Y(n_16086)
);

INVx1_ASAP7_75t_L g16087 ( 
.A(n_16015),
.Y(n_16087)
);

OR2x6_ASAP7_75t_L g16088 ( 
.A(n_16071),
.B(n_3787),
.Y(n_16088)
);

INVx1_ASAP7_75t_L g16089 ( 
.A(n_16077),
.Y(n_16089)
);

NOR3xp33_ASAP7_75t_L g16090 ( 
.A(n_16067),
.B(n_3788),
.C(n_3789),
.Y(n_16090)
);

O2A1O1Ixp33_ASAP7_75t_L g16091 ( 
.A1(n_16087),
.A2(n_3793),
.B(n_3791),
.C(n_3792),
.Y(n_16091)
);

XNOR2xp5_ASAP7_75t_L g16092 ( 
.A(n_16021),
.B(n_3792),
.Y(n_16092)
);

HB1xp67_ASAP7_75t_L g16093 ( 
.A(n_16083),
.Y(n_16093)
);

NAND3xp33_ASAP7_75t_L g16094 ( 
.A(n_16018),
.B(n_3794),
.C(n_3795),
.Y(n_16094)
);

XOR2xp5_ASAP7_75t_L g16095 ( 
.A(n_16031),
.B(n_3794),
.Y(n_16095)
);

AOI21xp33_ASAP7_75t_SL g16096 ( 
.A1(n_16020),
.A2(n_16023),
.B(n_16028),
.Y(n_16096)
);

NAND4xp25_ASAP7_75t_L g16097 ( 
.A(n_16036),
.B(n_16046),
.C(n_16037),
.D(n_16062),
.Y(n_16097)
);

INVx1_ASAP7_75t_L g16098 ( 
.A(n_16052),
.Y(n_16098)
);

XNOR2xp5_ASAP7_75t_L g16099 ( 
.A(n_16053),
.B(n_3796),
.Y(n_16099)
);

AO22x2_ASAP7_75t_L g16100 ( 
.A1(n_16038),
.A2(n_3798),
.B1(n_3796),
.B2(n_3797),
.Y(n_16100)
);

AOI211xp5_ASAP7_75t_L g16101 ( 
.A1(n_16059),
.A2(n_3800),
.B(n_3797),
.C(n_3799),
.Y(n_16101)
);

OAI22xp5_ASAP7_75t_L g16102 ( 
.A1(n_16082),
.A2(n_16034),
.B1(n_16044),
.B2(n_16049),
.Y(n_16102)
);

OAI22x1_ASAP7_75t_SL g16103 ( 
.A1(n_16057),
.A2(n_3802),
.B1(n_3799),
.B2(n_3801),
.Y(n_16103)
);

INVx2_ASAP7_75t_L g16104 ( 
.A(n_16078),
.Y(n_16104)
);

INVx2_ASAP7_75t_L g16105 ( 
.A(n_16048),
.Y(n_16105)
);

INVx2_ASAP7_75t_L g16106 ( 
.A(n_16035),
.Y(n_16106)
);

AOI22xp5_ASAP7_75t_L g16107 ( 
.A1(n_16030),
.A2(n_3803),
.B1(n_3801),
.B2(n_3802),
.Y(n_16107)
);

NOR2x1_ASAP7_75t_L g16108 ( 
.A(n_16050),
.B(n_3803),
.Y(n_16108)
);

INVx2_ASAP7_75t_SL g16109 ( 
.A(n_16019),
.Y(n_16109)
);

INVx1_ASAP7_75t_L g16110 ( 
.A(n_16043),
.Y(n_16110)
);

AND2x4_ASAP7_75t_L g16111 ( 
.A(n_16041),
.B(n_3804),
.Y(n_16111)
);

AOI22xp5_ASAP7_75t_L g16112 ( 
.A1(n_16047),
.A2(n_3806),
.B1(n_3804),
.B2(n_3805),
.Y(n_16112)
);

INVx1_ASAP7_75t_L g16113 ( 
.A(n_16055),
.Y(n_16113)
);

INVx2_ASAP7_75t_L g16114 ( 
.A(n_16025),
.Y(n_16114)
);

AOI222xp33_ASAP7_75t_SL g16115 ( 
.A1(n_16054),
.A2(n_16080),
.B1(n_16061),
.B2(n_16045),
.C1(n_16058),
.C2(n_16063),
.Y(n_16115)
);

OAI22xp5_ASAP7_75t_L g16116 ( 
.A1(n_16024),
.A2(n_3807),
.B1(n_3805),
.B2(n_3806),
.Y(n_16116)
);

AOI22xp5_ASAP7_75t_L g16117 ( 
.A1(n_16033),
.A2(n_3809),
.B1(n_3807),
.B2(n_3808),
.Y(n_16117)
);

AND2x2_ASAP7_75t_L g16118 ( 
.A(n_16055),
.B(n_3808),
.Y(n_16118)
);

AO22x2_ASAP7_75t_L g16119 ( 
.A1(n_16042),
.A2(n_3811),
.B1(n_3809),
.B2(n_3810),
.Y(n_16119)
);

NAND3xp33_ASAP7_75t_L g16120 ( 
.A(n_16051),
.B(n_3811),
.C(n_3812),
.Y(n_16120)
);

NOR2xp33_ASAP7_75t_R g16121 ( 
.A(n_16040),
.B(n_4095),
.Y(n_16121)
);

INVx1_ASAP7_75t_L g16122 ( 
.A(n_16027),
.Y(n_16122)
);

BUFx2_ASAP7_75t_L g16123 ( 
.A(n_16064),
.Y(n_16123)
);

INVx2_ASAP7_75t_L g16124 ( 
.A(n_16066),
.Y(n_16124)
);

AOI211xp5_ASAP7_75t_L g16125 ( 
.A1(n_16085),
.A2(n_3814),
.B(n_3812),
.C(n_3813),
.Y(n_16125)
);

XNOR2x1_ASAP7_75t_L g16126 ( 
.A(n_16039),
.B(n_3813),
.Y(n_16126)
);

AOI21xp5_ASAP7_75t_L g16127 ( 
.A1(n_16079),
.A2(n_3815),
.B(n_3816),
.Y(n_16127)
);

OAI22xp33_ASAP7_75t_L g16128 ( 
.A1(n_16072),
.A2(n_16056),
.B1(n_16084),
.B2(n_16073),
.Y(n_16128)
);

OAI22xp5_ASAP7_75t_L g16129 ( 
.A1(n_16039),
.A2(n_3817),
.B1(n_3815),
.B2(n_3816),
.Y(n_16129)
);

OAI22xp5_ASAP7_75t_L g16130 ( 
.A1(n_16074),
.A2(n_3820),
.B1(n_3818),
.B2(n_3819),
.Y(n_16130)
);

NOR2xp33_ASAP7_75t_L g16131 ( 
.A(n_16081),
.B(n_4101),
.Y(n_16131)
);

AOI21xp5_ASAP7_75t_L g16132 ( 
.A1(n_16032),
.A2(n_3819),
.B(n_3820),
.Y(n_16132)
);

INVx1_ASAP7_75t_SL g16133 ( 
.A(n_16093),
.Y(n_16133)
);

OAI22xp5_ASAP7_75t_SL g16134 ( 
.A1(n_16098),
.A2(n_16086),
.B1(n_16065),
.B2(n_16076),
.Y(n_16134)
);

AOI211x1_ASAP7_75t_L g16135 ( 
.A1(n_16089),
.A2(n_16029),
.B(n_16070),
.C(n_16060),
.Y(n_16135)
);

INVx1_ASAP7_75t_L g16136 ( 
.A(n_16096),
.Y(n_16136)
);

INVx2_ASAP7_75t_L g16137 ( 
.A(n_16104),
.Y(n_16137)
);

INVx1_ASAP7_75t_L g16138 ( 
.A(n_16110),
.Y(n_16138)
);

BUFx6f_ASAP7_75t_L g16139 ( 
.A(n_16105),
.Y(n_16139)
);

INVx2_ASAP7_75t_L g16140 ( 
.A(n_16123),
.Y(n_16140)
);

NAND3xp33_ASAP7_75t_L g16141 ( 
.A(n_16097),
.B(n_16113),
.C(n_16114),
.Y(n_16141)
);

INVx1_ASAP7_75t_L g16142 ( 
.A(n_16102),
.Y(n_16142)
);

NAND3x1_ASAP7_75t_L g16143 ( 
.A(n_16122),
.B(n_16022),
.C(n_16069),
.Y(n_16143)
);

INVx1_ASAP7_75t_L g16144 ( 
.A(n_16106),
.Y(n_16144)
);

INVx2_ASAP7_75t_L g16145 ( 
.A(n_16126),
.Y(n_16145)
);

INVx2_ASAP7_75t_L g16146 ( 
.A(n_16124),
.Y(n_16146)
);

INVx2_ASAP7_75t_L g16147 ( 
.A(n_16111),
.Y(n_16147)
);

INVx2_ASAP7_75t_L g16148 ( 
.A(n_16118),
.Y(n_16148)
);

OAI22xp5_ASAP7_75t_SL g16149 ( 
.A1(n_16109),
.A2(n_16092),
.B1(n_16131),
.B2(n_16095),
.Y(n_16149)
);

INVx3_ASAP7_75t_L g16150 ( 
.A(n_16088),
.Y(n_16150)
);

NAND2xp5_ASAP7_75t_L g16151 ( 
.A(n_16128),
.B(n_16026),
.Y(n_16151)
);

XNOR2x1_ASAP7_75t_L g16152 ( 
.A(n_16108),
.B(n_16075),
.Y(n_16152)
);

BUFx2_ASAP7_75t_L g16153 ( 
.A(n_16121),
.Y(n_16153)
);

HB1xp67_ASAP7_75t_L g16154 ( 
.A(n_16099),
.Y(n_16154)
);

INVxp33_ASAP7_75t_SL g16155 ( 
.A(n_16116),
.Y(n_16155)
);

NOR3x1_ASAP7_75t_L g16156 ( 
.A(n_16120),
.B(n_16075),
.C(n_16068),
.Y(n_16156)
);

XNOR2xp5_ASAP7_75t_L g16157 ( 
.A(n_16125),
.B(n_3822),
.Y(n_16157)
);

INVx1_ASAP7_75t_L g16158 ( 
.A(n_16119),
.Y(n_16158)
);

INVx1_ASAP7_75t_L g16159 ( 
.A(n_16119),
.Y(n_16159)
);

INVx1_ASAP7_75t_L g16160 ( 
.A(n_16112),
.Y(n_16160)
);

XOR2x2_ASAP7_75t_L g16161 ( 
.A(n_16117),
.B(n_3821),
.Y(n_16161)
);

BUFx2_ASAP7_75t_L g16162 ( 
.A(n_16088),
.Y(n_16162)
);

CKINVDCx20_ASAP7_75t_R g16163 ( 
.A(n_16133),
.Y(n_16163)
);

AO21x1_ASAP7_75t_L g16164 ( 
.A1(n_16136),
.A2(n_16129),
.B(n_16132),
.Y(n_16164)
);

INVx2_ASAP7_75t_L g16165 ( 
.A(n_16140),
.Y(n_16165)
);

NAND4xp25_ASAP7_75t_L g16166 ( 
.A(n_16141),
.B(n_16127),
.C(n_16090),
.D(n_16107),
.Y(n_16166)
);

INVx1_ASAP7_75t_L g16167 ( 
.A(n_16138),
.Y(n_16167)
);

INVxp67_ASAP7_75t_SL g16168 ( 
.A(n_16139),
.Y(n_16168)
);

HB1xp67_ASAP7_75t_L g16169 ( 
.A(n_16139),
.Y(n_16169)
);

AOI21x1_ASAP7_75t_L g16170 ( 
.A1(n_16146),
.A2(n_16130),
.B(n_16094),
.Y(n_16170)
);

AND5x1_ASAP7_75t_L g16171 ( 
.A(n_16137),
.B(n_16115),
.C(n_16091),
.D(n_16101),
.E(n_16103),
.Y(n_16171)
);

HB1xp67_ASAP7_75t_L g16172 ( 
.A(n_16147),
.Y(n_16172)
);

INVx3_ASAP7_75t_SL g16173 ( 
.A(n_16148),
.Y(n_16173)
);

INVx1_ASAP7_75t_L g16174 ( 
.A(n_16144),
.Y(n_16174)
);

INVx1_ASAP7_75t_L g16175 ( 
.A(n_16142),
.Y(n_16175)
);

NAND3xp33_ASAP7_75t_L g16176 ( 
.A(n_16162),
.B(n_16100),
.C(n_3821),
.Y(n_16176)
);

XNOR2xp5_ASAP7_75t_L g16177 ( 
.A(n_16152),
.B(n_16100),
.Y(n_16177)
);

NOR2xp33_ASAP7_75t_L g16178 ( 
.A(n_16150),
.B(n_3823),
.Y(n_16178)
);

AOI22xp5_ASAP7_75t_L g16179 ( 
.A1(n_16158),
.A2(n_3824),
.B1(n_3822),
.B2(n_3823),
.Y(n_16179)
);

INVx1_ASAP7_75t_L g16180 ( 
.A(n_16159),
.Y(n_16180)
);

INVx1_ASAP7_75t_L g16181 ( 
.A(n_16151),
.Y(n_16181)
);

NAND2xp5_ASAP7_75t_L g16182 ( 
.A(n_16145),
.B(n_3824),
.Y(n_16182)
);

INVx2_ASAP7_75t_L g16183 ( 
.A(n_16153),
.Y(n_16183)
);

AOI22xp5_ASAP7_75t_L g16184 ( 
.A1(n_16149),
.A2(n_16154),
.B1(n_16155),
.B2(n_16143),
.Y(n_16184)
);

OAI22xp33_ASAP7_75t_L g16185 ( 
.A1(n_16165),
.A2(n_16160),
.B1(n_16156),
.B2(n_16135),
.Y(n_16185)
);

INVx1_ASAP7_75t_L g16186 ( 
.A(n_16169),
.Y(n_16186)
);

HB1xp67_ASAP7_75t_L g16187 ( 
.A(n_16175),
.Y(n_16187)
);

BUFx2_ASAP7_75t_L g16188 ( 
.A(n_16163),
.Y(n_16188)
);

OAI31xp33_ASAP7_75t_SL g16189 ( 
.A1(n_16168),
.A2(n_16157),
.A3(n_16134),
.B(n_16161),
.Y(n_16189)
);

AOI22xp33_ASAP7_75t_L g16190 ( 
.A1(n_16167),
.A2(n_3827),
.B1(n_3825),
.B2(n_3826),
.Y(n_16190)
);

AOI22xp5_ASAP7_75t_L g16191 ( 
.A1(n_16174),
.A2(n_3827),
.B1(n_3825),
.B2(n_3826),
.Y(n_16191)
);

AOI22xp33_ASAP7_75t_L g16192 ( 
.A1(n_16172),
.A2(n_3830),
.B1(n_3828),
.B2(n_3829),
.Y(n_16192)
);

INVx1_ASAP7_75t_L g16193 ( 
.A(n_16181),
.Y(n_16193)
);

AOI22xp5_ASAP7_75t_L g16194 ( 
.A1(n_16183),
.A2(n_3831),
.B1(n_3828),
.B2(n_3829),
.Y(n_16194)
);

AOI22xp33_ASAP7_75t_L g16195 ( 
.A1(n_16173),
.A2(n_3833),
.B1(n_3831),
.B2(n_3832),
.Y(n_16195)
);

HB1xp67_ASAP7_75t_L g16196 ( 
.A(n_16180),
.Y(n_16196)
);

AOI22xp5_ASAP7_75t_L g16197 ( 
.A1(n_16184),
.A2(n_3834),
.B1(n_3832),
.B2(n_3833),
.Y(n_16197)
);

HB1xp67_ASAP7_75t_L g16198 ( 
.A(n_16177),
.Y(n_16198)
);

INVx1_ASAP7_75t_L g16199 ( 
.A(n_16176),
.Y(n_16199)
);

OR2x2_ASAP7_75t_L g16200 ( 
.A(n_16182),
.B(n_3835),
.Y(n_16200)
);

INVx2_ASAP7_75t_L g16201 ( 
.A(n_16170),
.Y(n_16201)
);

OAI22xp5_ASAP7_75t_L g16202 ( 
.A1(n_16178),
.A2(n_16179),
.B1(n_16171),
.B2(n_16164),
.Y(n_16202)
);

AOI22xp5_ASAP7_75t_L g16203 ( 
.A1(n_16166),
.A2(n_3837),
.B1(n_3835),
.B2(n_3836),
.Y(n_16203)
);

HB1xp67_ASAP7_75t_L g16204 ( 
.A(n_16169),
.Y(n_16204)
);

HB1xp67_ASAP7_75t_L g16205 ( 
.A(n_16169),
.Y(n_16205)
);

BUFx8_ASAP7_75t_L g16206 ( 
.A(n_16165),
.Y(n_16206)
);

AO21x2_ASAP7_75t_L g16207 ( 
.A1(n_16193),
.A2(n_3844),
.B(n_3836),
.Y(n_16207)
);

OAI21x1_ASAP7_75t_SL g16208 ( 
.A1(n_16186),
.A2(n_4115),
.B(n_3837),
.Y(n_16208)
);

NAND2xp5_ASAP7_75t_L g16209 ( 
.A(n_16204),
.B(n_3838),
.Y(n_16209)
);

AOI22xp33_ASAP7_75t_L g16210 ( 
.A1(n_16205),
.A2(n_3840),
.B1(n_3838),
.B2(n_3839),
.Y(n_16210)
);

INVx2_ASAP7_75t_L g16211 ( 
.A(n_16206),
.Y(n_16211)
);

OAI22xp5_ASAP7_75t_L g16212 ( 
.A1(n_16187),
.A2(n_3850),
.B1(n_3858),
.B2(n_3839),
.Y(n_16212)
);

INVx1_ASAP7_75t_L g16213 ( 
.A(n_16206),
.Y(n_16213)
);

NAND2xp5_ASAP7_75t_L g16214 ( 
.A(n_16188),
.B(n_3840),
.Y(n_16214)
);

INVx1_ASAP7_75t_L g16215 ( 
.A(n_16196),
.Y(n_16215)
);

HB1xp67_ASAP7_75t_L g16216 ( 
.A(n_16201),
.Y(n_16216)
);

OAI22x1_ASAP7_75t_L g16217 ( 
.A1(n_16198),
.A2(n_3843),
.B1(n_3841),
.B2(n_3842),
.Y(n_16217)
);

OAI21x1_ASAP7_75t_L g16218 ( 
.A1(n_16202),
.A2(n_3841),
.B(n_3843),
.Y(n_16218)
);

INVx1_ASAP7_75t_L g16219 ( 
.A(n_16185),
.Y(n_16219)
);

AOI221xp5_ASAP7_75t_L g16220 ( 
.A1(n_16199),
.A2(n_3849),
.B1(n_3845),
.B2(n_3846),
.C(n_3851),
.Y(n_16220)
);

INVx1_ASAP7_75t_SL g16221 ( 
.A(n_16200),
.Y(n_16221)
);

OAI21xp5_ASAP7_75t_L g16222 ( 
.A1(n_16203),
.A2(n_3849),
.B(n_3851),
.Y(n_16222)
);

NAND3xp33_ASAP7_75t_L g16223 ( 
.A(n_16189),
.B(n_3860),
.C(n_3852),
.Y(n_16223)
);

OAI21x1_ASAP7_75t_L g16224 ( 
.A1(n_16195),
.A2(n_3852),
.B(n_3853),
.Y(n_16224)
);

HB1xp67_ASAP7_75t_L g16225 ( 
.A(n_16215),
.Y(n_16225)
);

OAI22xp33_ASAP7_75t_L g16226 ( 
.A1(n_16219),
.A2(n_16197),
.B1(n_16194),
.B2(n_16191),
.Y(n_16226)
);

OAI22xp5_ASAP7_75t_SL g16227 ( 
.A1(n_16213),
.A2(n_16190),
.B1(n_16192),
.B2(n_3855),
.Y(n_16227)
);

OAI22xp5_ASAP7_75t_L g16228 ( 
.A1(n_16216),
.A2(n_3855),
.B1(n_3853),
.B2(n_3854),
.Y(n_16228)
);

INVxp67_ASAP7_75t_L g16229 ( 
.A(n_16211),
.Y(n_16229)
);

HB1xp67_ASAP7_75t_L g16230 ( 
.A(n_16221),
.Y(n_16230)
);

AOI22xp5_ASAP7_75t_L g16231 ( 
.A1(n_16207),
.A2(n_3858),
.B1(n_3856),
.B2(n_3857),
.Y(n_16231)
);

BUFx2_ASAP7_75t_L g16232 ( 
.A(n_16222),
.Y(n_16232)
);

OAI22xp5_ASAP7_75t_SL g16233 ( 
.A1(n_16214),
.A2(n_3860),
.B1(n_3857),
.B2(n_3859),
.Y(n_16233)
);

CKINVDCx5p33_ASAP7_75t_R g16234 ( 
.A(n_16209),
.Y(n_16234)
);

OAI22xp5_ASAP7_75t_L g16235 ( 
.A1(n_16223),
.A2(n_3862),
.B1(n_3859),
.B2(n_3861),
.Y(n_16235)
);

INVx4_ASAP7_75t_L g16236 ( 
.A(n_16208),
.Y(n_16236)
);

BUFx2_ASAP7_75t_L g16237 ( 
.A(n_16218),
.Y(n_16237)
);

NAND5xp2_ASAP7_75t_L g16238 ( 
.A(n_16220),
.B(n_3863),
.C(n_3861),
.D(n_3862),
.E(n_3864),
.Y(n_16238)
);

NAND2xp5_ASAP7_75t_SL g16239 ( 
.A(n_16229),
.B(n_16217),
.Y(n_16239)
);

NAND2xp5_ASAP7_75t_L g16240 ( 
.A(n_16225),
.B(n_16224),
.Y(n_16240)
);

AOI22xp33_ASAP7_75t_L g16241 ( 
.A1(n_16230),
.A2(n_16212),
.B1(n_16210),
.B2(n_3866),
.Y(n_16241)
);

AOI22xp33_ASAP7_75t_L g16242 ( 
.A1(n_16237),
.A2(n_3866),
.B1(n_3863),
.B2(n_3865),
.Y(n_16242)
);

NOR2xp33_ASAP7_75t_L g16243 ( 
.A(n_16236),
.B(n_3865),
.Y(n_16243)
);

OAI22xp5_ASAP7_75t_L g16244 ( 
.A1(n_16236),
.A2(n_3869),
.B1(n_3867),
.B2(n_3868),
.Y(n_16244)
);

HB1xp67_ASAP7_75t_L g16245 ( 
.A(n_16234),
.Y(n_16245)
);

OAI21xp5_ASAP7_75t_L g16246 ( 
.A1(n_16226),
.A2(n_3876),
.B(n_3868),
.Y(n_16246)
);

AOI22xp33_ASAP7_75t_L g16247 ( 
.A1(n_16232),
.A2(n_3871),
.B1(n_3869),
.B2(n_3870),
.Y(n_16247)
);

AOI22xp33_ASAP7_75t_L g16248 ( 
.A1(n_16233),
.A2(n_3872),
.B1(n_3870),
.B2(n_3871),
.Y(n_16248)
);

NAND2xp5_ASAP7_75t_L g16249 ( 
.A(n_16231),
.B(n_4115),
.Y(n_16249)
);

INVx2_ASAP7_75t_L g16250 ( 
.A(n_16245),
.Y(n_16250)
);

INVx1_ASAP7_75t_L g16251 ( 
.A(n_16240),
.Y(n_16251)
);

XOR2xp5_ASAP7_75t_L g16252 ( 
.A(n_16239),
.B(n_16227),
.Y(n_16252)
);

INVx1_ASAP7_75t_L g16253 ( 
.A(n_16249),
.Y(n_16253)
);

OAI22x1_ASAP7_75t_L g16254 ( 
.A1(n_16243),
.A2(n_16238),
.B1(n_16235),
.B2(n_16228),
.Y(n_16254)
);

AOI22xp5_ASAP7_75t_L g16255 ( 
.A1(n_16241),
.A2(n_3880),
.B1(n_3888),
.B2(n_3872),
.Y(n_16255)
);

AOI31xp33_ASAP7_75t_L g16256 ( 
.A1(n_16251),
.A2(n_16248),
.A3(n_16246),
.B(n_16244),
.Y(n_16256)
);

NAND2xp5_ASAP7_75t_L g16257 ( 
.A(n_16250),
.B(n_16242),
.Y(n_16257)
);

OAI21xp5_ASAP7_75t_L g16258 ( 
.A1(n_16252),
.A2(n_16253),
.B(n_16255),
.Y(n_16258)
);

AOI22xp33_ASAP7_75t_L g16259 ( 
.A1(n_16254),
.A2(n_16247),
.B1(n_3875),
.B2(n_3873),
.Y(n_16259)
);

AOI22xp33_ASAP7_75t_L g16260 ( 
.A1(n_16250),
.A2(n_3875),
.B1(n_3873),
.B2(n_3874),
.Y(n_16260)
);

NAND2xp5_ASAP7_75t_L g16261 ( 
.A(n_16250),
.B(n_3874),
.Y(n_16261)
);

AOI21xp5_ASAP7_75t_L g16262 ( 
.A1(n_16257),
.A2(n_3876),
.B(n_3877),
.Y(n_16262)
);

CKINVDCx20_ASAP7_75t_R g16263 ( 
.A(n_16258),
.Y(n_16263)
);

OAI22xp5_ASAP7_75t_L g16264 ( 
.A1(n_16259),
.A2(n_3879),
.B1(n_3877),
.B2(n_3878),
.Y(n_16264)
);

OAI22xp33_ASAP7_75t_L g16265 ( 
.A1(n_16256),
.A2(n_3880),
.B1(n_3878),
.B2(n_3879),
.Y(n_16265)
);

INVx1_ASAP7_75t_L g16266 ( 
.A(n_16263),
.Y(n_16266)
);

OAI21xp5_ASAP7_75t_L g16267 ( 
.A1(n_16264),
.A2(n_16261),
.B(n_16260),
.Y(n_16267)
);

AOI22xp33_ASAP7_75t_L g16268 ( 
.A1(n_16266),
.A2(n_16262),
.B1(n_16265),
.B2(n_3883),
.Y(n_16268)
);

AOI322xp5_ASAP7_75t_L g16269 ( 
.A1(n_16267),
.A2(n_3886),
.A3(n_3885),
.B1(n_3883),
.B2(n_3881),
.C1(n_3882),
.C2(n_3884),
.Y(n_16269)
);

OR2x6_ASAP7_75t_L g16270 ( 
.A(n_16268),
.B(n_4100),
.Y(n_16270)
);

NAND2xp5_ASAP7_75t_L g16271 ( 
.A(n_16269),
.B(n_3881),
.Y(n_16271)
);

AOI22xp5_ASAP7_75t_L g16272 ( 
.A1(n_16270),
.A2(n_3886),
.B1(n_3882),
.B2(n_3885),
.Y(n_16272)
);

AOI22xp33_ASAP7_75t_SL g16273 ( 
.A1(n_16271),
.A2(n_3893),
.B1(n_3895),
.B2(n_3887),
.Y(n_16273)
);

AOI22xp5_ASAP7_75t_L g16274 ( 
.A1(n_16273),
.A2(n_3890),
.B1(n_3887),
.B2(n_3889),
.Y(n_16274)
);

AOI211xp5_ASAP7_75t_L g16275 ( 
.A1(n_16274),
.A2(n_16272),
.B(n_3891),
.C(n_3889),
.Y(n_16275)
);


endmodule