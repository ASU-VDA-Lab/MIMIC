module real_jpeg_6185_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_1),
.A2(n_151),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_1),
.A2(n_250),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_1),
.A2(n_124),
.B1(n_250),
.B2(n_364),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_1),
.A2(n_250),
.B1(n_386),
.B2(n_389),
.Y(n_385)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_53),
.B1(n_121),
.B2(n_124),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_3),
.A2(n_53),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_3),
.B(n_70),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_3),
.A2(n_352),
.B(n_354),
.C(n_358),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_3),
.B(n_376),
.C(n_378),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_3),
.B(n_21),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_3),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_3),
.B(n_109),
.Y(n_415)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_5),
.Y(n_198)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_5),
.Y(n_403)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_5),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_6),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_7),
.Y(n_281)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_9),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_10),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_11),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_12),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_12),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_12),
.A2(n_92),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_12),
.A2(n_92),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_12),
.A2(n_92),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_13),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_13),
.A2(n_87),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_87),
.B1(n_210),
.B2(n_214),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_13),
.A2(n_87),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_448),
.B(n_451),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_167),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_165),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_18),
.B(n_141),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_96),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_55),
.B1(n_56),
.B2(n_95),
.Y(n_19)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_20),
.A2(n_95),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_33),
.B(n_49),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_21),
.B(n_129),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_21),
.A2(n_127),
.B(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_21),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_22),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_25),
.Y(n_356)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_27),
.Y(n_188)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_27),
.Y(n_215)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_27),
.Y(n_366)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_29),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_32),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_33),
.A2(n_157),
.B(n_163),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_33),
.B(n_49),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_33),
.B(n_269),
.Y(n_296)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_34),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_41),
.Y(n_159)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_42),
.Y(n_134)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_42),
.Y(n_279)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_49),
.Y(n_136)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_53),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_53),
.B(n_153),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g354 ( 
.A1(n_53),
.A2(n_355),
.B(n_357),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_80),
.B(n_88),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_57),
.A2(n_139),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_58),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_58),
.B(n_249),
.Y(n_248)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_70),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_68),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_63),
.Y(n_287)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_70),
.B(n_150),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_70),
.B(n_249),
.Y(n_264)
);

AO22x1_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_73),
.Y(n_285)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_77),
.Y(n_271)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_88),
.B(n_248),
.Y(n_312)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_95),
.B(n_321),
.C(n_323),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_126),
.C(n_137),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_97),
.A2(n_126),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_97),
.B(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_97),
.A2(n_147),
.B1(n_266),
.B2(n_274),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_97),
.B(n_263),
.C(n_266),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_118),
.B(n_119),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_98),
.A2(n_209),
.B(n_216),
.Y(n_208)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_99),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_99),
.B(n_120),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_99),
.B(n_363),
.Y(n_362)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_110),
.B1(n_112),
.B2(n_116),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_108),
.Y(n_213)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_109),
.B(n_184),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_109),
.B(n_363),
.Y(n_380)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_113),
.Y(n_389)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_115),
.Y(n_242)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_117),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_117),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_118),
.B(n_119),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_118),
.A2(n_183),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_123),
.Y(n_374)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_134),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_135),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_140),
.B(n_264),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.C(n_155),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_142),
.A2(n_143),
.B1(n_148),
.B2(n_175),
.Y(n_254)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.C(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_149),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_152),
.Y(n_283)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_155),
.B(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_158),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_164),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_164),
.B(n_296),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_256),
.B(n_444),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_252),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_220),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_171),
.B(n_220),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_190),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_178),
.B2(n_179),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_174),
.B(n_178),
.C(n_190),
.Y(n_255)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_180),
.B(n_189),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_181),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_183),
.B(n_380),
.Y(n_424)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_217),
.B(n_218),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_192),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_208),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_217),
.B1(n_218),
.B2(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_193),
.A2(n_208),
.B1(n_217),
.B2(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_193),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_193),
.A2(n_217),
.B1(n_351),
.B2(n_427),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_199),
.B(n_202),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_194),
.B(n_202),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_194),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_194),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_197),
.B(n_238),
.Y(n_301)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_205),
.Y(n_388)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_208),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g307 ( 
.A(n_216),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_216),
.B(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.C(n_227),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_221),
.A2(n_225),
.B1(n_226),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_221),
.Y(n_336)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_227),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_244),
.C(n_246),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_228),
.A2(n_229),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_243),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_230),
.B(n_243),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_231),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

INVx3_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_236),
.B(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_237),
.A2(n_289),
.B(n_293),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_244),
.B(n_246),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_245),
.B(n_268),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_252),
.A2(n_446),
.B(n_447),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_253),
.B(n_255),
.Y(n_447)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_436),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_325),
.C(n_341),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_315),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_302),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_261),
.B(n_302),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_275),
.C(n_294),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_262),
.B(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_275),
.A2(n_276),
.B1(n_294),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_288),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_277),
.B(n_288),
.Y(n_310)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_280),
.A3(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_301),
.B(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.C(n_299),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_299),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_300),
.B(n_401),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_301),
.B(n_384),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_302),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_302),
.B(n_316),
.Y(n_440)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.CI(n_309),
.CON(n_302),
.SN(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_307),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_308),
.B(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_315),
.A2(n_439),
.B(n_440),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_319),
.C(n_320),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_337),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_326),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_334),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_327),
.B(n_334),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.C(n_333),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_331),
.Y(n_339)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_338),
.B(n_340),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_367),
.B(n_435),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_346),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_343),
.B(n_346),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.C(n_359),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_347),
.B(n_431),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_350),
.A2(n_359),
.B1(n_360),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_429),
.B(n_434),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_419),
.B(n_428),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_395),
.B(n_418),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_381),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_381),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_379),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_372),
.A2(n_373),
.B1(n_379),
.B2(n_398),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_390),
.Y(n_381)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_391),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_391),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_392),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_393),
.C(n_421),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_396),
.A2(n_404),
.B(n_417),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_399),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_399),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_413),
.B(n_416),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_412),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_414),
.B(n_415),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_422),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_425),
.C(n_426),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_433),
.Y(n_434)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g436 ( 
.A1(n_437),
.A2(n_438),
.B(n_441),
.C(n_442),
.D(n_443),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_452),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx13_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);


endmodule