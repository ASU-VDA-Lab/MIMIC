module fake_netlist_1_2051_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
INVx1_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVxp67_ASAP7_75t_SL g4 ( .A(n_2), .Y(n_4) );
AND2x4_ASAP7_75t_L g5 ( .A(n_1), .B(n_0), .Y(n_5) );
AO31x2_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .A3(n_1), .B(n_5), .Y(n_6) );
AO31x2_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .A3(n_5), .B(n_4), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_5), .Y(n_8) );
BUFx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_5), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
NAND2xp33_ASAP7_75t_SL g13 ( .A(n_12), .B(n_7), .Y(n_13) );
AND3x1_ASAP7_75t_L g14 ( .A(n_12), .B(n_6), .C(n_11), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_13), .B(n_6), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_6), .Y(n_16) );
INVx3_ASAP7_75t_SL g17 ( .A(n_16), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
endmodule