module real_jpeg_5512_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_0),
.A2(n_52),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_0),
.A2(n_52),
.B1(n_201),
.B2(n_391),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_0),
.A2(n_52),
.B1(n_358),
.B2(n_404),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_1),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_1),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_1),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_2),
.A2(n_167),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_2),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_2),
.A2(n_202),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_2),
.A2(n_202),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_2),
.A2(n_202),
.B1(n_431),
.B2(n_433),
.Y(n_430)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_3),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_3),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g432 ( 
.A(n_3),
.Y(n_432)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_3),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_4),
.A2(n_60),
.B1(n_340),
.B2(n_343),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_4),
.A2(n_60),
.B1(n_162),
.B2(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_4),
.A2(n_60),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_5),
.A2(n_115),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_5),
.A2(n_169),
.B1(n_188),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_5),
.A2(n_169),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_5),
.A2(n_49),
.B1(n_169),
.B2(n_354),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_6),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_6),
.A2(n_92),
.B1(n_135),
.B2(n_140),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_6),
.A2(n_92),
.B1(n_376),
.B2(n_378),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_6),
.A2(n_92),
.B1(n_114),
.B2(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_8),
.Y(n_535)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_13),
.A2(n_160),
.B1(n_162),
.B2(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_13),
.B(n_117),
.C(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_13),
.B(n_79),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_13),
.B(n_128),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_13),
.B(n_89),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_179),
.B1(n_180),
.B2(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_14),
.A2(n_114),
.B1(n_184),
.B2(n_246),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_14),
.A2(n_184),
.B1(n_358),
.B2(n_360),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_14),
.A2(n_184),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_15),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_16),
.A2(n_43),
.B1(n_95),
.B2(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_16),
.A2(n_98),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_16),
.A2(n_58),
.B1(n_98),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_16),
.A2(n_98),
.B1(n_217),
.B2(n_384),
.Y(n_383)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_18),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_18),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_18),
.A2(n_201),
.B1(n_267),
.B2(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_18),
.A2(n_267),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_L g460 ( 
.A1(n_18),
.A2(n_267),
.B1(n_322),
.B2(n_431),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_534),
.B(n_536),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_149),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_147),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_144),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_23),
.B(n_144),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_133),
.C(n_141),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_24),
.A2(n_25),
.B1(n_530),
.B2(n_531),
.Y(n_529)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_61),
.C(n_99),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_26),
.B(n_522),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_53),
.B1(n_55),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_27),
.A2(n_53),
.B1(n_134),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_27),
.A2(n_352),
.B(n_407),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_27),
.A2(n_38),
.B1(n_407),
.B2(n_430),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_27),
.A2(n_48),
.B1(n_53),
.B2(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_28),
.A2(n_350),
.B(n_351),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_28),
.B(n_353),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_38),
.B(n_164),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_46),
.Y(n_38)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_39),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_41),
.Y(n_258)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_41),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_42),
.Y(n_330)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_42),
.Y(n_401)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_42),
.Y(n_404)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_43),
.A2(n_319),
.A3(n_323),
.B1(n_325),
.B2(n_331),
.Y(n_318)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_47),
.Y(n_327)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_SL g350 ( 
.A1(n_50),
.A2(n_164),
.B(n_331),
.Y(n_350)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_51),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_53),
.A2(n_430),
.B(n_461),
.Y(n_471)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_54),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_54),
.B(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_57),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_57),
.Y(n_354)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_61),
.A2(n_99),
.B1(n_100),
.B2(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_61),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_62),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_62),
.A2(n_93),
.B1(n_293),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_62),
.A2(n_93),
.B1(n_399),
.B2(n_405),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_62),
.A2(n_88),
.B1(n_93),
.B2(n_511),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_79),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_66),
.Y(n_276)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_68),
.Y(n_282)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_71),
.Y(n_363)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_77),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_78),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_78),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_78),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_78),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_79),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_79),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g435 ( 
.A1(n_79),
.A2(n_142),
.B1(n_300),
.B2(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_79),
.A2(n_142),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_83),
.Y(n_279)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_83),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_85),
.Y(n_396)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_93),
.B(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_93),
.A2(n_293),
.B(n_299),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_99),
.A2(n_100),
.B1(n_509),
.B2(n_510),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_99),
.B(n_506),
.C(n_509),
.Y(n_517)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_127),
.B(n_129),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_159),
.B(n_165),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_101),
.A2(n_127),
.B1(n_199),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_101),
.A2(n_165),
.B(n_245),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_101),
.A2(n_127),
.B1(n_365),
.B2(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_102),
.B(n_166),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_102),
.A2(n_128),
.B1(n_390),
.B2(n_394),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_102),
.A2(n_128),
.B1(n_394),
.B2(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_102),
.A2(n_128),
.B1(n_413),
.B2(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_116),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_110),
.B2(n_114),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_106),
.Y(n_248)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_116),
.A2(n_199),
.B(n_203),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_121),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_123),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_123),
.Y(n_343)
);

BUFx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_124),
.Y(n_388)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_127),
.A2(n_203),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_129),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_132),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_133),
.B(n_141),
.Y(n_531)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_140),
.B(n_164),
.Y(n_331)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_140),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_142),
.A2(n_251),
.B(n_255),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_142),
.B(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_142),
.A2(n_255),
.B(n_474),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_528),
.B(n_533),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_500),
.B(n_525),
.Y(n_150)
);

OAI311xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_369),
.A3(n_476),
.B1(n_494),
.C1(n_495),
.Y(n_151)
);

AOI21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_312),
.B(n_368),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_284),
.B(n_311),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_239),
.B(n_283),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_206),
.B(n_238),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_176),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_157),
.B(n_176),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_170),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_158),
.A2(n_170),
.B1(n_171),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_164),
.A2(n_185),
.B(n_191),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_SL g251 ( 
.A1(n_164),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_167),
.Y(n_274)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_175),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_196),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_197),
.C(n_205),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_185),
.B(n_191),
.Y(n_177)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_183),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_185),
.A2(n_334),
.B1(n_335),
.B2(n_338),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_185),
.A2(n_375),
.B1(n_380),
.B2(n_383),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_185),
.A2(n_383),
.B(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_194),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_186),
.A2(n_265),
.B1(n_304),
.B2(n_309),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_186),
.A2(n_339),
.B1(n_419),
.B2(n_427),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_190),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_193),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_204),
.B2(n_205),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_228),
.B(n_237),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_214),
.B(n_227),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_212),
.Y(n_337)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_212),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_226),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_226),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_222),
.B(n_225),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_225),
.A2(n_264),
.B(n_271),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_235),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_241),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_262),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_249),
.B2(n_250),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_249),
.C(n_262),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_248),
.Y(n_416)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI32xp33_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_273),
.A3(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_272)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_272),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_285),
.B(n_286),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_310),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_290),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_302),
.C(n_303),
.Y(n_344)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

INVx4_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_313),
.B(n_314),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_347),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_315)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_332),
.B2(n_333),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_318),
.B(n_332),
.Y(n_472)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_344),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_344),
.B(n_345),
.C(n_347),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_355),
.B2(n_367),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_348),
.B(n_356),
.C(n_364),
.Y(n_485)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_364),
.Y(n_355)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_462),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_SL g495 ( 
.A1(n_370),
.A2(n_462),
.B(n_496),
.C(n_499),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_437),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_371),
.B(n_437),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_410),
.C(n_422),
.Y(n_371)
);

FAx1_ASAP7_75t_SL g475 ( 
.A(n_372),
.B(n_410),
.CI(n_422),
.CON(n_475),
.SN(n_475)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_397),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_373),
.B(n_398),
.C(n_406),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_389),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_374),
.B(n_389),
.Y(n_468)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_375),
.Y(n_427)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_406),
.Y(n_397)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_405),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_417),
.B2(n_421),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_417),
.Y(n_455)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_417),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_417),
.A2(n_421),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_417),
.A2(n_455),
.B(n_458),
.Y(n_503)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_428),
.C(n_435),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_423),
.B(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_426),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_428),
.A2(n_429),
.B1(n_435),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx8_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_435),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_438),
.B(n_441),
.C(n_453),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_453),
.B2(n_454),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_449),
.B(n_452),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_450),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_452),
.B(n_503),
.CI(n_504),
.CON(n_502),
.SN(n_502)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_452),
.B(n_503),
.C(n_504),
.Y(n_524)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_461),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_460),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_475),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_475),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.C(n_469),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_464),
.A2(n_465),
.B1(n_468),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_487),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.C(n_473),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_470),
.A2(n_471),
.B1(n_473),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_475),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_489),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_497),
.B(n_498),
.Y(n_496)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_486),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_486),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_483),
.C(n_485),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_492),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_483),
.A2(n_484),
.B1(n_485),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_485),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_491),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_514),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_513),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_502),
.B(n_513),
.Y(n_526)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_502),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_508),
.B2(n_512),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_505),
.A2(n_506),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_516),
.C(n_520),
.Y(n_532)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_508),
.Y(n_512)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_514),
.A2(n_526),
.B(n_527),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_524),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_524),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_532),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_532),
.Y(n_533)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx8_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx13_ASAP7_75t_L g537 ( 
.A(n_535),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_538),
.Y(n_536)
);


endmodule