module real_aes_17247_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_845, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_845;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g110 ( .A(n_0), .B(n_111), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_1), .A2(n_4), .B1(n_146), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_2), .A2(n_42), .B1(n_153), .B2(n_189), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_3), .A2(n_24), .B1(n_189), .B2(n_231), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_5), .A2(n_16), .B1(n_143), .B2(n_220), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_6), .A2(n_61), .B1(n_203), .B2(n_233), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_7), .A2(n_17), .B1(n_153), .B2(n_174), .Y(n_625) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_9), .A2(n_477), .B(n_834), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_10), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_11), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_12), .A2(n_18), .B1(n_202), .B2(n_205), .Y(n_201) );
BUFx2_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
OR2x2_ASAP7_75t_L g472 ( .A(n_13), .B(n_37), .Y(n_472) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_15), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_19), .A2(n_101), .B1(n_143), .B2(n_146), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_20), .A2(n_38), .B1(n_178), .B2(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_21), .B(n_144), .Y(n_175) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_22), .A2(n_57), .B(n_162), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_23), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_25), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_26), .B(n_150), .Y(n_545) );
INVx4_ASAP7_75t_R g593 ( .A(n_27), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_28), .A2(n_47), .B1(n_191), .B2(n_192), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_29), .A2(n_54), .B1(n_143), .B2(n_192), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_30), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_31), .B(n_178), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_32), .Y(n_254) );
INVx1_ASAP7_75t_L g524 ( .A(n_33), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_34), .B(n_189), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_SL g536 ( .A1(n_35), .A2(n_149), .B(n_153), .C(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_36), .A2(n_55), .B1(n_153), .B2(n_192), .Y(n_513) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_37), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_39), .A2(n_88), .B1(n_153), .B2(n_230), .Y(n_229) );
XOR2x2_ASAP7_75t_L g827 ( .A(n_40), .B(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_41), .A2(n_45), .B1(n_153), .B2(n_174), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_43), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_44), .A2(n_59), .B1(n_143), .B2(n_152), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_46), .A2(n_73), .B1(n_829), .B2(n_830), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_46), .Y(n_830) );
INVx1_ASAP7_75t_L g548 ( .A(n_48), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_49), .B(n_153), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_50), .Y(n_565) );
INVx2_ASAP7_75t_L g485 ( .A(n_51), .Y(n_485) );
INVx1_ASAP7_75t_L g113 ( .A(n_52), .Y(n_113) );
BUFx3_ASAP7_75t_L g494 ( .A(n_52), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_53), .A2(n_122), .B(n_473), .Y(n_121) );
AOI31xp33_ASAP7_75t_L g473 ( .A1(n_53), .A2(n_474), .A3(n_476), .B(n_477), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_56), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_58), .A2(n_89), .B1(n_153), .B2(n_192), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_60), .A2(n_68), .B1(n_125), .B2(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_60), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_62), .A2(n_77), .B1(n_152), .B2(n_191), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_63), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_64), .A2(n_79), .B1(n_153), .B2(n_174), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_65), .A2(n_100), .B1(n_143), .B2(n_205), .Y(n_251) );
AND2x4_ASAP7_75t_L g139 ( .A(n_66), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g162 ( .A(n_67), .Y(n_162) );
INVx1_ASAP7_75t_L g125 ( .A(n_68), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_69), .A2(n_92), .B1(n_191), .B2(n_192), .Y(n_520) );
AO22x1_ASAP7_75t_L g582 ( .A1(n_70), .A2(n_78), .B1(n_217), .B2(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g140 ( .A(n_71), .Y(n_140) );
AND2x2_ASAP7_75t_L g540 ( .A(n_72), .B(n_184), .Y(n_540) );
INVx1_ASAP7_75t_L g829 ( .A(n_73), .Y(n_829) );
INVx1_ASAP7_75t_L g842 ( .A(n_74), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_75), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_76), .B(n_233), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_80), .B(n_189), .Y(n_566) );
INVx2_ASAP7_75t_L g150 ( .A(n_81), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_82), .B(n_184), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_83), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_84), .A2(n_99), .B1(n_192), .B2(n_233), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_85), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_86), .B(n_160), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_87), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_90), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_91), .B(n_184), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_93), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_94), .B(n_184), .Y(n_562) );
INVx1_ASAP7_75t_L g115 ( .A(n_95), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_95), .B(n_470), .Y(n_469) );
NAND2xp33_ASAP7_75t_L g180 ( .A(n_96), .B(n_144), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g588 ( .A1(n_97), .A2(n_208), .B(n_233), .C(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g595 ( .A(n_98), .B(n_596), .Y(n_595) );
NAND2xp33_ASAP7_75t_L g570 ( .A(n_102), .B(n_179), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_120), .B(n_841), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx12f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx4_ASAP7_75t_L g843 ( .A(n_106), .Y(n_843) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_116), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .C(n_114), .Y(n_108) );
INVx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g470 ( .A(n_113), .Y(n_470) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g500 ( .A(n_115), .Y(n_500) );
NOR2x1p5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_481), .B(n_486), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_466), .Y(n_122) );
INVx1_ASAP7_75t_L g476 ( .A(n_123), .Y(n_476) );
XOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
INVx2_ASAP7_75t_L g501 ( .A(n_127), .Y(n_501) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_369), .Y(n_127) );
NAND4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_293), .C(n_324), .D(n_353), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_260), .Y(n_129) );
OAI322xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_196), .A3(n_225), .B1(n_238), .B2(n_246), .C1(n_255), .C2(n_257), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_132), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_166), .Y(n_132) );
AND2x2_ASAP7_75t_L g290 ( .A(n_133), .B(n_291), .Y(n_290) );
INVx4_ASAP7_75t_L g326 ( .A(n_133), .Y(n_326) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g301 ( .A(n_134), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g304 ( .A(n_134), .B(n_198), .Y(n_304) );
AND2x2_ASAP7_75t_L g321 ( .A(n_134), .B(n_214), .Y(n_321) );
AND2x2_ASAP7_75t_L g419 ( .A(n_134), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g242 ( .A(n_135), .Y(n_242) );
AND2x4_ASAP7_75t_L g425 ( .A(n_135), .B(n_420), .Y(n_425) );
AO31x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_141), .A3(n_157), .B(n_163), .Y(n_135) );
AO31x2_ASAP7_75t_L g249 ( .A1(n_136), .A2(n_209), .A3(n_250), .B(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_137), .A2(n_588), .B(n_591), .Y(n_587) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_138), .A2(n_187), .A3(n_193), .B(n_194), .Y(n_186) );
AO31x2_ASAP7_75t_L g199 ( .A1(n_138), .A2(n_200), .A3(n_209), .B(n_211), .Y(n_199) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_138), .A2(n_215), .A3(n_222), .B(n_223), .Y(n_214) );
AO31x2_ASAP7_75t_L g623 ( .A1(n_138), .A2(n_165), .A3(n_624), .B(n_627), .Y(n_623) );
BUFx10_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
BUFx10_ASAP7_75t_L g515 ( .A(n_139), .Y(n_515) );
INVx1_ASAP7_75t_L g539 ( .A(n_139), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_148), .B1(n_151), .B2(n_154), .Y(n_141) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_144), .Y(n_583) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g147 ( .A(n_145), .Y(n_147) );
INVx3_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_145), .Y(n_179) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
INVx1_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
INVx1_ASAP7_75t_L g218 ( .A(n_145), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_145), .Y(n_221) );
INVx2_ASAP7_75t_L g231 ( .A(n_145), .Y(n_231) );
INVx1_ASAP7_75t_L g233 ( .A(n_145), .Y(n_233) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_147), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_148), .A2(n_177), .B(n_180), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_148), .A2(n_154), .B1(n_188), .B2(n_190), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_148), .A2(n_201), .B1(n_206), .B2(n_207), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_148), .A2(n_154), .B1(n_216), .B2(n_219), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_148), .A2(n_229), .B1(n_232), .B2(n_234), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_148), .A2(n_207), .B1(n_251), .B2(n_252), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_148), .A2(n_154), .B1(n_270), .B2(n_271), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_148), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_148), .A2(n_234), .B1(n_520), .B2(n_521), .Y(n_519) );
OAI22x1_ASAP7_75t_L g624 ( .A1(n_148), .A2(n_234), .B1(n_625), .B2(n_626), .Y(n_624) );
INVx6_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
O2A1O1Ixp5_ASAP7_75t_L g172 ( .A1(n_149), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_149), .A2(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_149), .B(n_582), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_149), .A2(n_578), .B(n_582), .C(n_585), .Y(n_639) );
BUFx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
INVx1_ASAP7_75t_L g535 ( .A(n_150), .Y(n_535) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx1_ASAP7_75t_L g205 ( .A(n_153), .Y(n_205) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g514 ( .A(n_155), .Y(n_514) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g568 ( .A(n_156), .Y(n_568) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_157), .A2(n_235), .A3(n_269), .B(n_272), .Y(n_268) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_157), .A2(n_587), .B(n_595), .Y(n_586) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_159), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_159), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g165 ( .A(n_160), .Y(n_165) );
INVx2_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
OAI21xp33_ASAP7_75t_L g585 ( .A1(n_160), .A2(n_539), .B(n_580), .Y(n_585) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_161), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_165), .B(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g430 ( .A(n_166), .B(n_331), .Y(n_430) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g259 ( .A(n_167), .Y(n_259) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_167), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_185), .Y(n_167) );
AND2x2_ASAP7_75t_L g247 ( .A(n_168), .B(n_186), .Y(n_247) );
INVx1_ASAP7_75t_L g288 ( .A(n_168), .Y(n_288) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_183), .Y(n_168) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_169), .A2(n_171), .B(n_183), .Y(n_283) );
INVx2_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_170), .B(n_195), .Y(n_194) );
BUFx3_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_170), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_170), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g552 ( .A(n_170), .B(n_515), .Y(n_552) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_176), .B(n_181), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_174), .A2(n_565), .B(n_566), .C(n_567), .Y(n_564) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g191 ( .A(n_179), .Y(n_191) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_179), .A2(n_221), .B1(n_593), .B2(n_594), .Y(n_592) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_SL g235 ( .A(n_182), .Y(n_235) );
INVx2_ASAP7_75t_L g193 ( .A(n_184), .Y(n_193) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_184), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g279 ( .A(n_185), .Y(n_279) );
AND2x2_ASAP7_75t_L g343 ( .A(n_185), .B(n_282), .Y(n_343) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g297 ( .A(n_186), .Y(n_297) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_186), .Y(n_350) );
OR2x2_ASAP7_75t_L g421 ( .A(n_186), .B(n_227), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_189), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g522 ( .A(n_192), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_192), .B(n_547), .Y(n_546) );
AO31x2_ASAP7_75t_L g510 ( .A1(n_193), .A2(n_511), .A3(n_515), .B(n_516), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g299 ( .A(n_196), .B(n_300), .C(n_303), .D(n_305), .Y(n_299) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g437 ( .A(n_197), .B(n_425), .Y(n_437) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_213), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_198), .B(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g291 ( .A(n_198), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_198), .Y(n_311) );
INVx1_ASAP7_75t_L g328 ( .A(n_198), .Y(n_328) );
INVx1_ASAP7_75t_L g336 ( .A(n_198), .Y(n_336) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_198), .Y(n_450) );
INVx4_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_199), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g368 ( .A(n_199), .B(n_268), .Y(n_368) );
AND2x2_ASAP7_75t_L g376 ( .A(n_199), .B(n_214), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_199), .B(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g441 ( .A(n_199), .Y(n_441) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_204), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g234 ( .A(n_208), .Y(n_234) );
AO31x2_ASAP7_75t_L g518 ( .A1(n_209), .A2(n_235), .A3(n_519), .B(n_523), .Y(n_518) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_209), .A2(n_528), .B(n_540), .Y(n_527) );
BUFx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_210), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_210), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g596 ( .A(n_210), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_210), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g245 ( .A(n_214), .Y(n_245) );
OR2x2_ASAP7_75t_L g306 ( .A(n_214), .B(n_268), .Y(n_306) );
INVx2_ASAP7_75t_L g313 ( .A(n_214), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_214), .B(n_266), .Y(n_337) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_214), .Y(n_424) );
OAI21xp33_ASAP7_75t_SL g544 ( .A1(n_217), .A2(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AO31x2_ASAP7_75t_L g227 ( .A1(n_222), .A2(n_228), .A3(n_235), .B(n_236), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_225), .B(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g248 ( .A(n_227), .B(n_249), .Y(n_248) );
BUFx2_ASAP7_75t_L g258 ( .A(n_227), .Y(n_258) );
INVx2_ASAP7_75t_L g276 ( .A(n_227), .Y(n_276) );
AND2x4_ASAP7_75t_L g308 ( .A(n_227), .B(n_280), .Y(n_308) );
OR2x2_ASAP7_75t_L g388 ( .A(n_227), .B(n_288), .Y(n_388) );
INVx2_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_231), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_234), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_243), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_240), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g305 ( .A(n_240), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_240), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_241), .B(n_311), .Y(n_319) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g264 ( .A(n_242), .Y(n_264) );
OR2x2_ASAP7_75t_L g357 ( .A(n_242), .B(n_267), .Y(n_357) );
INVx1_ASAP7_75t_L g284 ( .A(n_243), .Y(n_284) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g256 ( .A(n_244), .Y(n_256) );
INVx1_ASAP7_75t_L g292 ( .A(n_245), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
OAI322xp33_ASAP7_75t_L g260 ( .A1(n_247), .A2(n_261), .A3(n_274), .B1(n_277), .B2(n_284), .C1(n_285), .C2(n_289), .Y(n_260) );
AND2x4_ASAP7_75t_L g307 ( .A(n_247), .B(n_308), .Y(n_307) );
AOI211xp5_ASAP7_75t_SL g338 ( .A1(n_247), .A2(n_339), .B(n_340), .C(n_344), .Y(n_338) );
AND2x2_ASAP7_75t_L g358 ( .A(n_247), .B(n_248), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_247), .B(n_275), .Y(n_364) );
AND2x4_ASAP7_75t_SL g286 ( .A(n_248), .B(n_287), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_248), .B(n_304), .C(n_332), .Y(n_377) );
AND2x2_ASAP7_75t_L g408 ( .A(n_248), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g275 ( .A(n_249), .B(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g280 ( .A(n_249), .Y(n_280) );
BUFx2_ASAP7_75t_L g348 ( .A(n_249), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_258), .B(n_282), .Y(n_281) );
NAND2x1_ASAP7_75t_L g322 ( .A(n_258), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g341 ( .A(n_258), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_259), .B(n_275), .Y(n_406) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g349 ( .A(n_264), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_268), .Y(n_302) );
AND2x4_ASAP7_75t_L g312 ( .A(n_268), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g399 ( .A(n_268), .Y(n_399) );
INVx2_ASAP7_75t_L g420 ( .A(n_268), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g432 ( .A1(n_274), .A2(n_433), .B1(n_435), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g344 ( .A(n_275), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g298 ( .A(n_276), .B(n_282), .Y(n_298) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g317 ( .A(n_278), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x4_ASAP7_75t_L g287 ( .A(n_279), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g409 ( .A(n_279), .Y(n_409) );
INVx2_ASAP7_75t_L g295 ( .A(n_280), .Y(n_295) );
AND2x2_ASAP7_75t_L g323 ( .A(n_280), .B(n_282), .Y(n_323) );
INVx3_ASAP7_75t_L g331 ( .A(n_280), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_280), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
OAI222xp33_ASAP7_75t_L g455 ( .A1(n_285), .A2(n_445), .B1(n_456), .B2(n_459), .C1(n_461), .C2(n_463), .Y(n_455) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g396 ( .A(n_287), .Y(n_396) );
AND2x2_ASAP7_75t_L g460 ( .A(n_287), .B(n_330), .Y(n_460) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_290), .B(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_299), .B1(n_307), .B2(n_309), .C(n_314), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g382 ( .A(n_295), .Y(n_382) );
INVx2_ASAP7_75t_L g444 ( .A(n_296), .Y(n_444) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
AND2x2_ASAP7_75t_L g381 ( .A(n_297), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g347 ( .A(n_298), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g373 ( .A(n_298), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g462 ( .A(n_298), .Y(n_462) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g411 ( .A(n_302), .Y(n_411) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g434 ( .A(n_304), .B(n_312), .Y(n_434) );
AND2x2_ASAP7_75t_L g457 ( .A(n_304), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g318 ( .A(n_306), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g453 ( .A(n_306), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_307), .A2(n_361), .B1(n_395), .B2(n_397), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_307), .A2(n_423), .B(n_426), .Y(n_422) );
INVxp67_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
INVx2_ASAP7_75t_SL g443 ( .A(n_308), .Y(n_443) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
OR2x2_ASAP7_75t_L g356 ( .A(n_310), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g454 ( .A(n_310), .B(n_453), .Y(n_454) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g327 ( .A(n_312), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_312), .B(n_336), .Y(n_352) );
INVx2_ASAP7_75t_L g379 ( .A(n_312), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B1(n_320), .B2(n_322), .Y(n_314) );
NOR2xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_316), .A2(n_390), .B1(n_403), .B2(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g412 ( .A(n_321), .B(n_413), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_329), .B(n_333), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g393 ( .A(n_326), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_326), .B(n_376), .Y(n_404) );
INVx1_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_330), .B(n_343), .Y(n_435) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI21xp33_ASAP7_75t_L g448 ( .A1(n_331), .A2(n_449), .B(n_451), .Y(n_448) );
OAI21xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_338), .B(n_346), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g392 ( .A(n_337), .Y(n_392) );
INVx1_ASAP7_75t_L g458 ( .A(n_337), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g431 ( .A(n_341), .Y(n_431) );
OR2x2_ASAP7_75t_L g442 ( .A(n_342), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .C(n_351), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_347), .A2(n_408), .B1(n_410), .B2(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_349), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_352), .B(n_356), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_352), .A2(n_415), .B1(n_418), .B2(n_421), .C(n_422), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_358), .B(n_359), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g363 ( .A(n_357), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .B1(n_365), .B2(n_845), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g446 ( .A(n_368), .B(n_424), .Y(n_446) );
NAND4xp25_ASAP7_75t_L g369 ( .A(n_370), .B(n_400), .C(n_427), .D(n_447), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_383), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B1(n_377), .B2(n_378), .C(n_380), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_373), .A2(n_430), .B1(n_452), .B2(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g426 ( .A(n_375), .Y(n_426) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g410 ( .A(n_376), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_376), .B(n_419), .Y(n_418) );
NAND2x1_ASAP7_75t_L g463 ( .A(n_376), .B(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_378), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g385 ( .A(n_382), .B(n_386), .Y(n_385) );
OAI21xp33_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_389), .B(n_394), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g413 ( .A(n_399), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_399), .A2(n_428), .B(n_432), .C(n_438), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_414), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_402), .B(n_407), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g461 ( .A(n_409), .B(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx3_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI22xp33_ASAP7_75t_R g438 ( .A1(n_439), .A2(n_442), .B1(n_444), .B2(n_445), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g452 ( .A(n_441), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_455), .Y(n_447) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx5_ASAP7_75t_L g475 ( .A(n_468), .Y(n_475) );
INVx5_ASAP7_75t_L g480 ( .A(n_468), .Y(n_480) );
AND2x6_ASAP7_75t_SL g468 ( .A(n_469), .B(n_471), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_471), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR2x1_ASAP7_75t_L g840 ( .A(n_472), .B(n_494), .Y(n_840) );
BUFx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
NOR2xp67_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
BUFx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx8_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g491 ( .A(n_485), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_485), .B(n_838), .Y(n_837) );
OAI321xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_495), .A3(n_826), .B1(n_831), .B2(n_832), .C(n_833), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_488), .B(n_826), .Y(n_832) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx6_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x6_ASAP7_75t_SL g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g831 ( .A(n_495), .Y(n_831) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_499), .Y(n_502) );
BUFx8_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g839 ( .A(n_500), .B(n_840), .Y(n_839) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_718), .Y(n_503) );
NOR2xp67_ASAP7_75t_L g504 ( .A(n_505), .B(n_660), .Y(n_504) );
NAND3xp33_ASAP7_75t_SL g505 ( .A(n_506), .B(n_597), .C(n_642), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_553), .B(n_574), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_507), .A2(n_598), .B1(n_617), .B2(n_629), .Y(n_597) );
AOI22x1_ASAP7_75t_L g722 ( .A1(n_507), .A2(n_723), .B1(n_727), .B2(n_728), .Y(n_722) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_525), .Y(n_508) );
OR2x2_ASAP7_75t_L g683 ( .A(n_509), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_518), .Y(n_509) );
OR2x2_ASAP7_75t_L g558 ( .A(n_510), .B(n_518), .Y(n_558) );
AND2x2_ASAP7_75t_L g601 ( .A(n_510), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g609 ( .A(n_510), .Y(n_609) );
BUFx2_ASAP7_75t_L g659 ( .A(n_510), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_514), .A2(n_550), .B(n_551), .Y(n_549) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_514), .A2(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g573 ( .A(n_515), .Y(n_573) );
AND2x2_ASAP7_75t_L g604 ( .A(n_518), .B(n_541), .Y(n_604) );
INVx1_ASAP7_75t_L g611 ( .A(n_518), .Y(n_611) );
INVx1_ASAP7_75t_L g616 ( .A(n_518), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_518), .B(n_609), .Y(n_678) );
INVx1_ASAP7_75t_L g699 ( .A(n_518), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_518), .B(n_602), .Y(n_769) );
INVx1_ASAP7_75t_L g662 ( .A(n_525), .Y(n_662) );
OR2x2_ASAP7_75t_L g714 ( .A(n_525), .B(n_678), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_541), .Y(n_525) );
AND2x2_ASAP7_75t_L g559 ( .A(n_526), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g607 ( .A(n_526), .B(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g613 ( .A(n_526), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_526), .B(n_556), .Y(n_690) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g602 ( .A(n_527), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_536), .B(n_539), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_532), .B(n_534), .Y(n_529) );
BUFx4f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_535), .B(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g556 ( .A(n_541), .Y(n_556) );
INVx1_ASAP7_75t_L g656 ( .A(n_541), .Y(n_656) );
AND2x2_ASAP7_75t_L g658 ( .A(n_541), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g676 ( .A(n_541), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g698 ( .A(n_541), .B(n_699), .Y(n_698) );
NAND2x1p5_ASAP7_75t_SL g709 ( .A(n_541), .B(n_685), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_541), .B(n_616), .Y(n_799) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_549), .B(n_552), .Y(n_543) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_554), .A2(n_738), .B1(n_739), .B2(n_741), .Y(n_737) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_555), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_555), .B(n_794), .Y(n_793) );
OR2x2_ASAP7_75t_L g816 ( .A(n_555), .B(n_674), .Y(n_816) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g615 ( .A(n_556), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_556), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g704 ( .A(n_556), .B(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g655 ( .A(n_557), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g745 ( .A(n_558), .Y(n_745) );
OR2x2_ASAP7_75t_L g819 ( .A(n_558), .B(n_746), .Y(n_819) );
INVx1_ASAP7_75t_L g650 ( .A(n_559), .Y(n_650) );
INVx3_ASAP7_75t_L g654 ( .A(n_560), .Y(n_654) );
BUFx2_ASAP7_75t_L g665 ( .A(n_560), .Y(n_665) );
BUFx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g635 ( .A(n_561), .B(n_586), .Y(n_635) );
INVx2_ASAP7_75t_L g681 ( .A(n_561), .Y(n_681) );
INVx1_ASAP7_75t_L g713 ( .A(n_561), .Y(n_713) );
AND2x2_ASAP7_75t_L g726 ( .A(n_561), .B(n_623), .Y(n_726) );
AND2x2_ASAP7_75t_L g748 ( .A(n_561), .B(n_647), .Y(n_748) );
NAND2x1p5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_569), .B(n_572), .Y(n_563) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g739 ( .A(n_575), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_575), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g764 ( .A(n_575), .B(n_632), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_575), .B(n_766), .Y(n_765) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_586), .Y(n_575) );
INVx2_ASAP7_75t_L g621 ( .A(n_576), .Y(n_621) );
AND2x2_ASAP7_75t_L g648 ( .A(n_576), .B(n_649), .Y(n_648) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B(n_584), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g622 ( .A(n_586), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g641 ( .A(n_586), .Y(n_641) );
INVx2_ASAP7_75t_L g649 ( .A(n_586), .Y(n_649) );
OR2x2_ASAP7_75t_L g669 ( .A(n_586), .B(n_623), .Y(n_669) );
AND2x2_ASAP7_75t_L g680 ( .A(n_586), .B(n_681), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_603), .B1(n_605), .B2(n_610), .C(n_612), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI32xp33_ASAP7_75t_L g710 ( .A1(n_600), .A2(n_614), .A3(n_711), .B1(n_714), .B2(n_715), .Y(n_710) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g700 ( .A(n_601), .Y(n_700) );
AND2x2_ASAP7_75t_L g736 ( .A(n_601), .B(n_615), .Y(n_736) );
INVx1_ASAP7_75t_L g800 ( .A(n_601), .Y(n_800) );
OR2x2_ASAP7_75t_L g674 ( .A(n_602), .B(n_609), .Y(n_674) );
INVx2_ASAP7_75t_L g685 ( .A(n_602), .Y(n_685) );
BUFx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g824 ( .A(n_604), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_L g811 ( .A(n_607), .Y(n_811) );
INVx1_ASAP7_75t_L g825 ( .A(n_607), .Y(n_825) );
OR2x2_ASAP7_75t_L g705 ( .A(n_608), .B(n_685), .Y(n_705) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_610), .B(n_705), .Y(n_727) );
INVx1_ASAP7_75t_L g758 ( .A(n_610), .Y(n_758) );
BUFx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g792 ( .A(n_611), .Y(n_792) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2x1_ASAP7_75t_L g761 ( .A(n_613), .B(n_762), .Y(n_761) );
OAI21xp5_ASAP7_75t_SL g783 ( .A1(n_614), .A2(n_784), .B(n_789), .Y(n_783) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
AND2x2_ASAP7_75t_L g693 ( .A(n_619), .B(n_635), .Y(n_693) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_619), .Y(n_823) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g725 ( .A(n_620), .Y(n_725) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g707 ( .A(n_621), .B(n_681), .Y(n_707) );
AND2x2_ASAP7_75t_L g778 ( .A(n_621), .B(n_649), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_622), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g706 ( .A(n_622), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g785 ( .A(n_622), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g634 ( .A(n_623), .Y(n_634) );
INVx2_ASAP7_75t_L g647 ( .A(n_623), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_623), .B(n_638), .Y(n_695) );
AND2x2_ASAP7_75t_L g755 ( .A(n_623), .B(n_649), .Y(n_755) );
NAND2xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_636), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g730 ( .A(n_633), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_633), .B(n_713), .Y(n_805) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g637 ( .A(n_634), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g766 ( .A(n_634), .B(n_681), .Y(n_766) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_640), .Y(n_636) );
OR2x2_ASAP7_75t_L g711 ( .A(n_637), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g668 ( .A(n_638), .Y(n_668) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g694 ( .A(n_641), .B(n_695), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_655), .B1(n_657), .B2(n_658), .Y(n_642) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_650), .B(n_651), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g657 ( .A(n_645), .B(n_654), .Y(n_657) );
BUFx2_ASAP7_75t_L g675 ( .A(n_645), .Y(n_675) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g686 ( .A(n_646), .Y(n_686) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g701 ( .A(n_648), .B(n_665), .Y(n_701) );
INVx2_ASAP7_75t_L g717 ( .A(n_648), .Y(n_717) );
AND2x2_ASAP7_75t_L g759 ( .A(n_648), .B(n_681), .Y(n_759) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g734 ( .A(n_654), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g781 ( .A(n_655), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g812 ( .A(n_656), .Y(n_812) );
INVx2_ASAP7_75t_L g751 ( .A(n_659), .Y(n_751) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_670), .C(n_687), .D(n_702), .Y(n_660) );
NAND2xp33_ASAP7_75t_SL g661 ( .A(n_662), .B(n_663), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_663), .A2(n_741), .B1(n_757), .B2(n_759), .C(n_760), .Y(n_756) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g738 ( .A(n_667), .Y(n_738) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx2_ASAP7_75t_L g731 ( .A(n_668), .Y(n_731) );
INVx2_ASAP7_75t_L g803 ( .A(n_669), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B1(n_676), .B2(n_679), .C1(n_682), .C2(n_686), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g757 ( .A(n_673), .B(n_758), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_673), .A2(n_785), .B(n_787), .Y(n_784) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g796 ( .A(n_674), .B(n_740), .Y(n_796) );
OAI21xp33_ASAP7_75t_SL g770 ( .A1(n_675), .A2(n_696), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g689 ( .A(n_678), .B(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_SL g741 ( .A(n_678), .Y(n_741) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g740 ( .A(n_681), .Y(n_740) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g746 ( .A(n_685), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_691), .B1(n_696), .B2(n_701), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_693), .A2(n_703), .B1(n_706), .B2(n_708), .C(n_710), .Y(n_702) );
INVx3_ASAP7_75t_R g817 ( .A(n_694), .Y(n_817) );
INVx1_ASAP7_75t_L g735 ( .A(n_695), .Y(n_735) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_698), .Y(n_752) );
INVx1_ASAP7_75t_L g762 ( .A(n_698), .Y(n_762) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_707), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g780 ( .A(n_707), .Y(n_780) );
AND2x2_ASAP7_75t_L g808 ( .A(n_707), .B(n_755), .Y(n_808) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g802 ( .A(n_712), .B(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_774), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_756), .C(n_770), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_732), .C(n_742), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI21xp33_ASAP7_75t_L g733 ( .A1(n_723), .A2(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g773 ( .A(n_725), .Y(n_773) );
AND2x2_ASAP7_75t_L g814 ( .A(n_725), .B(n_803), .Y(n_814) );
NAND2x1_ASAP7_75t_L g772 ( .A(n_726), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g794 ( .A(n_731), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_737), .Y(n_732) );
INVx1_ASAP7_75t_L g786 ( .A(n_740), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_747), .B1(n_749), .B2(n_753), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g782 ( .A(n_746), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_748), .B(n_778), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g821 ( .A(n_754), .Y(n_821) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI22xp33_ASAP7_75t_SL g760 ( .A1(n_761), .A2(n_763), .B1(n_765), .B2(n_767), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_801), .Y(n_774) );
O2A1O1Ixp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_779), .B(n_781), .C(n_783), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OAI21xp33_ASAP7_75t_L g790 ( .A1(n_777), .A2(n_791), .B(n_793), .Y(n_790) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
O2A1O1Ixp5_ASAP7_75t_SL g801 ( .A1(n_781), .A2(n_802), .B(n_804), .C(n_806), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_785), .A2(n_790), .B1(n_795), .B2(n_797), .Y(n_789) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OR2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI211xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_809), .B(n_813), .C(n_820), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_813) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI21xp5_ASAP7_75t_SL g820 ( .A1(n_821), .A2(n_822), .B(n_824), .Y(n_820) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
BUFx10_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_R g841 ( .A(n_842), .B(n_843), .Y(n_841) );
endmodule