module fake_netlist_1_235_n_702 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_702);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_702;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_40), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_44), .Y(n_81) );
BUFx6f_ASAP7_75t_L g82 ( .A(n_18), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_65), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_34), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_46), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_28), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx4_ASAP7_75t_R g89 ( .A(n_27), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_36), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_72), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_9), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_59), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_32), .Y(n_94) );
BUFx10_ASAP7_75t_L g95 ( .A(n_49), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_17), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_0), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_73), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_48), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_54), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_67), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_55), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_4), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_68), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_77), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_62), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_19), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_1), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_31), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_45), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_13), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_42), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g116 ( .A(n_53), .B(n_10), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_78), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_23), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_66), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_76), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_56), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_70), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_22), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_64), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_12), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_52), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_29), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_24), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_113), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_113), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_125), .B(n_90), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_125), .B(n_2), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_122), .A2(n_96), .B1(n_110), .B2(n_88), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_97), .B(n_4), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_115), .B(n_5), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_110), .B(n_5), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_106), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
AOI22x1_ASAP7_75t_SL g147 ( .A1(n_103), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_98), .B(n_38), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_91), .B(n_10), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_108), .B(n_11), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_95), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_100), .B(n_11), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_98), .B(n_12), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_95), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g157 ( .A1(n_101), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_101), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_102), .A2(n_17), .B1(n_20), .B2(n_21), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_80), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_80), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_102), .A2(n_25), .B1(n_26), .B2(n_30), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_99), .B(n_33), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_105), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_105), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_127), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_107), .B(n_79), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_107), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_81), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
INVx4_ASAP7_75t_SL g174 ( .A(n_148), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_156), .B(n_112), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_151), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_131), .A2(n_118), .B1(n_117), .B2(n_111), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_156), .B(n_114), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_152), .B(n_118), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_170), .B(n_114), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_129), .A2(n_116), .B1(n_117), .B2(n_111), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_132), .B(n_104), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_159), .A2(n_127), .B1(n_126), .B2(n_83), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_153), .B(n_126), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_152), .B(n_104), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_152), .B(n_123), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_130), .B(n_93), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_134), .Y(n_197) );
BUFx10_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_136), .A2(n_81), .B1(n_83), .B2(n_84), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_156), .B(n_124), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_162), .B(n_121), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_170), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_153), .B(n_94), .Y(n_207) );
AND2x6_ASAP7_75t_L g208 ( .A(n_139), .B(n_94), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
INVx4_ASAP7_75t_SL g211 ( .A(n_148), .Y(n_211) );
XOR2xp5_ASAP7_75t_L g212 ( .A(n_147), .B(n_93), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_163), .B(n_120), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_167), .B(n_109), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_169), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_134), .Y(n_219) );
INVx4_ASAP7_75t_SL g220 ( .A(n_138), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_133), .B(n_85), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g223 ( .A1(n_157), .A2(n_160), .B1(n_143), .B2(n_161), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_172), .B(n_119), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_158), .Y(n_225) );
NAND2xp33_ASAP7_75t_L g226 ( .A(n_149), .B(n_87), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_166), .A2(n_171), .B1(n_168), .B2(n_145), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_144), .B(n_85), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_150), .B(n_84), .Y(n_229) );
INVx6_ASAP7_75t_L g230 ( .A(n_138), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_166), .B(n_87), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_168), .B(n_171), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_140), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_140), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_165), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_165), .B(n_87), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_188), .B(n_164), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_223), .B(n_147), .C(n_89), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_188), .B(n_87), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_231), .Y(n_240) );
INVxp67_ASAP7_75t_SL g241 ( .A(n_192), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_180), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_233), .B(n_234), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_217), .B(n_87), .Y(n_245) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_191), .A2(n_82), .B(n_142), .C(n_138), .Y(n_246) );
AND2x6_ASAP7_75t_SL g247 ( .A(n_221), .B(n_82), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_232), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_202), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_189), .B(n_142), .Y(n_250) );
AND2x6_ASAP7_75t_SL g251 ( .A(n_221), .B(n_142), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_191), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_208), .A2(n_142), .B1(n_138), .B2(n_39), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_198), .B(n_35), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_209), .B(n_37), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_192), .Y(n_257) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_186), .B(n_41), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_181), .B(n_43), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_186), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_215), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_222), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_208), .A2(n_47), .B1(n_50), .B2(n_51), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_193), .B(n_57), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
NOR2x2_ASAP7_75t_L g266 ( .A(n_221), .B(n_75), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_228), .B(n_58), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_SL g268 ( .A1(n_176), .A2(n_61), .B(n_63), .C(n_69), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_208), .A2(n_71), .B1(n_74), .B2(n_204), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_198), .B(n_218), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_228), .B(n_176), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_194), .B(n_207), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_182), .A2(n_179), .B(n_236), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_178), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_201), .B(n_174), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_207), .B(n_208), .Y(n_277) );
NAND3xp33_ASAP7_75t_SL g278 ( .A(n_212), .B(n_199), .C(n_190), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_177), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_185), .A2(n_196), .B1(n_177), .B2(n_175), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_235), .B(n_200), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_201), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_195), .B(n_183), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_205), .B(n_206), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_225), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_179), .B(n_190), .Y(n_286) );
OAI22xp5_ASAP7_75t_SL g287 ( .A1(n_223), .A2(n_187), .B1(n_227), .B2(n_203), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_210), .B(n_174), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_203), .B(n_214), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_184), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_173), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_226), .B(n_227), .C(n_182), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_174), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_229), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_216), .B(n_224), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_211), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_173), .Y(n_297) );
AO22x1_ASAP7_75t_L g298 ( .A1(n_211), .A2(n_187), .B1(n_226), .B2(n_213), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_211), .B(n_220), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_220), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_230), .A2(n_197), .B1(n_213), .B2(n_219), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_220), .B(n_197), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_219), .Y(n_304) );
O2A1O1Ixp5_ASAP7_75t_L g305 ( .A1(n_188), .A2(n_191), .B(n_182), .C(n_233), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_243), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_287), .A2(n_270), .B1(n_241), .B2(n_278), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_252), .B(n_274), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_257), .Y(n_309) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_238), .B(n_274), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_284), .A2(n_295), .B(n_286), .Y(n_311) );
NAND3xp33_ASAP7_75t_SL g312 ( .A(n_275), .B(n_289), .C(n_281), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_294), .B(n_248), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_247), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_248), .B(n_272), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_244), .A2(n_283), .B(n_271), .C(n_273), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_277), .A2(n_280), .B1(n_256), .B2(n_290), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_261), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_256), .B(n_285), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_252), .B(n_282), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_251), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_275), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_237), .B(n_279), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_285), .A2(n_292), .B(n_305), .C(n_261), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_262), .B(n_249), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_262), .B(n_265), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_260), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_250), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_249), .A2(n_240), .B(n_255), .C(n_267), .Y(n_329) );
INVx8_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_293), .B(n_252), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_265), .B(n_242), .Y(n_332) );
BUFx4f_ASAP7_75t_L g333 ( .A(n_258), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_265), .B(n_242), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_240), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_260), .B(n_282), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_269), .A2(n_258), .B1(n_263), .B2(n_264), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_258), .A2(n_259), .B1(n_245), .B2(n_253), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_298), .A2(n_288), .B1(n_239), .B2(n_276), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_298), .B(n_288), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_254), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_301), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_268), .A2(n_246), .B(n_297), .C(n_291), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_266), .B(n_293), .Y(n_344) );
NAND3xp33_ASAP7_75t_SL g345 ( .A(n_266), .B(n_302), .C(n_300), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_293), .A2(n_296), .B1(n_299), .B2(n_300), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_296), .B(n_254), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_291), .A2(n_297), .B(n_303), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_254), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_303), .A2(n_304), .B(n_254), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_284), .B(n_295), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_254), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_304), .A2(n_284), .B(n_295), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_SL g354 ( .A1(n_304), .A2(n_264), .B(n_259), .C(n_268), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_304), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_261), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_SL g357 ( .A1(n_255), .A2(n_244), .B(n_179), .C(n_283), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_270), .B(n_243), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_295), .B(n_294), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_357), .A2(n_359), .B(n_316), .C(n_313), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_315), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_306), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_312), .B(n_358), .Y(n_364) );
BUFx2_ASAP7_75t_SL g365 ( .A(n_314), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_343), .A2(n_338), .B(n_337), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_351), .A2(n_353), .B(n_311), .Y(n_367) );
OAI22x1_ASAP7_75t_SL g368 ( .A1(n_322), .A2(n_310), .B1(n_321), .B2(n_309), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_SL g369 ( .A1(n_329), .A2(n_324), .B(n_345), .C(n_351), .Y(n_369) );
CKINVDCx11_ASAP7_75t_R g370 ( .A(n_330), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_307), .B(n_344), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_317), .A2(n_319), .B1(n_328), .B2(n_311), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_325), .B(n_354), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_316), .B(n_323), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_343), .A2(n_348), .B(n_350), .Y(n_375) );
AO31x2_ASAP7_75t_L g376 ( .A1(n_340), .A2(n_348), .A3(n_318), .B(n_356), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_SL g377 ( .A1(n_346), .A2(n_336), .B(n_355), .C(n_347), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_333), .B(n_327), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_334), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_330), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_SL g384 ( .A1(n_320), .A2(n_339), .B(n_350), .C(n_333), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_332), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_331), .A2(n_308), .B(n_352), .C(n_327), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_349), .B(n_330), .Y(n_387) );
BUFx2_ASAP7_75t_R g388 ( .A(n_341), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_327), .A2(n_311), .B(n_316), .C(n_313), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_311), .A2(n_359), .B(n_191), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_359), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_359), .B(n_270), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g393 ( .A1(n_311), .A2(n_316), .B(n_313), .C(n_351), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_364), .A2(n_391), .B1(n_371), .B2(n_365), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_361), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_391), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g397 ( .A1(n_360), .A2(n_374), .B(n_362), .C(n_393), .Y(n_397) );
AO21x2_ASAP7_75t_L g398 ( .A1(n_367), .A2(n_366), .B(n_373), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_366), .A2(n_389), .B(n_393), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_392), .A2(n_363), .B1(n_378), .B2(n_382), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_381), .B(n_361), .Y(n_401) );
AO31x2_ASAP7_75t_L g402 ( .A1(n_389), .A2(n_386), .A3(n_390), .B(n_369), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_382), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_385), .B(n_379), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_386), .B(n_380), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_369), .B(n_384), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_376), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_377), .A2(n_384), .B(n_375), .Y(n_408) );
OA21x2_ASAP7_75t_L g409 ( .A1(n_376), .A2(n_377), .B(n_387), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_376), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_368), .A2(n_382), .B1(n_383), .B2(n_370), .C(n_376), .Y(n_411) );
INVx4_ASAP7_75t_L g412 ( .A(n_370), .Y(n_412) );
AO21x2_ASAP7_75t_L g413 ( .A1(n_388), .A2(n_367), .B(n_366), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_391), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_361), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_391), .B(n_362), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_364), .B(n_312), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_362), .B1(n_313), .B2(n_307), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_366), .A2(n_367), .B(n_375), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_361), .Y(n_421) );
BUFx2_ASAP7_75t_R g422 ( .A(n_365), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_397), .B(n_418), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_419), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_421), .B(n_407), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_407), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_414), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_395), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_395), .B(n_415), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_421), .B(n_410), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_406), .A2(n_408), .B(n_410), .Y(n_431) );
OR2x6_ASAP7_75t_L g432 ( .A(n_406), .B(n_419), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_415), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_417), .A2(n_405), .B(n_416), .Y(n_434) );
AO21x1_ASAP7_75t_L g435 ( .A1(n_421), .A2(n_401), .B(n_404), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_409), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_416), .B(n_401), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_399), .A2(n_398), .B(n_413), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_414), .B(n_396), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_414), .B(n_396), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_411), .A2(n_399), .B(n_398), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_399), .B(n_409), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_399), .A2(n_398), .B(n_420), .Y(n_446) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_398), .A2(n_413), .B(n_420), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_420), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_394), .B(n_400), .Y(n_449) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_413), .A2(n_420), .B(n_402), .Y(n_450) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_413), .A2(n_402), .B(n_419), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_402), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_402), .B(n_403), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_403), .A2(n_402), .B(n_412), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_402), .B(n_403), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_426), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_425), .B(n_412), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
AOI33xp33_ASAP7_75t_L g461 ( .A1(n_438), .A2(n_412), .A3(n_422), .B1(n_445), .B2(n_455), .B3(n_433), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_425), .B(n_412), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_425), .B(n_430), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_425), .B(n_430), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_448), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_428), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_430), .B(n_437), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_430), .B(n_437), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_427), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_445), .B(n_455), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_448), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_427), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_433), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_445), .B(n_455), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_424), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_435), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_438), .B(n_441), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_441), .B(n_442), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_455), .B(n_452), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_455), .B(n_452), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_435), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_453), .B(n_446), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_435), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_427), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_453), .B(n_446), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_423), .A2(n_449), .B1(n_442), .B2(n_434), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_453), .B(n_446), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_446), .B(n_444), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_454), .B(n_432), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_446), .B(n_444), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_446), .B(n_444), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_444), .B(n_439), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_429), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_427), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_432), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_444), .B(n_439), .Y(n_498) );
AND2x4_ASAP7_75t_SL g499 ( .A(n_432), .B(n_449), .Y(n_499) );
NOR2x1p5_ASAP7_75t_L g500 ( .A(n_473), .B(n_423), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_471), .B(n_444), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_467), .B(n_454), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_481), .B(n_432), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_495), .B(n_434), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_460), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_471), .B(n_439), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_471), .B(n_439), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_476), .B(n_439), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_488), .A2(n_436), .B1(n_440), .B2(n_443), .C(n_450), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_476), .B(n_450), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_466), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_476), .B(n_450), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_466), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_469), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_473), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_463), .B(n_450), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_457), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_467), .B(n_450), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_463), .B(n_447), .Y(n_520) );
BUFx2_ASAP7_75t_L g521 ( .A(n_469), .Y(n_521) );
INVx5_ASAP7_75t_L g522 ( .A(n_470), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_457), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_474), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_463), .B(n_447), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_473), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_464), .B(n_447), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_468), .B(n_480), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_468), .B(n_447), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_480), .B(n_447), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_464), .B(n_451), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_464), .B(n_451), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_457), .B(n_462), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_481), .B(n_451), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_479), .B(n_451), .Y(n_536) );
INVx4_ASAP7_75t_L g537 ( .A(n_462), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_481), .B(n_451), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_462), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_482), .B(n_431), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_475), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_474), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_472), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_472), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_479), .B(n_431), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_458), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_458), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_482), .B(n_431), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_459), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_477), .Y(n_551) );
INVxp67_ASAP7_75t_L g552 ( .A(n_470), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_537), .B(n_482), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_508), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_520), .B(n_487), .Y(n_555) );
OAI31xp33_ASAP7_75t_SL g556 ( .A1(n_523), .A2(n_488), .A3(n_456), .B(n_486), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_537), .B(n_491), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_508), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_529), .B(n_489), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_529), .B(n_487), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_504), .A2(n_461), .B(n_485), .Y(n_561) );
NAND2x1_ASAP7_75t_SL g562 ( .A(n_537), .B(n_478), .Y(n_562) );
NAND2x1_ASAP7_75t_L g563 ( .A(n_516), .B(n_491), .Y(n_563) );
NAND2x1_ASAP7_75t_L g564 ( .A(n_516), .B(n_491), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_520), .B(n_487), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_525), .B(n_484), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_524), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_534), .B(n_496), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_524), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_547), .B(n_489), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_522), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_503), .B(n_491), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_531), .B(n_489), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_543), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_525), .B(n_484), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_548), .B(n_484), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_505), .B(n_490), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_512), .B(n_490), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_527), .B(n_490), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_510), .B(n_478), .C(n_483), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_527), .B(n_492), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_516), .Y(n_584) );
OAI21xp33_ASAP7_75t_L g585 ( .A1(n_506), .A2(n_498), .B(n_494), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_511), .B(n_492), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_511), .B(n_492), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_538), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_513), .B(n_493), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_551), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_550), .Y(n_591) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_526), .B(n_499), .Y(n_592) );
OR2x6_ASAP7_75t_L g593 ( .A(n_500), .B(n_526), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_551), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_528), .Y(n_595) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_515), .B(n_499), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_544), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_522), .A2(n_499), .B(n_470), .C(n_496), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_544), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_506), .B(n_493), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_595), .B(n_540), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_560), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_590), .Y(n_605) );
AOI22x1_ASAP7_75t_SL g606 ( .A1(n_556), .A2(n_486), .B1(n_456), .B2(n_542), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_593), .A2(n_518), .B1(n_517), .B2(n_513), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_586), .B(n_509), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_584), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_555), .B(n_539), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_586), .B(n_509), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_597), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_555), .B(n_539), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_590), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_584), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_591), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_571), .B(n_522), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_587), .B(n_507), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_559), .B(n_518), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_587), .B(n_507), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_598), .A2(n_496), .B(n_522), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_589), .B(n_517), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g624 ( .A1(n_585), .A2(n_501), .B1(n_535), .B2(n_541), .C1(n_549), .C2(n_533), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_565), .B(n_535), .Y(n_625) );
NOR2xp67_ASAP7_75t_SL g626 ( .A(n_571), .B(n_522), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_563), .A2(n_552), .B(n_521), .C(n_515), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_565), .B(n_533), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g629 ( .A1(n_598), .A2(n_557), .B(n_553), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_582), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_566), .B(n_532), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_566), .B(n_532), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_554), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_597), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_594), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_553), .A2(n_491), .B1(n_557), .B2(n_503), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_589), .B(n_501), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_558), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_622), .B(n_601), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_603), .B(n_580), .Y(n_641) );
AOI21xp33_ASAP7_75t_SL g642 ( .A1(n_629), .A2(n_593), .B(n_592), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_624), .B(n_581), .C(n_561), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_609), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_615), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_604), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_627), .A2(n_564), .B(n_563), .C(n_562), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_606), .B(n_485), .C(n_483), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_628), .B(n_580), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_627), .A2(n_593), .B(n_574), .C(n_564), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_630), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_616), .B(n_583), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_617), .B(n_592), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_610), .A2(n_576), .A3(n_583), .B1(n_568), .B2(n_557), .C1(n_596), .C2(n_549), .Y(n_654) );
AOI32xp33_ASAP7_75t_L g655 ( .A1(n_619), .A2(n_576), .A3(n_572), .B1(n_521), .B2(n_574), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_633), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_638), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_639), .Y(n_658) );
AOI32xp33_ASAP7_75t_L g659 ( .A1(n_636), .A2(n_572), .A3(n_541), .B1(n_503), .B2(n_570), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_628), .B(n_577), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_610), .B(n_572), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_612), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_617), .A2(n_593), .B(n_596), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_653), .A2(n_621), .B(n_607), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_643), .A2(n_602), .B(n_608), .C(n_620), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_642), .A2(n_663), .B1(n_655), .B2(n_647), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_646), .B(n_631), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_650), .A2(n_626), .B(n_562), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_662), .Y(n_669) );
OAI32xp33_ASAP7_75t_L g670 ( .A1(n_644), .A2(n_606), .A3(n_637), .B1(n_618), .B2(n_611), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_648), .A2(n_502), .B1(n_494), .B2(n_498), .Y(n_671) );
AO21x1_ASAP7_75t_L g672 ( .A1(n_651), .A2(n_612), .B(n_634), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_652), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g674 ( .A1(n_645), .A2(n_626), .B(n_502), .C(n_531), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_652), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_641), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_659), .A2(n_579), .B(n_578), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_666), .B(n_654), .C(n_640), .D(n_641), .Y(n_678) );
AOI311xp33_ASAP7_75t_L g679 ( .A1(n_664), .A2(n_658), .A3(n_657), .B(n_656), .C(n_649), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_671), .A2(n_660), .B(n_623), .C(n_536), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_665), .A2(n_613), .B1(n_625), .B2(n_631), .C(n_632), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_671), .A2(n_536), .B(n_530), .C(n_519), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_665), .A2(n_613), .B1(n_625), .B2(n_632), .C(n_661), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_670), .A2(n_634), .B1(n_573), .B2(n_569), .C(n_575), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_677), .A2(n_635), .B1(n_614), .B2(n_605), .C(n_600), .Y(n_685) );
AND4x1_ASAP7_75t_L g686 ( .A(n_679), .B(n_668), .C(n_674), .D(n_676), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_684), .A2(n_675), .B(n_673), .C(n_667), .Y(n_687) );
AOI211xp5_ASAP7_75t_SL g688 ( .A1(n_680), .A2(n_685), .B(n_682), .C(n_683), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_678), .B(n_669), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_681), .B(n_542), .C(n_635), .Y(n_690) );
OAI21x1_ASAP7_75t_L g691 ( .A1(n_689), .A2(n_672), .B(n_614), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_687), .A2(n_530), .B1(n_519), .B2(n_546), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_686), .B(n_605), .C(n_599), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_693), .B(n_688), .C(n_690), .D(n_546), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_691), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_695), .Y(n_696) );
INVx3_ASAP7_75t_SL g697 ( .A(n_694), .Y(n_697) );
OAI22x1_ASAP7_75t_SL g698 ( .A1(n_696), .A2(n_692), .B1(n_542), .B2(n_475), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_698), .B(n_697), .C(n_494), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g700 ( .A1(n_699), .A2(n_498), .B(n_493), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_700), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_475), .B1(n_497), .B2(n_588), .Y(n_702) );
endmodule