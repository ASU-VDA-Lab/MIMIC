module fake_jpeg_15736_n_113 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_0),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_71),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_44),
.B1(n_38),
.B2(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_52),
.B1(n_55),
.B2(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_1),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_56),
.B(n_41),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_76),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_77),
.B1(n_82),
.B2(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_43),
.B1(n_42),
.B2(n_48),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_16),
.B1(n_33),
.B2(n_32),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_4),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_13),
.B1(n_31),
.B2(n_30),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_79),
.C(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_70),
.A3(n_11),
.B1(n_19),
.B2(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_2),
.C(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_85),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_86),
.B1(n_80),
.B2(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_94),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_99),
.B(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_80),
.B1(n_89),
.B2(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_105),
.C(n_103),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_101),
.B(n_5),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_109)
);

OAI321xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_21),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.C(n_9),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_4),
.C(n_8),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_10),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_10),
.Y(n_113)
);


endmodule