module real_jpeg_25434_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx6_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_0),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_2),
.A2(n_62),
.B1(n_71),
.B2(n_72),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_62),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_71),
.B1(n_72),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_86),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

INVx8_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_7),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_71),
.B1(n_72),
.B2(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_8),
.B(n_42),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_8),
.B(n_67),
.C(n_71),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_28),
.B1(n_55),
.B2(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_8),
.B(n_60),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_87),
.B1(n_91),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_9),
.A2(n_27),
.B1(n_41),
.B2(n_51),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_9),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_9),
.A2(n_51),
.B1(n_71),
.B2(n_72),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_46),
.B1(n_71),
.B2(n_72),
.Y(n_170)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_13),
.A2(n_71),
.B1(n_72),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_15),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_75),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_15),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_20),
.B(n_106),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.C(n_93),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_21),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_49),
.C(n_63),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_28),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_28),
.B(n_70),
.Y(n_176)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_28),
.B(n_36),
.CON(n_185),
.SN(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_29),
.A2(n_33),
.B(n_36),
.C(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_31),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_32),
.A2(n_44),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_38)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_35),
.C(n_41),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_36),
.B1(n_54),
.B2(n_58),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_36),
.B(n_55),
.C(n_58),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_63),
.B2(n_64),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_52),
.A2(n_60),
.B1(n_96),
.B2(n_185),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_54),
.A2(n_56),
.B(n_185),
.C(n_186),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_56),
.B(n_142),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_60),
.B(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_61),
.Y(n_128)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_76),
.Y(n_64)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_65),
.A2(n_70),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_65),
.A2(n_70),
.B1(n_146),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_65),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_72),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_74),
.B(n_79),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_79),
.A2(n_117),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_80),
.B(n_93),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_83),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_89),
.B(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_87),
.A2(n_113),
.B1(n_163),
.B2(n_170),
.Y(n_177)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_88),
.Y(n_103)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_92),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.C(n_101),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_94),
.B(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_103),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_120),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_118),
.B2(n_119),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_112),
.A2(n_157),
.B(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_131),
.B2(n_132),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_131),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_212),
.B(n_216),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_197),
.B(n_211),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_181),
.B(n_196),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_158),
.B(n_180),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_167),
.B(n_179),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_165),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_175),
.B(n_178),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_195),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_195),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_191),
.C(n_194),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_199),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_206),
.C(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);


endmodule