module fake_jpeg_29957_n_351 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_351);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_59),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_30),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_67),
.B(n_71),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_27),
.B1(n_19),
.B2(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_69),
.A2(n_77),
.B1(n_82),
.B2(n_7),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_27),
.B1(n_39),
.B2(n_20),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_92),
.B1(n_104),
.B2(n_55),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_18),
.B(n_41),
.C(n_32),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_85),
.B1(n_89),
.B2(n_23),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_42),
.B1(n_19),
.B2(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_78),
.B(n_2),
.Y(n_133)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_18),
.B1(n_41),
.B2(n_20),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_80),
.A2(n_83),
.B1(n_106),
.B2(n_8),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_42),
.B1(n_40),
.B2(n_28),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_37),
.B1(n_24),
.B2(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_39),
.B1(n_26),
.B2(n_29),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_37),
.B1(n_26),
.B2(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_29),
.B1(n_36),
.B2(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_48),
.B(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_42),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_109),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_49),
.A2(n_21),
.B1(n_40),
.B2(n_28),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_21),
.B1(n_33),
.B2(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_35),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_64),
.B1(n_35),
.B2(n_33),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_111),
.A2(n_110),
.B1(n_12),
.B2(n_13),
.Y(n_179)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_105),
.Y(n_114)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_66),
.B(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_35),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_33),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_132),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_74),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_138),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_23),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_135),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_140),
.B1(n_145),
.B2(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_3),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_10),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_101),
.B(n_91),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_99),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_73),
.A2(n_99),
.B1(n_88),
.B2(n_72),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_107),
.B1(n_65),
.B2(n_103),
.Y(n_151)
);

CKINVDCx6p67_ASAP7_75t_R g142 ( 
.A(n_96),
.Y(n_142)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_8),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_73),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_81),
.Y(n_146)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

CKINVDCx12_ASAP7_75t_R g147 ( 
.A(n_65),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_97),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_79),
.B(n_9),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_11),
.C(n_13),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_156),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_90),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_160),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_146),
.B1(n_139),
.B2(n_123),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_162),
.B(n_16),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_128),
.A2(n_107),
.B1(n_97),
.B2(n_102),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_102),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_130),
.B(n_142),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_120),
.A2(n_98),
.B1(n_88),
.B2(n_75),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_130),
.B(n_114),
.C(n_138),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_98),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_75),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_157),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_11),
.B(n_13),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_185),
.B(n_14),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_185),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_116),
.A2(n_14),
.B(n_15),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_141),
.B(n_130),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_179),
.B(n_151),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_188),
.A2(n_194),
.B(n_201),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_171),
.B1(n_155),
.B2(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_197),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_199),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_148),
.B(n_119),
.C(n_127),
.D(n_117),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_146),
.Y(n_197)
);

NOR4xp25_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_161),
.C(n_162),
.D(n_174),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_215),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_127),
.B1(n_117),
.B2(n_119),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_169),
.B1(n_168),
.B2(n_178),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_160),
.B(n_15),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_203),
.B(n_218),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_208),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_112),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_211),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_151),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_167),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_217),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_157),
.A2(n_123),
.B(n_129),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_183),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_175),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_129),
.B(n_16),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_180),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_222),
.B(n_188),
.C(n_190),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_155),
.B1(n_153),
.B2(n_152),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_186),
.B1(n_190),
.B2(n_202),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_236),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_246),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_151),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_149),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_156),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_192),
.B1(n_190),
.B2(n_217),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_193),
.A2(n_182),
.B(n_158),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_243),
.B(n_245),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_205),
.A2(n_169),
.B1(n_158),
.B2(n_173),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_173),
.B1(n_154),
.B2(n_177),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_187),
.A2(n_154),
.B1(n_177),
.B2(n_183),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_154),
.C(n_177),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_215),
.C(n_200),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_256),
.B1(n_236),
.B2(n_241),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_201),
.B(n_213),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_245),
.B(n_221),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_195),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_269),
.C(n_230),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_225),
.B(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_199),
.B1(n_238),
.B2(n_229),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_270),
.B(n_216),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_199),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_227),
.C(n_247),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_275),
.C(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_276),
.B1(n_251),
.B2(n_254),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_227),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_222),
.B1(n_220),
.B2(n_235),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_235),
.C(n_243),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_268),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_250),
.B(n_244),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_188),
.B(n_219),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_279),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_190),
.B1(n_198),
.B2(n_240),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_287),
.B1(n_278),
.B2(n_272),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_260),
.B(n_244),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_199),
.C(n_204),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_259),
.C(n_263),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_282),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_293),
.A2(n_301),
.B(n_281),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_300),
.C(n_302),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_273),
.C(n_272),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_295),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_288),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_270),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_257),
.C(n_266),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_271),
.C(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

AOI321xp33_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_283),
.A3(n_253),
.B1(n_276),
.B2(n_278),
.C(n_274),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_305),
.A2(n_253),
.B(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_253),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_315),
.B(n_314),
.Y(n_327)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_314),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_302),
.C(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_317),
.B(n_295),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_249),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_319),
.Y(n_326)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_321),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_300),
.C(n_301),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_297),
.B1(n_286),
.B2(n_305),
.Y(n_323)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_323),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_293),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_311),
.C(n_316),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_208),
.Y(n_328)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_307),
.A2(n_318),
.B1(n_309),
.B2(n_315),
.Y(n_329)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

AOI31xp67_ASAP7_75t_SL g330 ( 
.A1(n_322),
.A2(n_316),
.A3(n_194),
.B(n_267),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_325),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_308),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_253),
.B(n_261),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_343),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_326),
.B(n_324),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_339),
.A2(n_340),
.B(n_341),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_332),
.A2(n_265),
.B(n_261),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_331),
.B(n_334),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_342),
.B(n_331),
.C(n_335),
.Y(n_344)
);

AOI322xp5_ASAP7_75t_L g348 ( 
.A1(n_344),
.A2(n_17),
.A3(n_204),
.B1(n_210),
.B2(n_212),
.C1(n_218),
.C2(n_346),
.Y(n_348)
);

OAI321xp33_ASAP7_75t_L g347 ( 
.A1(n_345),
.A2(n_199),
.A3(n_265),
.B1(n_249),
.B2(n_229),
.C(n_214),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_347),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_348),
.C(n_212),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_17),
.Y(n_351)
);


endmodule