module fake_netlist_1_10346_n_28 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_0), .B(n_1), .Y(n_17) );
CKINVDCx8_ASAP7_75t_R g18 ( .A(n_13), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
OAI22xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_15), .B1(n_16), .B2(n_12), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NAND5xp2_ASAP7_75t_SL g22 ( .A(n_21), .B(n_18), .C(n_17), .D(n_7), .E(n_9), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_4), .Y(n_23) );
XNOR2x1_ASAP7_75t_L g24 ( .A(n_23), .B(n_11), .Y(n_24) );
NAND2xp33_ASAP7_75t_R g25 ( .A(n_23), .B(n_5), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OR2x6_ASAP7_75t_L g27 ( .A(n_26), .B(n_25), .Y(n_27) );
BUFx3_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
endmodule