module fake_jpeg_22663_n_40 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_40);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_32;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_26),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_7),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_31),
.B(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_29),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_15),
.Y(n_40)
);


endmodule