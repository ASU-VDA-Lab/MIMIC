module fake_jpeg_19859_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_2),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_15),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_26),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_28),
.B1(n_32),
.B2(n_27),
.Y(n_49)
);

AOI22x1_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_55),
.B1(n_56),
.B2(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_32),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_58),
.C(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_19),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_31),
.B1(n_25),
.B2(n_15),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_30),
.B1(n_21),
.B2(n_22),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_35),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_16),
.C(n_14),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_48),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_55),
.B1(n_49),
.B2(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_35),
.C(n_14),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_58),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_53),
.B(n_50),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_77),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_79),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_61),
.C(n_67),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_56),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_72),
.C(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_64),
.B1(n_65),
.B2(n_59),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_80),
.B(n_74),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_86),
.B(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.C(n_91),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

OAI322xp33_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_19),
.A3(n_12),
.B1(n_13),
.B2(n_18),
.C1(n_22),
.C2(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_85),
.B(n_69),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_95),
.B(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_98),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_12),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_7),
.B(n_10),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_10),
.A3(n_13),
.B1(n_18),
.B2(n_24),
.C1(n_46),
.C2(n_100),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);


endmodule