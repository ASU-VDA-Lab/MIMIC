module fake_netlist_6_3297_n_5186 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5186);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5186;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_741;
wire n_1351;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2786;
wire n_1971;
wire n_1781;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_989;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_3277;
wire n_2548;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_1094;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_4334;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_757;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_847;
wire n_851;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_2995;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4192;
wire n_4109;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_4543;
wire n_740;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_1003;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_825;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_2323;
wire n_2784;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_3407;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_4330;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_2316;
wire n_1771;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_2771;
wire n_3020;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_975;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

INVx1_ASAP7_75t_L g706 ( 
.A(n_508),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_506),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_238),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_574),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_467),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_329),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_395),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_576),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_394),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_624),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_679),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_403),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_555),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_420),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_422),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_547),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_499),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_688),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_654),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_240),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_655),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_71),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_130),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_434),
.Y(n_729)
);

BUFx5_ASAP7_75t_L g730 ( 
.A(n_134),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_659),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_491),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_21),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_387),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_552),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_276),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_372),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_245),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_498),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_88),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_213),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_106),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_56),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_630),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_700),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_49),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_192),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_515),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_43),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_180),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_203),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_412),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_103),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_204),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_113),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_473),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_58),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_622),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_367),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_198),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_702),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_395),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_680),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_86),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_337),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_120),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_55),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_143),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_526),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_349),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_195),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_355),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_384),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_471),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_413),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_656),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_76),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_231),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_641),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_320),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_180),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_573),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_166),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_52),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_216),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_333),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_372),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_245),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_283),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_201),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_307),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_459),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_52),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_165),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_153),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_497),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_661),
.Y(n_798)
);

BUFx8_ASAP7_75t_SL g799 ( 
.A(n_377),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_524),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_624),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_208),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_458),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_570),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_217),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_100),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_237),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_695),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_619),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_159),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_190),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_170),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_614),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_155),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_618),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_547),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_557),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_494),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_641),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_125),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_429),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_398),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_128),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_387),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_98),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_426),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_678),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_9),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_255),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_437),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_78),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_167),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_445),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_168),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_616),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_610),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_321),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_76),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_357),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_42),
.Y(n_840)
);

BUFx5_ASAP7_75t_L g841 ( 
.A(n_59),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_160),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_509),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_164),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_617),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_493),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_75),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_90),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_84),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_616),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_117),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_456),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_464),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_439),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_551),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_337),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_62),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_112),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_128),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_591),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_210),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_544),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_108),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_552),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_74),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_670),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_56),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_39),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_642),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_472),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_566),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_84),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_610),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_642),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_606),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_254),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_217),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_262),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_492),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_62),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_295),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_440),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_638),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_316),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_284),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_35),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_150),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_210),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_623),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_517),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_665),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_541),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_316),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_386),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_188),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_499),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_188),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_635),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_379),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_672),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_214),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_111),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_692),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_149),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_415),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_205),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_205),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_671),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_102),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_493),
.Y(n_910)
);

CKINVDCx16_ASAP7_75t_R g911 ( 
.A(n_527),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_149),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_585),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_571),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_339),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_281),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_592),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_116),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_516),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_261),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_448),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_415),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_490),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_260),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_406),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_177),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_615),
.Y(n_927)
);

CKINVDCx16_ASAP7_75t_R g928 ( 
.A(n_233),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_157),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_57),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_407),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_173),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_453),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_138),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_199),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_412),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_574),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_465),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_7),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_520),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_324),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_307),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_451),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_95),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_485),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_506),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_328),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_643),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_687),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_388),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_631),
.Y(n_951)
);

BUFx2_ASAP7_75t_SL g952 ( 
.A(n_72),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_634),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_206),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_331),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_97),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_629),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_326),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_489),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_621),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_223),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_175),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_585),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_525),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_383),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_544),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_561),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_586),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_305),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_568),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_243),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_75),
.Y(n_972)
);

BUFx5_ASAP7_75t_L g973 ( 
.A(n_352),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_473),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_101),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_264),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_623),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_162),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_287),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_203),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_429),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_315),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_285),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_121),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_452),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_266),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_185),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_177),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_126),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_617),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_455),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_261),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_541),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_572),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_88),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_619),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_368),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_436),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_133),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_646),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_468),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_536),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_636),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_578),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_542),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_555),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_198),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_446),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_72),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_620),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_401),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_278),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_100),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_364),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_579),
.Y(n_1015)
);

BUFx5_ASAP7_75t_L g1016 ( 
.A(n_490),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_4),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_351),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_551),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_394),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_609),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_310),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_4),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_197),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_402),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_13),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_240),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_416),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_548),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_197),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_178),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_553),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_199),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_663),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_594),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_333),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_80),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_553),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_509),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_7),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_227),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_730),
.Y(n_1042)
);

NOR2xp67_ASAP7_75t_L g1043 ( 
.A(n_890),
.B(n_0),
.Y(n_1043)
);

INVxp67_ASAP7_75t_SL g1044 ( 
.A(n_826),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_716),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_799),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_730),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_845),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_730),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_718),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_730),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_730),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_730),
.Y(n_1053)
);

CKINVDCx16_ASAP7_75t_R g1054 ( 
.A(n_766),
.Y(n_1054)
);

CKINVDCx14_ASAP7_75t_R g1055 ( 
.A(n_724),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_730),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_758),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_799),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_769),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_768),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_841),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_841),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_722),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_841),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_841),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_911),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_841),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_841),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_L g1069 ( 
.A(n_922),
.B(n_0),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_841),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_973),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_815),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_928),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_908),
.B(n_2),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_973),
.Y(n_1075)
);

CKINVDCx16_ASAP7_75t_R g1076 ( 
.A(n_723),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_722),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_973),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_707),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_708),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_973),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_709),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_973),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_973),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_973),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1016),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1016),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_710),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1016),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_712),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1016),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_718),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_752),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1016),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1016),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1016),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_751),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_752),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_751),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_800),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_800),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1026),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1026),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_718),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_718),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_855),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_855),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_713),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_830),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_855),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_855),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_879),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_879),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_908),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_879),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_879),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_894),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_894),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_894),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_894),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_870),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_963),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_963),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_963),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_963),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_L g1126 ( 
.A(n_970),
.B(n_1),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_971),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_971),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_726),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_971),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_971),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_980),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_980),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_980),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_980),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1025),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_731),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_762),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1025),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_777),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1025),
.Y(n_1141)
);

INVxp33_ASAP7_75t_L g1142 ( 
.A(n_741),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1025),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_706),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_711),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_736),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_715),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_734),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_714),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_987),
.B(n_1),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_717),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_746),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_764),
.Y(n_1153)
);

CKINVDCx16_ASAP7_75t_R g1154 ( 
.A(n_723),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_733),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_753),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_719),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_735),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_737),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_740),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_741),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_736),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_743),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_745),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_748),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_753),
.Y(n_1166)
);

INVxp67_ASAP7_75t_SL g1167 ( 
.A(n_827),
.Y(n_1167)
);

INVxp67_ASAP7_75t_SL g1168 ( 
.A(n_866),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_756),
.Y(n_1169)
);

CKINVDCx16_ASAP7_75t_R g1170 ( 
.A(n_736),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_744),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_757),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_763),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_767),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_773),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_774),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_776),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_721),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_778),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_734),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_738),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_779),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_725),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_738),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_780),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_891),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_781),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_727),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_949),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_728),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_783),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_729),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_784),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_794),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_793),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_804),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_739),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_744),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_794),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_798),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_808),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_805),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_754),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_775),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_794),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_900),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_903),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_754),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1034),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_809),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_810),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_742),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_884),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_816),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_747),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_820),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_749),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_739),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_770),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_775),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_884),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_825),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_832),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_834),
.Y(n_1224)
);

CKINVDCx16_ASAP7_75t_R g1225 ( 
.A(n_884),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_837),
.Y(n_1226)
);

INVxp33_ASAP7_75t_L g1227 ( 
.A(n_770),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_788),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_750),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_788),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_755),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_838),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_840),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_759),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_760),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_765),
.Y(n_1236)
);

INVxp67_ASAP7_75t_SL g1237 ( 
.A(n_829),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_847),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_856),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_857),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_771),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_829),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_858),
.Y(n_1243)
);

INVxp33_ASAP7_75t_SL g1244 ( 
.A(n_874),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_871),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_874),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_931),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_931),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_859),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_862),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_882),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_871),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_901),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_732),
.B(n_2),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_906),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_772),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_782),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_907),
.Y(n_1258)
);

CKINVDCx16_ASAP7_75t_R g1259 ( 
.A(n_931),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_909),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_913),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_792),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_914),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_917),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_785),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_786),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_787),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_921),
.Y(n_1268)
);

NOR2xp67_ASAP7_75t_L g1269 ( 
.A(n_732),
.B(n_3),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_923),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_925),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_926),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_927),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_982),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1038),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_929),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_936),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_792),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_877),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_877),
.Y(n_1280)
);

XOR2xp5_ASAP7_75t_L g1281 ( 
.A(n_803),
.B(n_3),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_938),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_789),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_982),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_932),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_950),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_803),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_790),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_956),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_964),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_989),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_791),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1003),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1007),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1009),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1011),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1014),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_982),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1024),
.Y(n_1299)
);

INVxp33_ASAP7_75t_L g1300 ( 
.A(n_932),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1029),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_957),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_957),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_795),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_958),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_796),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_812),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_958),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_967),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_797),
.Y(n_1310)
);

INVxp33_ASAP7_75t_SL g1311 ( 
.A(n_1038),
.Y(n_1311)
);

BUFx5_ASAP7_75t_L g1312 ( 
.A(n_967),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1015),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1015),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_952),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_848),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_848),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_854),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_854),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_896),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_896),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_993),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_993),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_720),
.B(n_5),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_801),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_802),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_806),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_807),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_811),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_813),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_814),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1039),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_818),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_819),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_812),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_823),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_824),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_828),
.Y(n_1338)
);

INVxp33_ASAP7_75t_SL g1339 ( 
.A(n_1039),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_831),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_833),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_835),
.Y(n_1342)
);

CKINVDCx14_ASAP7_75t_R g1343 ( 
.A(n_817),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_836),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_839),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_842),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_843),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_844),
.Y(n_1348)
);

NOR2xp67_ASAP7_75t_L g1349 ( 
.A(n_846),
.B(n_5),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_849),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_851),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_852),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_853),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_817),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_860),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_821),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_863),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_865),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_867),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_868),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_821),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1040),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_869),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_872),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_875),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_876),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_878),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1040),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_880),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_881),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_883),
.Y(n_1371)
);

CKINVDCx14_ASAP7_75t_R g1372 ( 
.A(n_850),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_885),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_886),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_887),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_888),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_892),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_893),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_895),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_898),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_899),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_902),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_850),
.Y(n_1383)
);

INVxp67_ASAP7_75t_SL g1384 ( 
.A(n_761),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_904),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_905),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_910),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1041),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_912),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_916),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_918),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_920),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1041),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_924),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_930),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_861),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_933),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_934),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_822),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_889),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_935),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_939),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_940),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_942),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_943),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1059),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1212),
.B(n_944),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1092),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1335),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1130),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1063),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1137),
.Y(n_1412)
);

CKINVDCx16_ASAP7_75t_R g1413 ( 
.A(n_1076),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1215),
.B(n_945),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1138),
.Y(n_1415)
);

INVxp33_ASAP7_75t_SL g1416 ( 
.A(n_1058),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1104),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1063),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1105),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1352),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1106),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1110),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1384),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1077),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1399),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1111),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1217),
.B(n_946),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1219),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1140),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1112),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1400),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1113),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1077),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1093),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1093),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1114),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1115),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_SL g1438 ( 
.A(n_1348),
.Y(n_1438)
);

CKINVDCx16_ASAP7_75t_R g1439 ( 
.A(n_1154),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1200),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1116),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1180),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1229),
.B(n_947),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1201),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1231),
.B(n_948),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1207),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1117),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1059),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1118),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1098),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1209),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_1098),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1119),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1120),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1352),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1122),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1123),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1234),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1124),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1127),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1156),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1128),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1066),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1131),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1156),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1235),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1132),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1134),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1135),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1136),
.Y(n_1470)
);

INVxp67_ASAP7_75t_SL g1471 ( 
.A(n_1352),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1139),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1236),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1141),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1206),
.B(n_951),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1352),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1166),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1143),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1107),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1387),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1107),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1387),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1241),
.B(n_953),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1125),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1125),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1166),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1133),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1256),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1257),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1382),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1133),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1114),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1385),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1392),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1402),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1050),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1079),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1079),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1114),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1204),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1080),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1204),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1114),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1312),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1050),
.Y(n_1505)
);

INVxp67_ASAP7_75t_SL g1506 ( 
.A(n_1387),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1080),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1060),
.B(n_919),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1050),
.Y(n_1509)
);

CKINVDCx14_ASAP7_75t_R g1510 ( 
.A(n_1343),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1237),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1082),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1280),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1045),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1186),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1186),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1186),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_SL g1518 ( 
.A(n_1348),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1312),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1186),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1220),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1189),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1082),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1338),
.B(n_954),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1088),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1189),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1206),
.B(n_955),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1066),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1387),
.B(n_959),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1189),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1342),
.B(n_961),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1088),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1090),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1189),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1220),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1144),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1145),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1147),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1090),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1262),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1108),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1342),
.B(n_962),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_1054),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1108),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1184),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1325),
.B(n_965),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1151),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1342),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1149),
.B(n_966),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1197),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1149),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1155),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1158),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1159),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1160),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1306),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1157),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1262),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1163),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1146),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1218),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1164),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1157),
.B(n_968),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1178),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1178),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1278),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1165),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1183),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1246),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1169),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1278),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1183),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1172),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1188),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1170),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1173),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1312),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1188),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1190),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1174),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1175),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1176),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1148),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1177),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1073),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1287),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1190),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1192),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1287),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1181),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_R g1591 ( 
.A(n_1055),
.B(n_1033),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1192),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1179),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1275),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1332),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1307),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1312),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1265),
.B(n_974),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1182),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1185),
.Y(n_1600)
);

NOR2xp67_ASAP7_75t_L g1601 ( 
.A(n_1368),
.B(n_651),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1312),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1265),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1266),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1307),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1266),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1354),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1187),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1267),
.B(n_975),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1267),
.B(n_976),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1191),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1283),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1193),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1195),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1362),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1196),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1073),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1202),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1283),
.B(n_977),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1210),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1328),
.B(n_1329),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1354),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1288),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1393),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1306),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1211),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1214),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1216),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1222),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1223),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1224),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1226),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1232),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1233),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1219),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1356),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1238),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1239),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1288),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1240),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1356),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1243),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1292),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1361),
.Y(n_1644)
);

CKINVDCx20_ASAP7_75t_R g1645 ( 
.A(n_1361),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_1383),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1249),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1292),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1383),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1304),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1250),
.Y(n_1651)
);

NOR2xp67_ASAP7_75t_L g1652 ( 
.A(n_1388),
.B(n_652),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1304),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1251),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1253),
.Y(n_1655)
);

BUFx10_ASAP7_75t_L g1656 ( 
.A(n_1046),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1255),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1258),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1330),
.B(n_978),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1260),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1261),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1284),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1396),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1263),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1264),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1310),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1268),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1270),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1310),
.B(n_979),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1338),
.B(n_981),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1271),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1272),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1273),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1276),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1219),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1326),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1326),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1277),
.Y(n_1678)
);

NOR2xp67_ASAP7_75t_L g1679 ( 
.A(n_1331),
.B(n_653),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1331),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1282),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1286),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1334),
.B(n_985),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1334),
.B(n_986),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1289),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1336),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1045),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1290),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1291),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1396),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1336),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1340),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1293),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1340),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1345),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1294),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1295),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1296),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1312),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1213),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1129),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1297),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1299),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1301),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1097),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_1343),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1099),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1345),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1100),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1101),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1333),
.B(n_988),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1496),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1496),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1548),
.B(n_1167),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1428),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1492),
.A2(n_1047),
.B(n_1042),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1549),
.A2(n_1347),
.B1(n_1357),
.B2(n_1351),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1420),
.B(n_1168),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1509),
.Y(n_1719)
);

AND2x2_ASAP7_75t_SL g1720 ( 
.A(n_1531),
.B(n_1074),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1509),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1563),
.A2(n_1347),
.B1(n_1357),
.B2(n_1351),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1705),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1479),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_L g1725 ( 
.A(n_1621),
.B(n_1254),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1598),
.A2(n_1360),
.B1(n_1371),
.B2(n_1365),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1514),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1707),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1455),
.B(n_1055),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1428),
.Y(n_1730)
);

INVx4_ASAP7_75t_L g1731 ( 
.A(n_1428),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1471),
.B(n_1350),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1428),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1514),
.B(n_1161),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1609),
.A2(n_1365),
.B1(n_1371),
.B2(n_1360),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1687),
.Y(n_1736)
);

OA21x2_ASAP7_75t_L g1737 ( 
.A1(n_1499),
.A2(n_1052),
.B(n_1051),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1709),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1635),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1481),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1484),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1476),
.B(n_1350),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1423),
.B(n_1327),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1687),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1662),
.Y(n_1745)
);

BUFx8_ASAP7_75t_L g1746 ( 
.A(n_1438),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1635),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1710),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1536),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1485),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1701),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1635),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1701),
.B(n_1161),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1480),
.B(n_1171),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1610),
.A2(n_1669),
.B1(n_1683),
.B2(n_1619),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1537),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1482),
.B(n_1353),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1408),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1635),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1538),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1436),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1506),
.B(n_1353),
.Y(n_1762)
);

AND2x6_ASAP7_75t_L g1763 ( 
.A(n_1524),
.B(n_1377),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1436),
.Y(n_1764)
);

AND2x2_ASAP7_75t_SL g1765 ( 
.A(n_1542),
.B(n_1324),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1601),
.B(n_1171),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1425),
.B(n_1327),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1431),
.A2(n_1311),
.B1(n_1339),
.B2(n_1244),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1487),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1436),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1675),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1410),
.B(n_1377),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1547),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1511),
.B(n_1244),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1675),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1556),
.A2(n_1339),
.B1(n_1311),
.B2(n_1057),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_L g1777 ( 
.A(n_1546),
.B(n_1312),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1491),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1504),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1552),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1529),
.B(n_1394),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1504),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1625),
.B(n_1394),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1675),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1560),
.B(n_1358),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1684),
.A2(n_1375),
.B1(n_1379),
.B2(n_1374),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1513),
.Y(n_1787)
);

BUFx12f_ASAP7_75t_L g1788 ( 
.A(n_1656),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1503),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1409),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1519),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1553),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1670),
.B(n_1358),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1515),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1554),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1706),
.A2(n_864),
.B1(n_873),
.B2(n_861),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1516),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1517),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1520),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1555),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1522),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1559),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1526),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1562),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1508),
.B(n_1369),
.Y(n_1805)
);

INVx6_ASAP7_75t_L g1806 ( 
.A(n_1543),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1652),
.B(n_1679),
.Y(n_1807)
);

INVx4_ASAP7_75t_L g1808 ( 
.A(n_1519),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1700),
.B(n_1369),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1475),
.B(n_1397),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1530),
.Y(n_1811)
);

AND2x6_ASAP7_75t_L g1812 ( 
.A(n_1577),
.B(n_1401),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1567),
.B(n_1198),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1442),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1534),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1577),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1597),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1545),
.B(n_1397),
.Y(n_1818)
);

CKINVDCx6p67_ASAP7_75t_R g1819 ( 
.A(n_1438),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1505),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1417),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1550),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1561),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1597),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1706),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1570),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1573),
.B(n_1198),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1659),
.B(n_1401),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1602),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1576),
.B(n_1203),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1407),
.A2(n_1375),
.B1(n_1379),
.B2(n_1374),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1580),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1581),
.B(n_1203),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1582),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1711),
.B(n_1337),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1584),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1419),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1602),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1593),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1569),
.B(n_1414),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1599),
.B(n_1208),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1527),
.B(n_1427),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1600),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1699),
.Y(n_1844)
);

CKINVDCx16_ASAP7_75t_R g1845 ( 
.A(n_1575),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1583),
.Y(n_1846)
);

INVx5_ASAP7_75t_L g1847 ( 
.A(n_1699),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1608),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1443),
.B(n_1445),
.Y(n_1849)
);

INVxp67_ASAP7_75t_SL g1850 ( 
.A(n_1611),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1613),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1483),
.B(n_1199),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1590),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1594),
.B(n_1199),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1595),
.B(n_1380),
.Y(n_1855)
);

CKINVDCx16_ASAP7_75t_R g1856 ( 
.A(n_1413),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1421),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1614),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1422),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1426),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1616),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1618),
.B(n_1208),
.Y(n_1862)
);

OAI21x1_ASAP7_75t_L g1863 ( 
.A1(n_1430),
.A2(n_1062),
.B(n_1049),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1432),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1437),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1441),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1447),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1449),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1453),
.Y(n_1869)
);

OA21x2_ASAP7_75t_L g1870 ( 
.A1(n_1454),
.A2(n_1056),
.B(n_1053),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1456),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1620),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1591),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1457),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1626),
.Y(n_1875)
);

OAI22x1_ASAP7_75t_R g1876 ( 
.A1(n_1411),
.A2(n_873),
.B1(n_897),
.B2(n_864),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1627),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1459),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1460),
.B(n_1341),
.Y(n_1879)
);

BUFx6f_ASAP7_75t_L g1880 ( 
.A(n_1462),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1628),
.B(n_1228),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1464),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1467),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1468),
.B(n_1344),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1615),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1469),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1629),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1470),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1630),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1472),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1624),
.A2(n_1069),
.B1(n_1126),
.B2(n_1043),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1631),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1632),
.B(n_1380),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1510),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1633),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1406),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1634),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1474),
.Y(n_1898)
);

CKINVDCx16_ASAP7_75t_R g1899 ( 
.A(n_1439),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1478),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1637),
.Y(n_1901)
);

OAI21x1_ASAP7_75t_L g1902 ( 
.A1(n_1638),
.A2(n_1062),
.B(n_1049),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1448),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_SL g1904 ( 
.A1(n_1411),
.A2(n_915),
.B1(n_969),
.B2(n_897),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1640),
.B(n_1346),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1642),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1647),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1651),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1654),
.Y(n_1909)
);

INVx6_ASAP7_75t_L g1910 ( 
.A(n_1656),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1418),
.A2(n_969),
.B1(n_972),
.B2(n_915),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1655),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1657),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1412),
.B(n_1404),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1658),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1660),
.Y(n_1916)
);

CKINVDCx16_ASAP7_75t_R g1917 ( 
.A(n_1510),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1661),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1664),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1665),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1667),
.B(n_1228),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1668),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1671),
.A2(n_1070),
.B(n_1067),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1591),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1672),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1673),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1674),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1678),
.B(n_1355),
.Y(n_1928)
);

OA21x2_ASAP7_75t_L g1929 ( 
.A1(n_1681),
.A2(n_1064),
.B(n_1061),
.Y(n_1929)
);

OA22x2_ASAP7_75t_SL g1930 ( 
.A1(n_1518),
.A2(n_1048),
.B1(n_1044),
.B2(n_1372),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1682),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1685),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1688),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1689),
.B(n_1359),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1693),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1696),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1639),
.B(n_1404),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1697),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1698),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1415),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1702),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1703),
.Y(n_1942)
);

OAI21x1_ASAP7_75t_L g1943 ( 
.A1(n_1704),
.A2(n_1070),
.B(n_1067),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1650),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1691),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1429),
.B(n_1405),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1440),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1444),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1458),
.B(n_1405),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1463),
.B(n_1230),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1528),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1446),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1585),
.B(n_1230),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1466),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1473),
.B(n_1363),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1617),
.Y(n_1956)
);

AOI22x1_ASAP7_75t_SL g1957 ( 
.A1(n_1418),
.A2(n_984),
.B1(n_1021),
.B2(n_972),
.Y(n_1957)
);

BUFx2_ASAP7_75t_L g1958 ( 
.A(n_1424),
.Y(n_1958)
);

BUFx12f_ASAP7_75t_L g1959 ( 
.A(n_1656),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1451),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1488),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1489),
.B(n_1205),
.Y(n_1962)
);

XOR2xp5_ASAP7_75t_L g1963 ( 
.A(n_1424),
.B(n_1372),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1433),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1490),
.B(n_1364),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1497),
.B(n_1072),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1433),
.A2(n_1021),
.B1(n_1037),
.B2(n_984),
.Y(n_1967)
);

INVxp33_ASAP7_75t_SL g1968 ( 
.A(n_1498),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1493),
.B(n_1245),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1494),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1495),
.B(n_1366),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1501),
.B(n_1245),
.Y(n_1972)
);

AND2x6_ASAP7_75t_L g1973 ( 
.A(n_1518),
.B(n_1376),
.Y(n_1973)
);

OA21x2_ASAP7_75t_L g1974 ( 
.A1(n_1507),
.A2(n_1068),
.B(n_1065),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1512),
.A2(n_1150),
.B1(n_1370),
.B2(n_1367),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1523),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1525),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1532),
.B(n_1279),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1533),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1539),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1541),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1544),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1551),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1557),
.B(n_1373),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1564),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1565),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1568),
.B(n_1378),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1708),
.B(n_1381),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1572),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1574),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_SL g1991 ( 
.A1(n_1434),
.A2(n_1037),
.B1(n_1281),
.B2(n_1225),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1578),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1579),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1587),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1588),
.Y(n_1995)
);

AOI22x1_ASAP7_75t_SL g1996 ( 
.A1(n_1434),
.A2(n_991),
.B1(n_992),
.B2(n_990),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1592),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1603),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1604),
.B(n_1279),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1606),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1734),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1940),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_R g2003 ( 
.A(n_1894),
.B(n_1612),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1734),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_R g2005 ( 
.A(n_1894),
.B(n_1623),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1785),
.B(n_1643),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1940),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1948),
.Y(n_2008)
);

AND3x2_ASAP7_75t_L g2009 ( 
.A(n_1790),
.B(n_1121),
.C(n_1109),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1902),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1902),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1913),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1790),
.Y(n_2013)
);

AND3x2_ASAP7_75t_L g2014 ( 
.A(n_1745),
.B(n_1924),
.C(n_1873),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1734),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_R g2016 ( 
.A(n_1856),
.B(n_1899),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1948),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1842),
.B(n_1648),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1948),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1948),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1923),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1923),
.Y(n_2022)
);

NAND2xp33_ASAP7_75t_R g2023 ( 
.A(n_1958),
.B(n_1653),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1961),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1961),
.Y(n_2025)
);

BUFx3_ASAP7_75t_L g2026 ( 
.A(n_1727),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1849),
.B(n_1666),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1961),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1961),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1753),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_1845),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1753),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1968),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_SL g2034 ( 
.A(n_1990),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1968),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1917),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1943),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1964),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1788),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_1806),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1788),
.Y(n_2041)
);

INVx1_ASAP7_75t_SL g2042 ( 
.A(n_1805),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1753),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1813),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1943),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1863),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1959),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1959),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1863),
.Y(n_2049)
);

BUFx2_ASAP7_75t_L g2050 ( 
.A(n_1956),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1819),
.Y(n_2051)
);

CKINVDCx20_ASAP7_75t_R g2052 ( 
.A(n_1806),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1819),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1990),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1716),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1954),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1813),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1954),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1983),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1983),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1727),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1983),
.Y(n_2062)
);

CKINVDCx20_ASAP7_75t_R g2063 ( 
.A(n_1963),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1983),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1989),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1989),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1989),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1989),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1813),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1910),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_1808),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1910),
.Y(n_2072)
);

BUFx6f_ASAP7_75t_L g2073 ( 
.A(n_1913),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1827),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_R g2075 ( 
.A(n_1980),
.B(n_1676),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_1796),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1972),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1827),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1827),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1910),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1830),
.Y(n_2081)
);

CKINVDCx20_ASAP7_75t_R g2082 ( 
.A(n_1904),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1849),
.B(n_1677),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1854),
.B(n_1680),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1807),
.B(n_1386),
.Y(n_2085)
);

AOI21x1_ASAP7_75t_L g2086 ( 
.A1(n_1828),
.A2(n_1075),
.B(n_1071),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_1911),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1830),
.Y(n_2088)
);

CKINVDCx20_ASAP7_75t_R g2089 ( 
.A(n_1967),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1969),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1806),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1830),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1716),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1716),
.Y(n_2094)
);

CKINVDCx20_ASAP7_75t_R g2095 ( 
.A(n_1991),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1746),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1746),
.Y(n_2097)
);

NAND2xp33_ASAP7_75t_R g2098 ( 
.A(n_1974),
.B(n_1686),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_1966),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1737),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1746),
.Y(n_2101)
);

CKINVDCx20_ASAP7_75t_R g2102 ( 
.A(n_1876),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1993),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_1972),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1993),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1980),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1737),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1985),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1985),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1737),
.Y(n_2110)
);

CKINVDCx20_ASAP7_75t_R g2111 ( 
.A(n_1825),
.Y(n_2111)
);

CKINVDCx20_ASAP7_75t_R g2112 ( 
.A(n_1956),
.Y(n_2112)
);

NOR2xp67_ASAP7_75t_L g2113 ( 
.A(n_1717),
.B(n_1692),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1833),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1870),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_L g2116 ( 
.A(n_1755),
.B(n_1694),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_1962),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1870),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1807),
.B(n_1389),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1986),
.Y(n_2120)
);

NOR2xp67_ASAP7_75t_L g2121 ( 
.A(n_1722),
.B(n_1726),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1833),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1807),
.B(n_1720),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_1972),
.Y(n_2124)
);

INVxp33_ASAP7_75t_L g2125 ( 
.A(n_1774),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1833),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1986),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1994),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1870),
.Y(n_2129)
);

CKINVDCx20_ASAP7_75t_R g2130 ( 
.A(n_1962),
.Y(n_2130)
);

CKINVDCx20_ASAP7_75t_R g2131 ( 
.A(n_1914),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_1994),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_1997),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1997),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1947),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1947),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1736),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1720),
.B(n_1390),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1952),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1841),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_1952),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1841),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1970),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1970),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1960),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1949),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_1736),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1841),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1779),
.Y(n_2149)
);

INVxp67_ASAP7_75t_L g2150 ( 
.A(n_1814),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_1744),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1744),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1862),
.Y(n_2153)
);

CKINVDCx20_ASAP7_75t_R g2154 ( 
.A(n_1914),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1862),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1751),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1751),
.Y(n_2157)
);

CKINVDCx20_ASAP7_75t_R g2158 ( 
.A(n_1946),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1862),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1881),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1831),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1735),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1779),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1786),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1977),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1782),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1977),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1981),
.Y(n_2168)
);

BUFx2_ASAP7_75t_L g2169 ( 
.A(n_1846),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1881),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_1981),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1982),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_1982),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1881),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1995),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_1995),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1840),
.B(n_1695),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1765),
.B(n_1221),
.Y(n_2178)
);

HB1xp67_ASAP7_75t_L g2179 ( 
.A(n_1978),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1998),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1782),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_1808),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1998),
.Y(n_2183)
);

CKINVDCx20_ASAP7_75t_R g2184 ( 
.A(n_1946),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1976),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1921),
.Y(n_2186)
);

CKINVDCx20_ASAP7_75t_R g2187 ( 
.A(n_1957),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1979),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_R g2189 ( 
.A(n_1992),
.B(n_1435),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_2000),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1921),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_1978),
.Y(n_2192)
);

INVxp67_ASAP7_75t_L g2193 ( 
.A(n_1814),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1965),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1971),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_1973),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1973),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1852),
.B(n_1416),
.Y(n_2198)
);

AOI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_1765),
.A2(n_1416),
.B1(n_1391),
.B2(n_1398),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_1973),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1921),
.Y(n_2201)
);

CKINVDCx20_ASAP7_75t_R g2202 ( 
.A(n_1846),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_R g2203 ( 
.A(n_1725),
.B(n_1589),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1912),
.Y(n_2204)
);

CKINVDCx20_ASAP7_75t_R g2205 ( 
.A(n_1853),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1973),
.Y(n_2206)
);

CKINVDCx20_ASAP7_75t_R g2207 ( 
.A(n_1853),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1973),
.Y(n_2208)
);

CKINVDCx20_ASAP7_75t_R g2209 ( 
.A(n_1885),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1816),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_1978),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_1955),
.Y(n_2212)
);

BUFx2_ASAP7_75t_L g2213 ( 
.A(n_1885),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1999),
.B(n_1969),
.Y(n_2214)
);

CKINVDCx20_ASAP7_75t_R g2215 ( 
.A(n_1822),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_R g2216 ( 
.A(n_1725),
.B(n_1589),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1912),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1768),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_1988),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1776),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1816),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_1984),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1714),
.B(n_1248),
.Y(n_2223)
);

BUFx10_ASAP7_75t_L g2224 ( 
.A(n_1774),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1919),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_1987),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1817),
.Y(n_2227)
);

CKINVDCx16_ASAP7_75t_R g2228 ( 
.A(n_1937),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_1969),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_1822),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1817),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_1823),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_1823),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_R g2234 ( 
.A(n_1944),
.B(n_1605),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_1975),
.Y(n_2235)
);

BUFx3_ASAP7_75t_L g2236 ( 
.A(n_1848),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1919),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1999),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1935),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_R g2240 ( 
.A(n_1945),
.B(n_1605),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1935),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_1999),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_1848),
.B(n_1315),
.Y(n_2243)
);

BUFx10_ASAP7_75t_L g2244 ( 
.A(n_1893),
.Y(n_2244)
);

OA21x2_ASAP7_75t_L g2245 ( 
.A1(n_1824),
.A2(n_1083),
.B(n_1081),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1824),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_1855),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1893),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1996),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1809),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1829),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1829),
.Y(n_2252)
);

INVxp67_ASAP7_75t_L g2253 ( 
.A(n_1818),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1895),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1936),
.Y(n_2255)
);

CKINVDCx20_ASAP7_75t_R g2256 ( 
.A(n_1896),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1895),
.Y(n_2257)
);

NOR2xp67_ASAP7_75t_L g2258 ( 
.A(n_1896),
.B(n_1395),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_1793),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_1906),
.Y(n_2260)
);

INVxp67_ASAP7_75t_L g2261 ( 
.A(n_1743),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_1906),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1844),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1787),
.Y(n_2264)
);

BUFx10_ASAP7_75t_L g2265 ( 
.A(n_1950),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1787),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_R g2267 ( 
.A(n_1777),
.B(n_1644),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_1835),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_1767),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1936),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_1951),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_1913),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1758),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1939),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_1758),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1939),
.Y(n_2276)
);

CKINVDCx5p33_ASAP7_75t_R g2277 ( 
.A(n_1903),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_1903),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_1781),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_1950),
.Y(n_2280)
);

NOR2xp67_ASAP7_75t_L g2281 ( 
.A(n_1729),
.B(n_1403),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_1844),
.A2(n_1078),
.B(n_1084),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_R g2283 ( 
.A(n_1777),
.B(n_1646),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_1808),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_1891),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_1913),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1929),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_R g2288 ( 
.A(n_1920),
.B(n_1646),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_1950),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_1953),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1749),
.Y(n_2291)
);

NAND2xp33_ASAP7_75t_L g2292 ( 
.A(n_1763),
.B(n_1058),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_1953),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1929),
.Y(n_2294)
);

CKINVDCx16_ASAP7_75t_R g2295 ( 
.A(n_1953),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1783),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_1850),
.B(n_1259),
.Y(n_2297)
);

INVx3_ASAP7_75t_L g2298 ( 
.A(n_1929),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1724),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_1772),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_1905),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1763),
.B(n_1732),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_1928),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1756),
.Y(n_2304)
);

NOR2xp67_ASAP7_75t_L g2305 ( 
.A(n_1920),
.B(n_1162),
.Y(n_2305)
);

NAND2xp33_ASAP7_75t_R g2306 ( 
.A(n_1974),
.B(n_994),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1760),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1934),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_1915),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1915),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1773),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1780),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_1791),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1792),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_1850),
.B(n_1142),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1915),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_1974),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1724),
.Y(n_2318)
);

CKINVDCx5p33_ASAP7_75t_R g2319 ( 
.A(n_1915),
.Y(n_2319)
);

INVx3_ASAP7_75t_L g2320 ( 
.A(n_1791),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_1916),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_2026),
.B(n_2061),
.Y(n_2322)
);

NAND2x1p5_ASAP7_75t_L g2323 ( 
.A(n_2071),
.B(n_1932),
.Y(n_2323)
);

AOI22xp33_ASAP7_75t_L g2324 ( 
.A1(n_2123),
.A2(n_1763),
.B1(n_1812),
.B2(n_1754),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2149),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2317),
.A2(n_1763),
.B1(n_1812),
.B2(n_1269),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2268),
.B(n_1918),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2315),
.B(n_1763),
.Y(n_2328)
);

INVxp67_ASAP7_75t_SL g2329 ( 
.A(n_2071),
.Y(n_2329)
);

HB1xp67_ASAP7_75t_L g2330 ( 
.A(n_2013),
.Y(n_2330)
);

NAND3xp33_ASAP7_75t_L g2331 ( 
.A(n_2018),
.B(n_2116),
.C(n_2297),
.Y(n_2331)
);

CKINVDCx11_ASAP7_75t_R g2332 ( 
.A(n_2031),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2001),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2149),
.Y(n_2334)
);

INVx2_ASAP7_75t_SL g2335 ( 
.A(n_2169),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_2026),
.Y(n_2336)
);

INVx4_ASAP7_75t_L g2337 ( 
.A(n_2008),
.Y(n_2337)
);

BUFx2_ASAP7_75t_L g2338 ( 
.A(n_2215),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2279),
.B(n_1754),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_2213),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2138),
.A2(n_1810),
.B1(n_1757),
.B2(n_1762),
.Y(n_2341)
);

BUFx3_ASAP7_75t_L g2342 ( 
.A(n_2040),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2071),
.B(n_1754),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2163),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_2016),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2004),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2163),
.Y(n_2347)
);

BUFx4f_ASAP7_75t_L g2348 ( 
.A(n_2050),
.Y(n_2348)
);

OR2x6_ASAP7_75t_L g2349 ( 
.A(n_2038),
.B(n_1712),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2015),
.Y(n_2350)
);

INVx4_ASAP7_75t_L g2351 ( 
.A(n_2017),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2182),
.B(n_1742),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2166),
.Y(n_2353)
);

INVx3_ASAP7_75t_L g2354 ( 
.A(n_2012),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2182),
.B(n_2284),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2030),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2182),
.B(n_1718),
.Y(n_2357)
);

INVx6_ASAP7_75t_L g2358 ( 
.A(n_2265),
.Y(n_2358)
);

INVx4_ASAP7_75t_L g2359 ( 
.A(n_2019),
.Y(n_2359)
);

INVx2_ASAP7_75t_SL g2360 ( 
.A(n_2230),
.Y(n_2360)
);

OAI22xp33_ASAP7_75t_L g2361 ( 
.A1(n_2125),
.A2(n_1227),
.B1(n_1300),
.B2(n_1142),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2125),
.B(n_1435),
.Y(n_2362)
);

NAND2xp33_ASAP7_75t_L g2363 ( 
.A(n_2309),
.B(n_1812),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2032),
.Y(n_2364)
);

CKINVDCx20_ASAP7_75t_R g2365 ( 
.A(n_2031),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2042),
.B(n_2006),
.Y(n_2366)
);

INVx4_ASAP7_75t_L g2367 ( 
.A(n_2020),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2166),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_2248),
.B(n_1450),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2284),
.B(n_1791),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2214),
.Y(n_2371)
);

CKINVDCx5p33_ASAP7_75t_R g2372 ( 
.A(n_2002),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2043),
.Y(n_2373)
);

AOI22xp33_ASAP7_75t_L g2374 ( 
.A1(n_2121),
.A2(n_1812),
.B1(n_941),
.B2(n_960),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2284),
.B(n_1838),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2012),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2296),
.B(n_1838),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2300),
.B(n_1932),
.Y(n_2378)
);

BUFx2_ASAP7_75t_L g2379 ( 
.A(n_2215),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2261),
.B(n_2298),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2259),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_SL g2382 ( 
.A(n_2024),
.B(n_1812),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2044),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2057),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2069),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2298),
.B(n_1942),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2298),
.B(n_1942),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2012),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_2194),
.B(n_1450),
.Y(n_2389)
);

INVx1_ASAP7_75t_SL g2390 ( 
.A(n_2232),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2301),
.B(n_1820),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_2061),
.Y(n_2392)
);

INVx4_ASAP7_75t_L g2393 ( 
.A(n_2025),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2099),
.B(n_1713),
.Y(n_2394)
);

CKINVDCx20_ASAP7_75t_R g2395 ( 
.A(n_2052),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2181),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2303),
.B(n_1820),
.Y(n_2397)
);

INVx5_ASAP7_75t_L g2398 ( 
.A(n_2012),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2195),
.B(n_1452),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2074),
.Y(n_2400)
);

INVx4_ASAP7_75t_SL g2401 ( 
.A(n_2034),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2308),
.B(n_2219),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2181),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2078),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2084),
.B(n_1194),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2210),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2210),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2221),
.Y(n_2408)
);

INVx5_ASAP7_75t_L g2409 ( 
.A(n_2073),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2079),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2081),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2007),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2221),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2088),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2177),
.B(n_1298),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2092),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_2027),
.B(n_1452),
.Y(n_2417)
);

CKINVDCx20_ASAP7_75t_R g2418 ( 
.A(n_2003),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2264),
.B(n_1931),
.Y(n_2419)
);

INVx4_ASAP7_75t_SL g2420 ( 
.A(n_2034),
.Y(n_2420)
);

INVxp67_ASAP7_75t_SL g2421 ( 
.A(n_2073),
.Y(n_2421)
);

NAND2xp33_ASAP7_75t_L g2422 ( 
.A(n_2310),
.B(n_1916),
.Y(n_2422)
);

AOI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2204),
.A2(n_1918),
.B1(n_1922),
.B2(n_1916),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2083),
.B(n_1461),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_2202),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2266),
.B(n_1931),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2114),
.Y(n_2427)
);

NAND2xp33_ASAP7_75t_L g2428 ( 
.A(n_2316),
.B(n_1916),
.Y(n_2428)
);

AND2x6_ASAP7_75t_SL g2429 ( 
.A(n_2198),
.B(n_1316),
.Y(n_2429)
);

BUFx4f_ASAP7_75t_L g2430 ( 
.A(n_2090),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2227),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2115),
.B(n_1766),
.Y(n_2432)
);

NOR2x1p5_ASAP7_75t_L g2433 ( 
.A(n_2070),
.B(n_1213),
.Y(n_2433)
);

NAND2x1p5_ASAP7_75t_L g2434 ( 
.A(n_2073),
.B(n_1775),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2122),
.Y(n_2435)
);

AOI22xp33_ASAP7_75t_L g2436 ( 
.A1(n_2217),
.A2(n_1922),
.B1(n_1926),
.B2(n_1918),
.Y(n_2436)
);

INVx2_ASAP7_75t_SL g2437 ( 
.A(n_2233),
.Y(n_2437)
);

BUFx4f_ASAP7_75t_L g2438 ( 
.A(n_2243),
.Y(n_2438)
);

AND2x6_ASAP7_75t_L g2439 ( 
.A(n_2115),
.B(n_1719),
.Y(n_2439)
);

AOI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2118),
.A2(n_983),
.B1(n_998),
.B2(n_937),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2118),
.B(n_1766),
.Y(n_2441)
);

BUFx2_ASAP7_75t_L g2442 ( 
.A(n_2202),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2223),
.B(n_1461),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2126),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_2059),
.Y(n_2445)
);

BUFx3_ASAP7_75t_L g2446 ( 
.A(n_2091),
.Y(n_2446)
);

OAI22xp33_ASAP7_75t_SL g2447 ( 
.A1(n_2135),
.A2(n_1721),
.B1(n_1002),
.B2(n_1006),
.Y(n_2447)
);

INVx2_ASAP7_75t_SL g2448 ( 
.A(n_2060),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2077),
.B(n_1348),
.Y(n_2449)
);

OR2x6_ASAP7_75t_L g2450 ( 
.A(n_2104),
.B(n_1795),
.Y(n_2450)
);

OR2x2_ASAP7_75t_L g2451 ( 
.A(n_2295),
.B(n_1800),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2137),
.B(n_1927),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2129),
.B(n_1766),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2137),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2140),
.Y(n_2455)
);

NAND2xp33_ASAP7_75t_L g2456 ( 
.A(n_2319),
.B(n_1918),
.Y(n_2456)
);

INVx2_ASAP7_75t_SL g2457 ( 
.A(n_2062),
.Y(n_2457)
);

INVx4_ASAP7_75t_L g2458 ( 
.A(n_2028),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2236),
.B(n_1938),
.Y(n_2459)
);

INVx2_ASAP7_75t_SL g2460 ( 
.A(n_2064),
.Y(n_2460)
);

INVx4_ASAP7_75t_L g2461 ( 
.A(n_2029),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2273),
.B(n_1931),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2129),
.B(n_2287),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2142),
.Y(n_2464)
);

INVx5_ASAP7_75t_L g2465 ( 
.A(n_2073),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2227),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2275),
.B(n_1931),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2148),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2231),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2153),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2155),
.Y(n_2471)
);

BUFx2_ASAP7_75t_L g2472 ( 
.A(n_2205),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2065),
.Y(n_2473)
);

INVx4_ASAP7_75t_L g2474 ( 
.A(n_2321),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2231),
.Y(n_2475)
);

AND2x6_ASAP7_75t_L g2476 ( 
.A(n_2287),
.B(n_1802),
.Y(n_2476)
);

INVx4_ASAP7_75t_SL g2477 ( 
.A(n_2034),
.Y(n_2477)
);

INVx2_ASAP7_75t_SL g2478 ( 
.A(n_2066),
.Y(n_2478)
);

NAND2xp33_ASAP7_75t_L g2479 ( 
.A(n_2196),
.B(n_1922),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2246),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2136),
.B(n_1922),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2269),
.B(n_1465),
.Y(n_2482)
);

INVxp67_ASAP7_75t_SL g2483 ( 
.A(n_2272),
.Y(n_2483)
);

OR2x2_ASAP7_75t_L g2484 ( 
.A(n_2228),
.B(n_1804),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2246),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2272),
.Y(n_2486)
);

NAND2xp33_ASAP7_75t_L g2487 ( 
.A(n_2197),
.B(n_1926),
.Y(n_2487)
);

OAI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2162),
.A2(n_2164),
.B1(n_2161),
.B2(n_2220),
.Y(n_2488)
);

BUFx10_ASAP7_75t_L g2489 ( 
.A(n_2014),
.Y(n_2489)
);

BUFx2_ASAP7_75t_L g2490 ( 
.A(n_2205),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2224),
.B(n_1465),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2224),
.B(n_1477),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2124),
.B(n_1227),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_SL g2494 ( 
.A(n_2067),
.B(n_1001),
.Y(n_2494)
);

BUFx10_ASAP7_75t_L g2495 ( 
.A(n_2033),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_2272),
.Y(n_2496)
);

NAND3xp33_ASAP7_75t_L g2497 ( 
.A(n_2150),
.B(n_1832),
.C(n_1826),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2139),
.B(n_1926),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_2272),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2159),
.Y(n_2500)
);

INVx3_ASAP7_75t_L g2501 ( 
.A(n_2286),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2160),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_2207),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2224),
.B(n_1477),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2170),
.Y(n_2505)
);

INVx6_ASAP7_75t_L g2506 ( 
.A(n_2265),
.Y(n_2506)
);

BUFx4f_ASAP7_75t_L g2507 ( 
.A(n_2243),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2294),
.B(n_1834),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2141),
.B(n_1926),
.Y(n_2509)
);

AOI22xp33_ASAP7_75t_L g2510 ( 
.A1(n_2294),
.A2(n_1032),
.B1(n_1300),
.B2(n_1836),
.Y(n_2510)
);

CKINVDCx20_ASAP7_75t_R g2511 ( 
.A(n_2005),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2236),
.B(n_1925),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2193),
.B(n_1486),
.Y(n_2513)
);

AOI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_2285),
.A2(n_1843),
.B1(n_1851),
.B2(n_1839),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2174),
.Y(n_2515)
);

INVx4_ASAP7_75t_L g2516 ( 
.A(n_2068),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2186),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_SL g2518 ( 
.A(n_2072),
.B(n_1858),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2055),
.B(n_1861),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2277),
.B(n_2278),
.Y(n_2520)
);

INVx1_ASAP7_75t_SL g2521 ( 
.A(n_2207),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2251),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2286),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2055),
.B(n_1872),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2143),
.B(n_1933),
.Y(n_2525)
);

AND3x2_ASAP7_75t_L g2526 ( 
.A(n_2179),
.B(n_1930),
.C(n_1103),
.Y(n_2526)
);

AND2x2_ASAP7_75t_SL g2527 ( 
.A(n_2292),
.B(n_2192),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2253),
.B(n_1486),
.Y(n_2528)
);

INVx4_ASAP7_75t_SL g2529 ( 
.A(n_2286),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2191),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_2075),
.Y(n_2531)
);

BUFx2_ASAP7_75t_L g2532 ( 
.A(n_2209),
.Y(n_2532)
);

BUFx3_ASAP7_75t_L g2533 ( 
.A(n_2147),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2201),
.Y(n_2534)
);

INVxp33_ASAP7_75t_L g2535 ( 
.A(n_2234),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2178),
.B(n_1875),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2299),
.Y(n_2537)
);

INVx1_ASAP7_75t_SL g2538 ( 
.A(n_2209),
.Y(n_2538)
);

INVxp67_ASAP7_75t_SL g2539 ( 
.A(n_2286),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_2151),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2211),
.B(n_1247),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2112),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2299),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2313),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2251),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2318),
.Y(n_2546)
);

OR2x6_ASAP7_75t_L g2547 ( 
.A(n_2238),
.B(n_1877),
.Y(n_2547)
);

BUFx3_ASAP7_75t_L g2548 ( 
.A(n_2152),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2247),
.B(n_2250),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2222),
.B(n_1247),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2093),
.B(n_2094),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2226),
.B(n_1274),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2318),
.Y(n_2553)
);

INVx3_ASAP7_75t_L g2554 ( 
.A(n_2313),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_2265),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2093),
.B(n_1887),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2144),
.B(n_1933),
.Y(n_2557)
);

INVx1_ASAP7_75t_SL g2558 ( 
.A(n_2112),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2165),
.B(n_1500),
.Y(n_2559)
);

BUFx3_ASAP7_75t_L g2560 ( 
.A(n_2156),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_2167),
.B(n_1933),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2168),
.B(n_1933),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2252),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2171),
.B(n_1889),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2212),
.B(n_1274),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2172),
.B(n_1892),
.Y(n_2566)
);

OR2x2_ASAP7_75t_L g2567 ( 
.A(n_2103),
.B(n_1897),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2173),
.B(n_1500),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_L g2569 ( 
.A1(n_2094),
.A2(n_1907),
.B1(n_1908),
.B2(n_1901),
.Y(n_2569)
);

NOR2x1p5_ASAP7_75t_L g2570 ( 
.A(n_2080),
.B(n_1909),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2225),
.Y(n_2571)
);

INVx4_ASAP7_75t_L g2572 ( 
.A(n_2254),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2100),
.A2(n_1941),
.B1(n_1085),
.B2(n_1087),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2229),
.B(n_1102),
.Y(n_2574)
);

INVx5_ASAP7_75t_L g2575 ( 
.A(n_2037),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2175),
.B(n_1502),
.Y(n_2576)
);

INVx6_ASAP7_75t_L g2577 ( 
.A(n_2243),
.Y(n_2577)
);

BUFx2_ASAP7_75t_L g2578 ( 
.A(n_2288),
.Y(n_2578)
);

INVx6_ASAP7_75t_L g2579 ( 
.A(n_2244),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_SL g2580 ( 
.A(n_2176),
.B(n_1860),
.Y(n_2580)
);

OR2x6_ASAP7_75t_L g2581 ( 
.A(n_2113),
.B(n_1723),
.Y(n_2581)
);

BUFx10_ASAP7_75t_L g2582 ( 
.A(n_2035),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2252),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2237),
.Y(n_2584)
);

BUFx2_ASAP7_75t_L g2585 ( 
.A(n_2256),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2180),
.B(n_2183),
.Y(n_2586)
);

AOI22xp33_ASAP7_75t_SL g2587 ( 
.A1(n_2131),
.A2(n_1521),
.B1(n_1535),
.B2(n_1502),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2263),
.Y(n_2588)
);

BUFx6f_ASAP7_75t_L g2589 ( 
.A(n_2245),
.Y(n_2589)
);

OAI22xp5_ASAP7_75t_L g2590 ( 
.A1(n_2218),
.A2(n_1884),
.B1(n_1879),
.B2(n_1728),
.Y(n_2590)
);

BUFx10_ASAP7_75t_L g2591 ( 
.A(n_2039),
.Y(n_2591)
);

NAND3xp33_ASAP7_75t_L g2592 ( 
.A(n_2199),
.B(n_1748),
.C(n_1738),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2239),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2257),
.B(n_1860),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2313),
.Y(n_2595)
);

NAND3xp33_ASAP7_75t_L g2596 ( 
.A(n_2271),
.B(n_1859),
.C(n_1857),
.Y(n_2596)
);

NOR2x1p5_ASAP7_75t_L g2597 ( 
.A(n_2051),
.B(n_1317),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_2291),
.B(n_1869),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2241),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2255),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_SL g2601 ( 
.A(n_2260),
.B(n_1869),
.Y(n_2601)
);

INVxp33_ASAP7_75t_L g2602 ( 
.A(n_2240),
.Y(n_2602)
);

INVx4_ASAP7_75t_L g2603 ( 
.A(n_2262),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2320),
.Y(n_2604)
);

AOI22xp33_ASAP7_75t_L g2605 ( 
.A1(n_2100),
.A2(n_1086),
.B1(n_1091),
.B2(n_1089),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2242),
.B(n_1883),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2305),
.B(n_1521),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2320),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_SL g2609 ( 
.A(n_2244),
.B(n_1883),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_2244),
.B(n_1535),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_L g2611 ( 
.A(n_2280),
.B(n_1540),
.Y(n_2611)
);

INVx4_ASAP7_75t_L g2612 ( 
.A(n_2056),
.Y(n_2612)
);

BUFx8_ASAP7_75t_SL g2613 ( 
.A(n_2036),
.Y(n_2613)
);

INVx5_ASAP7_75t_L g2614 ( 
.A(n_2037),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2270),
.Y(n_2615)
);

BUFx10_ASAP7_75t_L g2616 ( 
.A(n_2041),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2274),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2320),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2276),
.Y(n_2619)
);

NOR3xp33_ASAP7_75t_L g2620 ( 
.A(n_2235),
.B(n_1886),
.C(n_1349),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2289),
.B(n_1540),
.Y(n_2621)
);

AOI22xp33_ASAP7_75t_L g2622 ( 
.A1(n_2304),
.A2(n_1837),
.B1(n_1864),
.B2(n_1821),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2307),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2107),
.B(n_1886),
.Y(n_2624)
);

XOR2xp5_ASAP7_75t_L g2625 ( 
.A(n_2063),
.B(n_1558),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2157),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2311),
.Y(n_2627)
);

INVx2_ASAP7_75t_SL g2628 ( 
.A(n_2290),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2312),
.Y(n_2629)
);

AND2x4_ASAP7_75t_L g2630 ( 
.A(n_2314),
.B(n_1857),
.Y(n_2630)
);

INVx4_ASAP7_75t_L g2631 ( 
.A(n_2058),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2263),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2245),
.Y(n_2633)
);

BUFx6f_ASAP7_75t_L g2634 ( 
.A(n_2245),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2282),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2282),
.Y(n_2636)
);

BUFx3_ASAP7_75t_L g2637 ( 
.A(n_2054),
.Y(n_2637)
);

AOI22xp33_ASAP7_75t_L g2638 ( 
.A1(n_2302),
.A2(n_1837),
.B1(n_1864),
.B2(n_1821),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2010),
.Y(n_2639)
);

INVxp67_ASAP7_75t_SL g2640 ( 
.A(n_2107),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2293),
.B(n_1558),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2281),
.B(n_1898),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2010),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2011),
.Y(n_2644)
);

BUFx3_ASAP7_75t_L g2645 ( 
.A(n_2111),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2011),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2021),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2110),
.B(n_1799),
.Y(n_2648)
);

AND2x2_ASAP7_75t_SL g2649 ( 
.A(n_2102),
.B(n_1566),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2110),
.B(n_1799),
.Y(n_2650)
);

AOI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2098),
.A2(n_1794),
.B1(n_1815),
.B2(n_1821),
.Y(n_2651)
);

INVxp67_ASAP7_75t_L g2652 ( 
.A(n_2085),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2021),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2022),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2119),
.B(n_2258),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_2037),
.Y(n_2656)
);

AND2x2_ASAP7_75t_SL g2657 ( 
.A(n_2102),
.B(n_1566),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2105),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2022),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2045),
.Y(n_2660)
);

AND3x2_ASAP7_75t_L g2661 ( 
.A(n_2076),
.B(n_1319),
.C(n_1318),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2045),
.B(n_1803),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2046),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2046),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2049),
.Y(n_2665)
);

AND2x6_ASAP7_75t_L g2666 ( 
.A(n_2049),
.B(n_1859),
.Y(n_2666)
);

INVx4_ASAP7_75t_L g2667 ( 
.A(n_2106),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_2145),
.B(n_1864),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2086),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2306),
.A2(n_2188),
.B1(n_2185),
.B2(n_2190),
.Y(n_2670)
);

BUFx3_ASAP7_75t_L g2671 ( 
.A(n_2111),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_2108),
.Y(n_2672)
);

NAND2xp33_ASAP7_75t_SL g2673 ( 
.A(n_2267),
.B(n_1571),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2109),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2120),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2127),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2128),
.B(n_2132),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2133),
.B(n_1571),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2134),
.Y(n_2679)
);

OR2x2_ASAP7_75t_L g2680 ( 
.A(n_2146),
.B(n_1865),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2640),
.B(n_1794),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2486),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2331),
.B(n_1586),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2652),
.B(n_1815),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2652),
.B(n_1865),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2438),
.B(n_2203),
.Y(n_2686)
);

BUFx3_ASAP7_75t_L g2687 ( 
.A(n_2473),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_SL g2688 ( 
.A(n_2438),
.B(n_2216),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2325),
.Y(n_2689)
);

NAND2xp33_ASAP7_75t_L g2690 ( 
.A(n_2555),
.B(n_2200),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2640),
.B(n_1803),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2329),
.B(n_1811),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2537),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2329),
.B(n_1811),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2543),
.Y(n_2695)
);

NOR2xp67_ASAP7_75t_L g2696 ( 
.A(n_2372),
.B(n_2053),
.Y(n_2696)
);

AOI221x1_ASAP7_75t_L g2697 ( 
.A1(n_2620),
.A2(n_2447),
.B1(n_2590),
.B2(n_2655),
.C(n_2328),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2380),
.B(n_1775),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_2507),
.B(n_2283),
.Y(n_2699)
);

NAND3xp33_ASAP7_75t_L g2700 ( 
.A(n_2417),
.B(n_2023),
.C(n_2256),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2380),
.B(n_1867),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2328),
.B(n_1867),
.Y(n_2702)
);

BUFx6f_ASAP7_75t_L g2703 ( 
.A(n_2486),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2366),
.B(n_2131),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2493),
.B(n_2154),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2508),
.B(n_2519),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2334),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2507),
.B(n_2378),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2508),
.B(n_1871),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2519),
.B(n_1871),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2546),
.Y(n_2711)
);

INVxp33_ASAP7_75t_L g2712 ( 
.A(n_2559),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2486),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2524),
.B(n_1874),
.Y(n_2714)
);

INVxp33_ASAP7_75t_L g2715 ( 
.A(n_2568),
.Y(n_2715)
);

NOR3xp33_ASAP7_75t_L g2716 ( 
.A(n_2402),
.B(n_2048),
.C(n_2047),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2553),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2415),
.B(n_1586),
.Y(n_2718)
);

OR2x6_ASAP7_75t_L g2719 ( 
.A(n_2445),
.B(n_1874),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2383),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2339),
.B(n_1878),
.Y(n_2721)
);

OR2x6_ASAP7_75t_L g2722 ( 
.A(n_2448),
.B(n_1878),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2384),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2339),
.B(n_1882),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2378),
.B(n_2154),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_L g2726 ( 
.A(n_2488),
.B(n_1596),
.Y(n_2726)
);

INVx2_ASAP7_75t_SL g2727 ( 
.A(n_2348),
.Y(n_2727)
);

AOI22xp33_ASAP7_75t_L g2728 ( 
.A1(n_2371),
.A2(n_2184),
.B1(n_2158),
.B2(n_2117),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2385),
.Y(n_2729)
);

AOI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2371),
.A2(n_2184),
.B1(n_2158),
.B2(n_2117),
.Y(n_2730)
);

INVx2_ASAP7_75t_SL g2731 ( 
.A(n_2348),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2344),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2400),
.Y(n_2733)
);

A2O1A1Ixp33_ASAP7_75t_L g2734 ( 
.A1(n_2655),
.A2(n_2208),
.B(n_2206),
.C(n_1888),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2404),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2446),
.Y(n_2736)
);

BUFx3_ASAP7_75t_L g2737 ( 
.A(n_2637),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2377),
.B(n_1882),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2410),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_SL g2740 ( 
.A(n_2391),
.B(n_2189),
.Y(n_2740)
);

OAI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2670),
.A2(n_2130),
.B1(n_2076),
.B2(n_2087),
.Y(n_2741)
);

INVxp67_ASAP7_75t_SL g2742 ( 
.A(n_2355),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_SL g2743 ( 
.A(n_2391),
.B(n_2130),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2335),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2377),
.B(n_2397),
.Y(n_2745)
);

BUFx6f_ASAP7_75t_L g2746 ( 
.A(n_2555),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2397),
.B(n_1821),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2357),
.B(n_1888),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2347),
.Y(n_2749)
);

INVx2_ASAP7_75t_SL g2750 ( 
.A(n_2340),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_SL g2751 ( 
.A(n_2494),
.B(n_1837),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2353),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2411),
.Y(n_2753)
);

INVx1_ASAP7_75t_SL g2754 ( 
.A(n_2340),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2322),
.B(n_1890),
.Y(n_2755)
);

INVxp67_ASAP7_75t_SL g2756 ( 
.A(n_2355),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2357),
.B(n_1890),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2488),
.B(n_1596),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2368),
.Y(n_2759)
);

AOI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2443),
.A2(n_2087),
.B1(n_2089),
.B2(n_2082),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2586),
.B(n_2494),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2414),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2623),
.B(n_1837),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_SL g2764 ( 
.A(n_2518),
.B(n_1864),
.Y(n_2764)
);

NOR2x1p5_ASAP7_75t_L g2765 ( 
.A(n_2337),
.B(n_2097),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_L g2766 ( 
.A(n_2424),
.B(n_1607),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2524),
.B(n_1866),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2555),
.Y(n_2768)
);

INVx2_ASAP7_75t_SL g2769 ( 
.A(n_2330),
.Y(n_2769)
);

AND2x4_ASAP7_75t_L g2770 ( 
.A(n_2322),
.B(n_1866),
.Y(n_2770)
);

BUFx8_ASAP7_75t_L g2771 ( 
.A(n_2338),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2396),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2627),
.B(n_1866),
.Y(n_2773)
);

NAND3xp33_ASAP7_75t_SL g2774 ( 
.A(n_2620),
.B(n_1622),
.C(n_1607),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2362),
.B(n_1622),
.Y(n_2775)
);

INVxp67_ASAP7_75t_L g2776 ( 
.A(n_2330),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2629),
.B(n_1866),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_2528),
.B(n_1636),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2341),
.B(n_1868),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2403),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2406),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2518),
.B(n_1868),
.Y(n_2782)
);

NAND2xp33_ASAP7_75t_L g2783 ( 
.A(n_2531),
.B(n_2096),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_2452),
.B(n_2459),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2590),
.B(n_1868),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2513),
.B(n_1636),
.Y(n_2786)
);

BUFx8_ASAP7_75t_L g2787 ( 
.A(n_2379),
.Y(n_2787)
);

NOR3xp33_ASAP7_75t_L g2788 ( 
.A(n_2389),
.B(n_2249),
.C(n_2101),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2416),
.B(n_1868),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2440),
.A2(n_2089),
.B1(n_2082),
.B2(n_2095),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2427),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2405),
.B(n_2009),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_2369),
.B(n_2399),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2452),
.B(n_1880),
.Y(n_2794)
);

NOR3xp33_ASAP7_75t_L g2795 ( 
.A(n_2611),
.B(n_1322),
.C(n_1321),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2435),
.Y(n_2796)
);

INVxp67_ASAP7_75t_L g2797 ( 
.A(n_2574),
.Y(n_2797)
);

NAND3xp33_ASAP7_75t_L g2798 ( 
.A(n_2576),
.B(n_2482),
.C(n_2520),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2390),
.B(n_1641),
.Y(n_2799)
);

INVxp33_ASAP7_75t_L g2800 ( 
.A(n_2621),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2444),
.Y(n_2801)
);

BUFx12f_ASAP7_75t_SL g2802 ( 
.A(n_2337),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2556),
.B(n_1880),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2556),
.B(n_1880),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2407),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2408),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2352),
.B(n_1880),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2413),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2352),
.B(n_1898),
.Y(n_2809)
);

OAI221xp5_ASAP7_75t_L g2810 ( 
.A1(n_2374),
.A2(n_997),
.B1(n_999),
.B2(n_996),
.C(n_995),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2463),
.B(n_1898),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_2390),
.B(n_1641),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2680),
.B(n_1898),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_SL g2814 ( 
.A(n_2474),
.B(n_1900),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2535),
.B(n_2602),
.Y(n_2815)
);

AOI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2577),
.A2(n_2095),
.B1(n_1645),
.B2(n_1649),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2677),
.B(n_1644),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2455),
.B(n_1900),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2381),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2464),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2468),
.Y(n_2821)
);

OAI22xp33_ASAP7_75t_L g2822 ( 
.A1(n_2567),
.A2(n_1649),
.B1(n_1690),
.B2(n_1663),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2470),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2431),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2466),
.Y(n_2825)
);

NAND2xp33_ASAP7_75t_L g2826 ( 
.A(n_2412),
.B(n_2336),
.Y(n_2826)
);

BUFx3_ASAP7_75t_L g2827 ( 
.A(n_2342),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2469),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2475),
.Y(n_2829)
);

INVxp67_ASAP7_75t_L g2830 ( 
.A(n_2381),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_SL g2831 ( 
.A(n_2474),
.B(n_1900),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2549),
.B(n_1645),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2471),
.B(n_1900),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_2457),
.B(n_1663),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2500),
.B(n_1740),
.Y(n_2835)
);

AOI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_2630),
.A2(n_1741),
.B1(n_1750),
.B2(n_1740),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2577),
.A2(n_1690),
.B1(n_2063),
.B2(n_1798),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2502),
.B(n_1741),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2505),
.B(n_1750),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2480),
.Y(n_2840)
);

NAND3xp33_ASAP7_75t_SL g2841 ( 
.A(n_2374),
.B(n_2187),
.C(n_1004),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2485),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2522),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2545),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2515),
.B(n_1769),
.Y(n_2845)
);

AOI22x1_ASAP7_75t_L g2846 ( 
.A1(n_2669),
.A2(n_1778),
.B1(n_1769),
.B2(n_1797),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2463),
.B(n_1778),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2517),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2551),
.B(n_1761),
.Y(n_2849)
);

INVxp67_ASAP7_75t_L g2850 ( 
.A(n_2394),
.Y(n_2850)
);

OR2x2_ASAP7_75t_L g2851 ( 
.A(n_2521),
.B(n_1320),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_2460),
.B(n_1797),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_SL g2853 ( 
.A(n_2478),
.B(n_1797),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2530),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2563),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2583),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2551),
.B(n_2624),
.Y(n_2857)
);

BUFx6f_ASAP7_75t_L g2858 ( 
.A(n_2336),
.Y(n_2858)
);

OAI22xp33_ASAP7_75t_L g2859 ( 
.A1(n_2536),
.A2(n_2187),
.B1(n_1005),
.B2(n_1008),
.Y(n_2859)
);

AOI221xp5_ASAP7_75t_L g2860 ( 
.A1(n_2440),
.A2(n_1012),
.B1(n_1013),
.B2(n_1010),
.C(n_1000),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2598),
.B(n_1797),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2588),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2632),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2624),
.B(n_1761),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2550),
.B(n_1129),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2569),
.B(n_1761),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2351),
.B(n_1798),
.Y(n_2867)
);

INVxp33_ASAP7_75t_L g2868 ( 
.A(n_2641),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2639),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2569),
.B(n_1761),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2534),
.B(n_1764),
.Y(n_2871)
);

AOI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2577),
.A2(n_1798),
.B1(n_1801),
.B2(n_1789),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2333),
.B(n_1764),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2336),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2643),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2598),
.B(n_1798),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2346),
.B(n_1764),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2350),
.B(n_1764),
.Y(n_2878)
);

BUFx6f_ASAP7_75t_L g2879 ( 
.A(n_2392),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2351),
.B(n_1801),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2647),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2653),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2359),
.B(n_1801),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2356),
.B(n_1770),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2664),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2364),
.Y(n_2886)
);

OAI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2386),
.A2(n_1733),
.B(n_1715),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2343),
.B(n_1770),
.Y(n_2888)
);

AOI221xp5_ASAP7_75t_L g2889 ( 
.A1(n_2361),
.A2(n_1019),
.B1(n_1020),
.B2(n_1018),
.C(n_1017),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2373),
.B(n_1770),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2459),
.B(n_1801),
.Y(n_2891)
);

INVxp67_ASAP7_75t_L g2892 ( 
.A(n_2484),
.Y(n_2892)
);

AOI22x1_ASAP7_75t_L g2893 ( 
.A1(n_2544),
.A2(n_1789),
.B1(n_1733),
.B2(n_1715),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2544),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2571),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2343),
.B(n_1770),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2554),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2552),
.B(n_1152),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2359),
.B(n_1771),
.Y(n_2899)
);

NOR3xp33_ASAP7_75t_L g2900 ( 
.A(n_2678),
.B(n_1023),
.C(n_1022),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2554),
.B(n_1771),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2630),
.B(n_1771),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2595),
.B(n_1771),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2584),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2593),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_SL g2906 ( 
.A(n_2367),
.B(n_1027),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2599),
.Y(n_2907)
);

NAND2xp33_ASAP7_75t_R g2908 ( 
.A(n_2607),
.B(n_657),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2510),
.B(n_1784),
.Y(n_2909)
);

AND2x4_ASAP7_75t_L g2910 ( 
.A(n_2512),
.B(n_1784),
.Y(n_2910)
);

BUFx6f_ASAP7_75t_L g2911 ( 
.A(n_2392),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2512),
.B(n_1784),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2510),
.B(n_1784),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2595),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_L g2915 ( 
.A(n_2367),
.B(n_1789),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2604),
.Y(n_2916)
);

INVx2_ASAP7_75t_SL g2917 ( 
.A(n_2451),
.Y(n_2917)
);

OAI22xp33_ASAP7_75t_L g2918 ( 
.A1(n_2360),
.A2(n_1030),
.B1(n_1031),
.B2(n_1028),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2604),
.B(n_1789),
.Y(n_2919)
);

OAI22xp33_ASAP7_75t_L g2920 ( 
.A1(n_2437),
.A2(n_1036),
.B1(n_1035),
.B2(n_1152),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2361),
.B(n_1153),
.Y(n_2921)
);

BUFx6f_ASAP7_75t_L g2922 ( 
.A(n_2392),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2514),
.B(n_1153),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2600),
.B(n_1847),
.Y(n_2924)
);

INVxp67_ASAP7_75t_L g2925 ( 
.A(n_2565),
.Y(n_2925)
);

NAND2xp33_ASAP7_75t_L g2926 ( 
.A(n_2454),
.B(n_1730),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2615),
.B(n_2617),
.Y(n_2927)
);

CKINVDCx11_ASAP7_75t_R g2928 ( 
.A(n_2332),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2608),
.Y(n_2929)
);

AOI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2327),
.A2(n_1731),
.B1(n_1739),
.B2(n_1730),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2619),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2573),
.B(n_1847),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2608),
.Y(n_2933)
);

NOR3xp33_ASAP7_75t_L g2934 ( 
.A(n_2587),
.B(n_1323),
.C(n_1320),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_SL g2935 ( 
.A(n_2454),
.B(n_2393),
.Y(n_2935)
);

INVx3_ASAP7_75t_L g2936 ( 
.A(n_2618),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2644),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2646),
.Y(n_2938)
);

INVxp67_ASAP7_75t_L g2939 ( 
.A(n_2425),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2654),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2573),
.B(n_1847),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2421),
.B(n_1847),
.Y(n_2942)
);

NOR2xp33_ASAP7_75t_L g2943 ( 
.A(n_2393),
.B(n_1731),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2618),
.Y(n_2944)
);

INVxp67_ASAP7_75t_L g2945 ( 
.A(n_2442),
.Y(n_2945)
);

OAI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2386),
.A2(n_1095),
.B(n_1094),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2659),
.Y(n_2947)
);

INVxp67_ASAP7_75t_L g2948 ( 
.A(n_2472),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2454),
.B(n_1730),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2660),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_2458),
.B(n_1730),
.Y(n_2951)
);

BUFx6f_ASAP7_75t_SL g2952 ( 
.A(n_2495),
.Y(n_2952)
);

INVx2_ASAP7_75t_SL g2953 ( 
.A(n_2349),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2421),
.B(n_1731),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2458),
.B(n_1739),
.Y(n_2955)
);

OAI21xp33_ASAP7_75t_L g2956 ( 
.A1(n_2587),
.A2(n_1323),
.B(n_1303),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2663),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_SL g2958 ( 
.A(n_2461),
.B(n_1739),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2665),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2387),
.B(n_1096),
.Y(n_2960)
);

NOR2xp33_ASAP7_75t_L g2961 ( 
.A(n_2461),
.B(n_1739),
.Y(n_2961)
);

BUFx5_ASAP7_75t_L g2962 ( 
.A(n_2666),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2387),
.B(n_1078),
.Y(n_2963)
);

AOI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2596),
.A2(n_1752),
.B1(n_1759),
.B2(n_1747),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2516),
.B(n_1747),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2450),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2516),
.B(n_1747),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_SL g2968 ( 
.A(n_2572),
.B(n_1285),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_2521),
.B(n_1747),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2635),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_2349),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2450),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2675),
.B(n_1752),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2538),
.B(n_2542),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2483),
.B(n_1752),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2450),
.Y(n_2976)
);

INVx1_ASAP7_75t_SL g2977 ( 
.A(n_2754),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2793),
.B(n_2538),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2745),
.B(n_2481),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2720),
.Y(n_2980)
);

INVxp33_ASAP7_75t_SL g2981 ( 
.A(n_2817),
.Y(n_2981)
);

AND2x2_ASAP7_75t_SL g2982 ( 
.A(n_2726),
.B(n_2649),
.Y(n_2982)
);

AO22x2_ASAP7_75t_L g2983 ( 
.A1(n_2697),
.A2(n_2558),
.B1(n_2542),
.B2(n_2592),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_L g2984 ( 
.A(n_2712),
.B(n_2558),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2886),
.Y(n_2985)
);

NAND2x1p5_ASAP7_75t_L g2986 ( 
.A(n_2736),
.B(n_2533),
.Y(n_2986)
);

AND2x4_ASAP7_75t_L g2987 ( 
.A(n_2737),
.B(n_2570),
.Y(n_2987)
);

NAND2xp33_ASAP7_75t_L g2988 ( 
.A(n_2746),
.B(n_2345),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2723),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2729),
.Y(n_2990)
);

INVxp67_ASAP7_75t_L g2991 ( 
.A(n_2974),
.Y(n_2991)
);

INVxp67_ASAP7_75t_L g2992 ( 
.A(n_2750),
.Y(n_2992)
);

BUFx2_ASAP7_75t_L g2993 ( 
.A(n_2754),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2733),
.Y(n_2994)
);

AO22x2_ASAP7_75t_L g2995 ( 
.A1(n_2790),
.A2(n_2420),
.B1(n_2477),
.B2(n_2401),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2735),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2715),
.B(n_2610),
.Y(n_2997)
);

CKINVDCx5p33_ASAP7_75t_R g2998 ( 
.A(n_2928),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2952),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2739),
.Y(n_3000)
);

AO22x2_ASAP7_75t_L g3001 ( 
.A1(n_2790),
.A2(n_2420),
.B1(n_2477),
.B2(n_2401),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2863),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2800),
.B(n_2491),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2753),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2762),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2947),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2791),
.Y(n_3007)
);

OAI221xp5_ASAP7_75t_L g3008 ( 
.A1(n_2766),
.A2(n_2673),
.B1(n_2504),
.B2(n_2492),
.C(n_2566),
.Y(n_3008)
);

OAI221xp5_ASAP7_75t_L g3009 ( 
.A1(n_2683),
.A2(n_2564),
.B1(n_2658),
.B2(n_2497),
.C(n_2449),
.Y(n_3009)
);

CKINVDCx5p33_ASAP7_75t_R g3010 ( 
.A(n_2952),
.Y(n_3010)
);

BUFx2_ASAP7_75t_L g3011 ( 
.A(n_2939),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2796),
.Y(n_3012)
);

NAND3xp33_ASAP7_75t_SL g3013 ( 
.A(n_2760),
.B(n_2900),
.C(n_2718),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2801),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2820),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2950),
.Y(n_3016)
);

AO22x2_ASAP7_75t_L g3017 ( 
.A1(n_2841),
.A2(n_2420),
.B1(n_2477),
.B2(n_2401),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2725),
.A2(n_2547),
.B1(n_2657),
.B2(n_2541),
.Y(n_3018)
);

AO22x2_ASAP7_75t_L g3019 ( 
.A1(n_2774),
.A2(n_2609),
.B1(n_2509),
.B2(n_2525),
.Y(n_3019)
);

BUFx3_ASAP7_75t_L g3020 ( 
.A(n_2687),
.Y(n_3020)
);

OAI221xp5_ASAP7_75t_L g3021 ( 
.A1(n_2761),
.A2(n_2786),
.B1(n_2797),
.B2(n_2758),
.C(n_2778),
.Y(n_3021)
);

AO22x2_ASAP7_75t_L g3022 ( 
.A1(n_2743),
.A2(n_2557),
.B1(n_2561),
.B2(n_2498),
.Y(n_3022)
);

NOR3xp33_ASAP7_75t_L g3023 ( 
.A(n_2798),
.B(n_2578),
.C(n_2668),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2957),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2821),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2823),
.Y(n_3026)
);

INVxp67_ASAP7_75t_L g3027 ( 
.A(n_2704),
.Y(n_3027)
);

INVx2_ASAP7_75t_SL g3028 ( 
.A(n_2744),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2848),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2854),
.Y(n_3030)
);

AND2x6_ASAP7_75t_L g3031 ( 
.A(n_2897),
.B(n_2651),
.Y(n_3031)
);

AO22x2_ASAP7_75t_L g3032 ( 
.A1(n_2700),
.A2(n_2562),
.B1(n_2625),
.B2(n_2674),
.Y(n_3032)
);

AO22x2_ASAP7_75t_L g3033 ( 
.A1(n_2785),
.A2(n_2676),
.B1(n_2580),
.B2(n_2426),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2937),
.Y(n_3034)
);

NOR2xp67_ASAP7_75t_L g3035 ( 
.A(n_2850),
.B(n_2612),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2721),
.B(n_2679),
.Y(n_3036)
);

AO22x2_ASAP7_75t_L g3037 ( 
.A1(n_2751),
.A2(n_2462),
.B1(n_2467),
.B2(n_2419),
.Y(n_3037)
);

AND2x4_ASAP7_75t_L g3038 ( 
.A(n_2827),
.B(n_2540),
.Y(n_3038)
);

AOI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2775),
.A2(n_2418),
.B1(n_2511),
.B2(n_2628),
.Y(n_3039)
);

NAND2x1_ASAP7_75t_L g3040 ( 
.A(n_2897),
.B(n_2354),
.Y(n_3040)
);

AO22x2_ASAP7_75t_L g3041 ( 
.A1(n_2764),
.A2(n_2636),
.B1(n_2633),
.B2(n_2612),
.Y(n_3041)
);

INVxp67_ASAP7_75t_L g3042 ( 
.A(n_2769),
.Y(n_3042)
);

AO22x2_ASAP7_75t_L g3043 ( 
.A1(n_2782),
.A2(n_2631),
.B1(n_2672),
.B2(n_2667),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2938),
.Y(n_3044)
);

AOI22xp5_ASAP7_75t_L g3045 ( 
.A1(n_2799),
.A2(n_2812),
.B1(n_2834),
.B2(n_2832),
.Y(n_3045)
);

NAND2x1_ASAP7_75t_L g3046 ( 
.A(n_2936),
.B(n_2354),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2895),
.Y(n_3047)
);

OR2x6_ASAP7_75t_L g3048 ( 
.A(n_2727),
.B(n_2572),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2940),
.Y(n_3049)
);

BUFx8_ASAP7_75t_L g3050 ( 
.A(n_2731),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2959),
.Y(n_3051)
);

AO22x2_ASAP7_75t_L g3052 ( 
.A1(n_2966),
.A2(n_2631),
.B1(n_2672),
.B2(n_2667),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2917),
.B(n_2868),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2904),
.Y(n_3054)
);

OAI221xp5_ASAP7_75t_L g3055 ( 
.A1(n_2860),
.A2(n_2547),
.B1(n_2585),
.B2(n_2606),
.C(n_2503),
.Y(n_3055)
);

CKINVDCx5p33_ASAP7_75t_R g3056 ( 
.A(n_2802),
.Y(n_3056)
);

BUFx8_ASAP7_75t_L g3057 ( 
.A(n_2705),
.Y(n_3057)
);

OAI221xp5_ASAP7_75t_L g3058 ( 
.A1(n_2728),
.A2(n_2547),
.B1(n_2532),
.B2(n_2490),
.C(n_2581),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2724),
.B(n_2594),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2822),
.B(n_2815),
.Y(n_3060)
);

INVx2_ASAP7_75t_SL g3061 ( 
.A(n_2858),
.Y(n_3061)
);

AND2x4_ASAP7_75t_L g3062 ( 
.A(n_2784),
.B(n_2548),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2905),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2907),
.Y(n_3064)
);

NOR2xp67_ASAP7_75t_L g3065 ( 
.A(n_2696),
.B(n_2603),
.Y(n_3065)
);

AND2x4_ASAP7_75t_L g3066 ( 
.A(n_2784),
.B(n_2560),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2931),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2741),
.B(n_2730),
.Y(n_3068)
);

HB1xp67_ASAP7_75t_L g3069 ( 
.A(n_2776),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2927),
.Y(n_3070)
);

AO22x2_ASAP7_75t_L g3071 ( 
.A1(n_2972),
.A2(n_2976),
.B1(n_2708),
.B2(n_2921),
.Y(n_3071)
);

AND2x4_ASAP7_75t_L g3072 ( 
.A(n_2953),
.B(n_2626),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2693),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2738),
.B(n_2601),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2695),
.Y(n_3075)
);

BUFx3_ASAP7_75t_L g3076 ( 
.A(n_2771),
.Y(n_3076)
);

OR2x2_ASAP7_75t_SL g3077 ( 
.A(n_2851),
.B(n_2579),
.Y(n_3077)
);

BUFx2_ASAP7_75t_L g3078 ( 
.A(n_2945),
.Y(n_3078)
);

AND2x2_ASAP7_75t_L g3079 ( 
.A(n_2865),
.B(n_2603),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2711),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2717),
.Y(n_3081)
);

AND2x4_ASAP7_75t_L g3082 ( 
.A(n_2971),
.B(n_2645),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2869),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2875),
.Y(n_3084)
);

AO22x2_ASAP7_75t_L g3085 ( 
.A1(n_2740),
.A2(n_2671),
.B1(n_2526),
.B2(n_2539),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2898),
.B(n_2349),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2881),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2706),
.B(n_2527),
.Y(n_3088)
);

OR2x2_ASAP7_75t_L g3089 ( 
.A(n_2892),
.B(n_2948),
.Y(n_3089)
);

BUFx8_ASAP7_75t_L g3090 ( 
.A(n_2792),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2882),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2885),
.Y(n_3092)
);

AO22x2_ASAP7_75t_L g3093 ( 
.A1(n_2970),
.A2(n_2526),
.B1(n_2539),
.B2(n_2483),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2689),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2707),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2732),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2749),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2752),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2759),
.Y(n_3099)
);

NOR3xp33_ASAP7_75t_SL g3100 ( 
.A(n_2908),
.B(n_2859),
.C(n_2918),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2772),
.Y(n_3101)
);

AO22x2_ASAP7_75t_L g3102 ( 
.A1(n_2747),
.A2(n_2656),
.B1(n_2429),
.B2(n_2662),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2780),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2706),
.B(n_2422),
.Y(n_3104)
);

AOI22xp5_ASAP7_75t_SL g3105 ( 
.A1(n_2925),
.A2(n_2365),
.B1(n_2395),
.B2(n_2661),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2685),
.B(n_2428),
.Y(n_3106)
);

NOR2xp33_ASAP7_75t_L g3107 ( 
.A(n_2819),
.B(n_2579),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2781),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2684),
.B(n_2456),
.Y(n_3109)
);

AO22x2_ASAP7_75t_L g3110 ( 
.A1(n_2934),
.A2(n_2656),
.B1(n_2662),
.B2(n_2642),
.Y(n_3110)
);

AO22x2_ASAP7_75t_L g3111 ( 
.A1(n_2779),
.A2(n_2441),
.B1(n_2453),
.B2(n_2432),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2805),
.Y(n_3112)
);

AO22x2_ASAP7_75t_L g3113 ( 
.A1(n_2813),
.A2(n_2441),
.B1(n_2453),
.B2(n_2432),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2806),
.Y(n_3114)
);

AO22x2_ASAP7_75t_L g3115 ( 
.A1(n_2686),
.A2(n_2529),
.B1(n_2650),
.B2(n_2648),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2808),
.Y(n_3116)
);

AO22x2_ASAP7_75t_L g3117 ( 
.A1(n_2688),
.A2(n_2529),
.B1(n_2650),
.B2(n_2648),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2748),
.B(n_2579),
.Y(n_3118)
);

AO22x2_ASAP7_75t_L g3119 ( 
.A1(n_2742),
.A2(n_2529),
.B1(n_2581),
.B2(n_2376),
.Y(n_3119)
);

AO22x2_ASAP7_75t_L g3120 ( 
.A1(n_2756),
.A2(n_2581),
.B1(n_2376),
.B2(n_2496),
.Y(n_3120)
);

BUFx3_ASAP7_75t_L g3121 ( 
.A(n_2771),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2824),
.Y(n_3122)
);

INVxp67_ASAP7_75t_L g3123 ( 
.A(n_2830),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2825),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2858),
.Y(n_3125)
);

BUFx8_ASAP7_75t_L g3126 ( 
.A(n_2858),
.Y(n_3126)
);

OAI221xp5_ASAP7_75t_L g3127 ( 
.A1(n_2889),
.A2(n_2430),
.B1(n_2324),
.B2(n_2638),
.C(n_2622),
.Y(n_3127)
);

INVx3_ASAP7_75t_L g3128 ( 
.A(n_2874),
.Y(n_3128)
);

AOI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2968),
.A2(n_2433),
.B1(n_2495),
.B2(n_2582),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2828),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2837),
.B(n_2582),
.Y(n_3131)
);

AO22x2_ASAP7_75t_L g3132 ( 
.A1(n_2923),
.A2(n_2388),
.B1(n_2499),
.B2(n_2496),
.Y(n_3132)
);

AO22x2_ASAP7_75t_L g3133 ( 
.A1(n_2909),
.A2(n_2388),
.B1(n_2501),
.B2(n_2499),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2829),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2840),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2757),
.B(n_2605),
.Y(n_3136)
);

OAI22xp5_ASAP7_75t_SL g3137 ( 
.A1(n_2816),
.A2(n_2506),
.B1(n_2358),
.B2(n_2661),
.Y(n_3137)
);

BUFx8_ASAP7_75t_L g3138 ( 
.A(n_2874),
.Y(n_3138)
);

NAND2x1p5_ASAP7_75t_L g3139 ( 
.A(n_2746),
.B(n_2398),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2709),
.B(n_2605),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2709),
.B(n_2430),
.Y(n_3141)
);

AO22x2_ASAP7_75t_L g3142 ( 
.A1(n_2913),
.A2(n_2501),
.B1(n_2523),
.B2(n_2370),
.Y(n_3142)
);

AO22x2_ASAP7_75t_L g3143 ( 
.A1(n_2788),
.A2(n_2523),
.B1(n_2370),
.B2(n_2375),
.Y(n_3143)
);

AO22x2_ASAP7_75t_L g3144 ( 
.A1(n_2699),
.A2(n_2375),
.B1(n_2476),
.B2(n_1302),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2842),
.Y(n_3145)
);

AO22x2_ASAP7_75t_L g3146 ( 
.A1(n_2866),
.A2(n_2476),
.B1(n_1305),
.B2(n_1309),
.Y(n_3146)
);

OAI221xp5_ASAP7_75t_L g3147 ( 
.A1(n_2810),
.A2(n_2326),
.B1(n_2436),
.B2(n_2423),
.C(n_2382),
.Y(n_3147)
);

AO22x2_ASAP7_75t_L g3148 ( 
.A1(n_2866),
.A2(n_2476),
.B1(n_1308),
.B2(n_1314),
.Y(n_3148)
);

INVxp67_ASAP7_75t_L g3149 ( 
.A(n_2787),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2843),
.Y(n_3150)
);

AOI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_2968),
.A2(n_2597),
.B1(n_2382),
.B2(n_2506),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2844),
.Y(n_3152)
);

AOI22xp5_ASAP7_75t_SL g3153 ( 
.A1(n_2755),
.A2(n_2476),
.B1(n_2439),
.B2(n_2666),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2710),
.B(n_2358),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2855),
.Y(n_3155)
);

INVxp67_ASAP7_75t_L g3156 ( 
.A(n_2787),
.Y(n_3156)
);

AO22x2_ASAP7_75t_L g3157 ( 
.A1(n_2870),
.A2(n_2476),
.B1(n_1313),
.B2(n_2326),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2856),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2862),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2835),
.Y(n_3160)
);

AO22x2_ASAP7_75t_L g3161 ( 
.A1(n_2870),
.A2(n_1285),
.B1(n_2439),
.B2(n_2489),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2838),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_2906),
.B(n_2613),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2710),
.B(n_2358),
.Y(n_3164)
);

INVx2_ASAP7_75t_SL g3165 ( 
.A(n_2874),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2714),
.B(n_2506),
.Y(n_3166)
);

OR2x6_ASAP7_75t_L g3167 ( 
.A(n_2746),
.B(n_2323),
.Y(n_3167)
);

AO22x2_ASAP7_75t_L g3168 ( 
.A1(n_2852),
.A2(n_2439),
.B1(n_2489),
.B2(n_2363),
.Y(n_3168)
);

OA22x2_ASAP7_75t_L g3169 ( 
.A1(n_2719),
.A2(n_2591),
.B1(n_2616),
.B2(n_1252),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2839),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2845),
.Y(n_3171)
);

AO22x2_ASAP7_75t_L g3172 ( 
.A1(n_2853),
.A2(n_2439),
.B1(n_2666),
.B2(n_9),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2714),
.B(n_2479),
.Y(n_3173)
);

AO22x2_ASAP7_75t_L g3174 ( 
.A1(n_2973),
.A2(n_2439),
.B1(n_2666),
.B2(n_10),
.Y(n_3174)
);

OAI221xp5_ASAP7_75t_L g3175 ( 
.A1(n_2956),
.A2(n_2487),
.B1(n_2323),
.B2(n_2434),
.C(n_1252),
.Y(n_3175)
);

OAI221xp5_ASAP7_75t_L g3176 ( 
.A1(n_2795),
.A2(n_2434),
.B1(n_1252),
.B2(n_2616),
.C(n_2591),
.Y(n_3176)
);

OAI221xp5_ASAP7_75t_L g3177 ( 
.A1(n_2716),
.A2(n_2589),
.B1(n_2634),
.B2(n_1242),
.C(n_1219),
.Y(n_3177)
);

AO22x2_ASAP7_75t_L g3178 ( 
.A1(n_2701),
.A2(n_2666),
.B1(n_10),
.B2(n_6),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2894),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_R g3180 ( 
.A(n_2826),
.B(n_2398),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2755),
.B(n_1242),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_2879),
.Y(n_3182)
);

NAND2x1p5_ASAP7_75t_L g3183 ( 
.A(n_2768),
.B(n_2398),
.Y(n_3183)
);

CKINVDCx5p33_ASAP7_75t_R g3184 ( 
.A(n_2765),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2914),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2916),
.Y(n_3186)
);

OAI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_2681),
.A2(n_2409),
.B1(n_2465),
.B2(n_2398),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2701),
.B(n_2589),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2929),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2933),
.Y(n_3190)
);

INVxp67_ASAP7_75t_L g3191 ( 
.A(n_2969),
.Y(n_3191)
);

AOI22xp5_ASAP7_75t_L g3192 ( 
.A1(n_2906),
.A2(n_2794),
.B1(n_2783),
.B2(n_2770),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2944),
.Y(n_3193)
);

AOI22xp5_ASAP7_75t_L g3194 ( 
.A1(n_2794),
.A2(n_2465),
.B1(n_2409),
.B2(n_2589),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2847),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2770),
.B(n_2634),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2936),
.Y(n_3197)
);

AO22x2_ASAP7_75t_L g3198 ( 
.A1(n_2814),
.A2(n_2831),
.B1(n_2809),
.B2(n_2807),
.Y(n_3198)
);

AO22x2_ASAP7_75t_L g3199 ( 
.A1(n_2807),
.A2(n_2809),
.B1(n_2803),
.B2(n_2804),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_L g3200 ( 
.A(n_2920),
.B(n_2634),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2847),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2763),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2773),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_3047),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3070),
.B(n_2978),
.Y(n_3205)
);

AOI21xp5_ASAP7_75t_L g3206 ( 
.A1(n_3104),
.A2(n_2691),
.B(n_2767),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2979),
.B(n_2910),
.Y(n_3207)
);

O2A1O1Ixp33_ASAP7_75t_L g3208 ( 
.A1(n_3068),
.A2(n_2734),
.B(n_2935),
.C(n_2951),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_3177),
.A2(n_3173),
.B(n_3140),
.Y(n_3209)
);

BUFx4f_ASAP7_75t_L g3210 ( 
.A(n_2986),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3136),
.A2(n_2691),
.B(n_2767),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2991),
.B(n_3036),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2985),
.Y(n_3213)
);

OAI21x1_ASAP7_75t_L g3214 ( 
.A1(n_3188),
.A2(n_2846),
.B(n_2887),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_3160),
.B(n_2910),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_3147),
.A2(n_2804),
.B(n_2803),
.Y(n_3216)
);

NAND3xp33_ASAP7_75t_L g3217 ( 
.A(n_3100),
.B(n_2722),
.C(n_2719),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3162),
.B(n_2867),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_3106),
.A2(n_2614),
.B(n_2575),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3027),
.B(n_2719),
.Y(n_3220)
);

A2O1A1Ixp33_ASAP7_75t_L g3221 ( 
.A1(n_3008),
.A2(n_2880),
.B(n_2915),
.C(n_2883),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_3021),
.A2(n_3045),
.B1(n_2981),
.B2(n_3060),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3170),
.B(n_2879),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_3195),
.A2(n_2614),
.B(n_2575),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_3002),
.Y(n_3225)
);

A2O1A1Ixp33_ASAP7_75t_L g3226 ( 
.A1(n_3200),
.A2(n_3013),
.B(n_3009),
.C(n_3088),
.Y(n_3226)
);

AOI21xp5_ASAP7_75t_L g3227 ( 
.A1(n_3201),
.A2(n_2614),
.B(n_2575),
.Y(n_3227)
);

A2O1A1Ixp33_ASAP7_75t_L g3228 ( 
.A1(n_3141),
.A2(n_2943),
.B(n_2899),
.C(n_2961),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2980),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_3111),
.A2(n_2614),
.B(n_2575),
.Y(n_3230)
);

AOI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_3111),
.A2(n_2926),
.B(n_2857),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3171),
.B(n_2879),
.Y(n_3232)
);

INVx1_ASAP7_75t_SL g3233 ( 
.A(n_2977),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3018),
.A2(n_2722),
.B1(n_2681),
.B2(n_2965),
.Y(n_3234)
);

OAI21x1_ASAP7_75t_L g3235 ( 
.A1(n_3154),
.A2(n_2887),
.B(n_2893),
.Y(n_3235)
);

BUFx8_ASAP7_75t_SL g3236 ( 
.A(n_2998),
.Y(n_3236)
);

INVxp67_ASAP7_75t_SL g3237 ( 
.A(n_3069),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_SL g3238 ( 
.A(n_2997),
.B(n_2768),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_SL g3239 ( 
.A(n_3003),
.B(n_2768),
.Y(n_3239)
);

CKINVDCx10_ASAP7_75t_R g3240 ( 
.A(n_3048),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3059),
.B(n_2911),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3006),
.Y(n_3242)
);

OAI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_3058),
.A2(n_2722),
.B1(n_2777),
.B2(n_2789),
.Y(n_3243)
);

INVxp33_ASAP7_75t_SL g3244 ( 
.A(n_3039),
.Y(n_3244)
);

O2A1O1Ixp5_ASAP7_75t_L g3245 ( 
.A1(n_3109),
.A2(n_2955),
.B(n_2967),
.C(n_2958),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2989),
.Y(n_3246)
);

NOR2xp67_ASAP7_75t_L g3247 ( 
.A(n_3074),
.B(n_2902),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3164),
.A2(n_2857),
.B(n_2694),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_3023),
.B(n_2911),
.Y(n_3249)
);

OAI22xp5_ASAP7_75t_L g3250 ( 
.A1(n_3191),
.A2(n_2872),
.B1(n_2891),
.B2(n_2833),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_3166),
.A2(n_2694),
.B(n_2692),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3079),
.B(n_2911),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_3020),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3199),
.A2(n_2692),
.B(n_2811),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_3016),
.Y(n_3255)
);

BUFx8_ASAP7_75t_SL g3256 ( 
.A(n_2999),
.Y(n_3256)
);

BUFx6f_ASAP7_75t_L g3257 ( 
.A(n_3125),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_2984),
.B(n_3053),
.Y(n_3258)
);

OAI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_3118),
.A2(n_3127),
.B(n_3176),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_3024),
.Y(n_3260)
);

BUFx2_ASAP7_75t_L g3261 ( 
.A(n_2993),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3083),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3199),
.A2(n_2811),
.B(n_2465),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2990),
.Y(n_3264)
);

OAI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3055),
.A2(n_2702),
.B(n_2946),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3091),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_3095),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_3157),
.A2(n_2465),
.B(n_2409),
.Y(n_3268)
);

BUFx6f_ASAP7_75t_L g3269 ( 
.A(n_3125),
.Y(n_3269)
);

O2A1O1Ixp33_ASAP7_75t_L g3270 ( 
.A1(n_3123),
.A2(n_2912),
.B(n_2876),
.C(n_2861),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_3096),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_2982),
.B(n_2922),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2994),
.Y(n_3273)
);

OAI21xp33_ASAP7_75t_L g3274 ( 
.A1(n_3032),
.A2(n_2836),
.B(n_2818),
.Y(n_3274)
);

OR2x2_ASAP7_75t_L g3275 ( 
.A(n_3089),
.B(n_2702),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3202),
.B(n_2922),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3203),
.B(n_2922),
.Y(n_3277)
);

NOR2xp33_ASAP7_75t_SL g3278 ( 
.A(n_3056),
.B(n_3163),
.Y(n_3278)
);

OAI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_3175),
.A2(n_2946),
.B(n_2960),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3157),
.A2(n_2409),
.B(n_2932),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3086),
.B(n_3181),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_3151),
.B(n_2962),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2996),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_3187),
.A2(n_2941),
.B(n_2954),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3000),
.Y(n_3285)
);

OAI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_3077),
.A2(n_2964),
.B1(n_2924),
.B2(n_2873),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_SL g3287 ( 
.A(n_3192),
.B(n_2962),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2992),
.B(n_2960),
.Y(n_3288)
);

INVxp67_ASAP7_75t_L g3289 ( 
.A(n_3011),
.Y(n_3289)
);

O2A1O1Ixp33_ASAP7_75t_L g3290 ( 
.A1(n_3042),
.A2(n_2690),
.B(n_2949),
.C(n_2877),
.Y(n_3290)
);

INVx3_ASAP7_75t_L g3291 ( 
.A(n_3167),
.Y(n_3291)
);

INVx3_ASAP7_75t_L g3292 ( 
.A(n_3167),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3032),
.B(n_2682),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3134),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3131),
.B(n_2682),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_3110),
.A2(n_2896),
.B(n_2888),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3004),
.Y(n_3297)
);

CKINVDCx20_ASAP7_75t_R g3298 ( 
.A(n_3057),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_SL g3299 ( 
.A(n_3105),
.B(n_2962),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3062),
.B(n_2698),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_3110),
.A2(n_2896),
.B(n_2888),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3066),
.B(n_2698),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3168),
.A2(n_2849),
.B(n_2963),
.Y(n_3303)
);

BUFx6f_ASAP7_75t_L g3304 ( 
.A(n_3038),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3168),
.A2(n_2849),
.B(n_2963),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_SL g3306 ( 
.A(n_3010),
.B(n_2987),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3005),
.Y(n_3307)
);

AOI22x1_ASAP7_75t_L g3308 ( 
.A1(n_3033),
.A2(n_2703),
.B1(n_2713),
.B2(n_2962),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_3145),
.B(n_2703),
.Y(n_3309)
);

INVx3_ASAP7_75t_L g3310 ( 
.A(n_3139),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3078),
.B(n_2703),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3155),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3115),
.A2(n_2942),
.B(n_2864),
.Y(n_3313)
);

OAI21x1_ASAP7_75t_L g3314 ( 
.A1(n_3040),
.A2(n_2864),
.B(n_2919),
.Y(n_3314)
);

AOI21x1_ASAP7_75t_L g3315 ( 
.A1(n_3041),
.A2(n_2919),
.B(n_2975),
.Y(n_3315)
);

OAI21xp33_ASAP7_75t_L g3316 ( 
.A1(n_3022),
.A2(n_2878),
.B(n_2871),
.Y(n_3316)
);

HB1xp67_ASAP7_75t_L g3317 ( 
.A(n_3028),
.Y(n_3317)
);

OAI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_3129),
.A2(n_2884),
.B1(n_2890),
.B2(n_2930),
.Y(n_3318)
);

OAI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_3137),
.A2(n_2901),
.B1(n_2903),
.B2(n_2713),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_3115),
.A2(n_2903),
.B(n_2901),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3007),
.B(n_2713),
.Y(n_3321)
);

NOR3xp33_ASAP7_75t_L g3322 ( 
.A(n_2988),
.B(n_2962),
.C(n_6),
.Y(n_3322)
);

O2A1O1Ixp33_ASAP7_75t_L g3323 ( 
.A1(n_3012),
.A2(n_12),
.B(n_8),
.C(n_11),
.Y(n_3323)
);

NOR2x1p5_ASAP7_75t_SL g3324 ( 
.A(n_3197),
.B(n_3158),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3014),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3159),
.Y(n_3326)
);

OAI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3065),
.A2(n_1759),
.B(n_1752),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_3117),
.A2(n_3113),
.B(n_3033),
.Y(n_3328)
);

AOI22xp5_ASAP7_75t_L g3329 ( 
.A1(n_3169),
.A2(n_1242),
.B1(n_1759),
.B2(n_12),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3015),
.Y(n_3330)
);

O2A1O1Ixp33_ASAP7_75t_L g3331 ( 
.A1(n_3025),
.A2(n_13),
.B(n_8),
.C(n_11),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_3117),
.A2(n_1759),
.B(n_1242),
.Y(n_3332)
);

NOR2xp33_ASAP7_75t_L g3333 ( 
.A(n_3082),
.B(n_3107),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3113),
.A2(n_705),
.B(n_660),
.Y(n_3334)
);

BUFx4f_ASAP7_75t_L g3335 ( 
.A(n_3048),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3198),
.A2(n_685),
.B(n_684),
.Y(n_3336)
);

OAI21xp5_ASAP7_75t_L g3337 ( 
.A1(n_3031),
.A2(n_14),
.B(n_15),
.Y(n_3337)
);

NOR2x1_ASAP7_75t_L g3338 ( 
.A(n_3035),
.B(n_658),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_3072),
.B(n_3149),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_SL g3340 ( 
.A(n_3180),
.B(n_14),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3026),
.B(n_15),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3029),
.B(n_16),
.Y(n_3342)
);

HB1xp67_ASAP7_75t_L g3343 ( 
.A(n_3128),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3030),
.B(n_16),
.Y(n_3344)
);

AOI21x1_ASAP7_75t_L g3345 ( 
.A1(n_3041),
.A2(n_664),
.B(n_662),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3054),
.Y(n_3346)
);

A2O1A1Ixp33_ASAP7_75t_L g3347 ( 
.A1(n_3153),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_3347)
);

AND2x4_ASAP7_75t_L g3348 ( 
.A(n_3182),
.B(n_666),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3198),
.A2(n_698),
.B(n_697),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3063),
.B(n_17),
.Y(n_3350)
);

BUFx6f_ASAP7_75t_L g3351 ( 
.A(n_3061),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_3156),
.B(n_667),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_3084),
.B(n_18),
.Y(n_3353)
);

INVx4_ASAP7_75t_L g3354 ( 
.A(n_3183),
.Y(n_3354)
);

NOR3xp33_ASAP7_75t_L g3355 ( 
.A(n_3184),
.B(n_19),
.C(n_20),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_3126),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3064),
.B(n_20),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3067),
.Y(n_3358)
);

OAI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_3022),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3031),
.B(n_22),
.Y(n_3360)
);

O2A1O1Ixp33_ASAP7_75t_L g3361 ( 
.A1(n_3034),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_3361)
);

OAI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3031),
.A2(n_24),
.B(n_25),
.Y(n_3362)
);

AOI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3142),
.A2(n_690),
.B(n_689),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3044),
.Y(n_3364)
);

BUFx6f_ASAP7_75t_L g3365 ( 
.A(n_3165),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3087),
.B(n_26),
.Y(n_3366)
);

CKINVDCx5p33_ASAP7_75t_R g3367 ( 
.A(n_3076),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3092),
.B(n_26),
.Y(n_3368)
);

NOR2xp67_ASAP7_75t_L g3369 ( 
.A(n_3094),
.B(n_668),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3097),
.B(n_27),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3049),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3098),
.B(n_27),
.Y(n_3372)
);

BUFx6f_ASAP7_75t_SL g3373 ( 
.A(n_3121),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3099),
.B(n_28),
.Y(n_3374)
);

OAI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3196),
.A2(n_28),
.B(n_29),
.Y(n_3375)
);

BUFx2_ASAP7_75t_L g3376 ( 
.A(n_3138),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3101),
.B(n_29),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3185),
.B(n_669),
.Y(n_3378)
);

O2A1O1Ixp33_ASAP7_75t_L g3379 ( 
.A1(n_3051),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_3379)
);

INVx1_ASAP7_75t_SL g3380 ( 
.A(n_3103),
.Y(n_3380)
);

NAND3xp33_ASAP7_75t_SL g3381 ( 
.A(n_3073),
.B(n_30),
.C(n_31),
.Y(n_3381)
);

OAI22xp5_ASAP7_75t_L g3382 ( 
.A1(n_3019),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_3186),
.B(n_673),
.Y(n_3383)
);

AOI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_3142),
.A2(n_3037),
.B(n_3144),
.Y(n_3384)
);

AOI21xp5_ASAP7_75t_L g3385 ( 
.A1(n_3037),
.A2(n_677),
.B(n_676),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3108),
.B(n_33),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3112),
.B(n_34),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_3144),
.A2(n_686),
.B(n_683),
.Y(n_3388)
);

BUFx6f_ASAP7_75t_L g3389 ( 
.A(n_3046),
.Y(n_3389)
);

AND2x6_ASAP7_75t_L g3390 ( 
.A(n_3194),
.B(n_674),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_3132),
.A2(n_3148),
.B(n_3146),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3132),
.A2(n_694),
.B(n_693),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_L g3393 ( 
.A(n_3179),
.B(n_675),
.Y(n_3393)
);

OAI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3114),
.A2(n_35),
.B(n_36),
.Y(n_3394)
);

OAI21xp5_ASAP7_75t_L g3395 ( 
.A1(n_3116),
.A2(n_36),
.B(n_37),
.Y(n_3395)
);

BUFx6f_ASAP7_75t_L g3396 ( 
.A(n_3075),
.Y(n_3396)
);

AOI22xp5_ASAP7_75t_L g3397 ( 
.A1(n_3019),
.A2(n_3102),
.B1(n_3043),
.B2(n_3052),
.Y(n_3397)
);

NAND3xp33_ASAP7_75t_L g3398 ( 
.A(n_3090),
.B(n_37),
.C(n_38),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_L g3399 ( 
.A(n_3189),
.B(n_3190),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3080),
.Y(n_3400)
);

A2O1A1Ixp33_ASAP7_75t_L g3401 ( 
.A1(n_3081),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3122),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3124),
.B(n_40),
.Y(n_3403)
);

O2A1O1Ixp5_ASAP7_75t_L g3404 ( 
.A1(n_3130),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_3404)
);

INVxp67_ASAP7_75t_L g3405 ( 
.A(n_3050),
.Y(n_3405)
);

A2O1A1Ixp33_ASAP7_75t_L g3406 ( 
.A1(n_3135),
.A2(n_45),
.B(n_41),
.C(n_44),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3150),
.Y(n_3407)
);

AOI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_3146),
.A2(n_682),
.B(n_681),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_L g3409 ( 
.A(n_3193),
.B(n_691),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3148),
.A2(n_3093),
.B(n_3120),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3093),
.A2(n_699),
.B(n_696),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_3152),
.B(n_701),
.Y(n_3412)
);

BUFx6f_ASAP7_75t_L g3413 ( 
.A(n_3052),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_3102),
.B(n_703),
.Y(n_3414)
);

AOI22xp5_ASAP7_75t_L g3415 ( 
.A1(n_3043),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_3133),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3205),
.B(n_2983),
.Y(n_3417)
);

AOI21xp5_ASAP7_75t_L g3418 ( 
.A1(n_3279),
.A2(n_3172),
.B(n_3174),
.Y(n_3418)
);

A2O1A1Ixp33_ASAP7_75t_L g3419 ( 
.A1(n_3226),
.A2(n_2983),
.B(n_3085),
.C(n_3172),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3209),
.A2(n_3174),
.B(n_3071),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3281),
.B(n_3085),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3229),
.Y(n_3422)
);

INVx3_ASAP7_75t_L g3423 ( 
.A(n_3396),
.Y(n_3423)
);

AOI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_3221),
.A2(n_3071),
.B(n_3143),
.Y(n_3424)
);

O2A1O1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_3222),
.A2(n_3143),
.B(n_3178),
.C(n_3120),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3212),
.B(n_3275),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_3244),
.B(n_2995),
.Y(n_3427)
);

NOR2x1_ASAP7_75t_L g3428 ( 
.A(n_3217),
.B(n_3017),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3204),
.Y(n_3429)
);

A2O1A1Ixp33_ASAP7_75t_L g3430 ( 
.A1(n_3337),
.A2(n_3178),
.B(n_3001),
.C(n_2995),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3300),
.B(n_3302),
.Y(n_3431)
);

NOR3xp33_ASAP7_75t_SL g3432 ( 
.A(n_3381),
.B(n_3017),
.C(n_3001),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3396),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3265),
.A2(n_3119),
.B(n_3133),
.Y(n_3434)
);

O2A1O1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_3362),
.A2(n_3119),
.B(n_3161),
.C(n_48),
.Y(n_3435)
);

OAI21xp33_ASAP7_75t_L g3436 ( 
.A1(n_3375),
.A2(n_3161),
.B(n_46),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3330),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3231),
.A2(n_704),
.B(n_47),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3218),
.B(n_47),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_L g3440 ( 
.A(n_3258),
.B(n_48),
.Y(n_3440)
);

NOR2x1_ASAP7_75t_L g3441 ( 
.A(n_3228),
.B(n_49),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3211),
.A2(n_638),
.B(n_637),
.Y(n_3442)
);

BUFx6f_ASAP7_75t_L g3443 ( 
.A(n_3304),
.Y(n_3443)
);

CKINVDCx5p33_ASAP7_75t_R g3444 ( 
.A(n_3236),
.Y(n_3444)
);

O2A1O1Ixp5_ASAP7_75t_L g3445 ( 
.A1(n_3385),
.A2(n_53),
.B(n_50),
.C(n_51),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3248),
.A2(n_639),
.B(n_637),
.Y(n_3446)
);

A2O1A1Ixp33_ASAP7_75t_L g3447 ( 
.A1(n_3208),
.A2(n_53),
.B(n_50),
.C(n_51),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_3206),
.A2(n_645),
.B(n_644),
.Y(n_3448)
);

OAI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3259),
.A2(n_54),
.B(n_55),
.Y(n_3449)
);

NOR3xp33_ASAP7_75t_SL g3450 ( 
.A(n_3414),
.B(n_645),
.C(n_644),
.Y(n_3450)
);

OAI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_3335),
.A2(n_58),
.B1(n_54),
.B2(n_57),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3216),
.A2(n_650),
.B(n_59),
.Y(n_3452)
);

BUFx12f_ASAP7_75t_L g3453 ( 
.A(n_3367),
.Y(n_3453)
);

INVxp67_ASAP7_75t_L g3454 ( 
.A(n_3261),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_3220),
.B(n_60),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3346),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3335),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_3457)
);

BUFx12f_ASAP7_75t_L g3458 ( 
.A(n_3356),
.Y(n_3458)
);

O2A1O1Ixp5_ASAP7_75t_SL g3459 ( 
.A1(n_3382),
.A2(n_64),
.B(n_61),
.C(n_63),
.Y(n_3459)
);

HB1xp67_ASAP7_75t_L g3460 ( 
.A(n_3237),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3207),
.B(n_64),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3288),
.B(n_65),
.Y(n_3462)
);

INVx4_ASAP7_75t_L g3463 ( 
.A(n_3210),
.Y(n_3463)
);

A2O1A1Ixp33_ASAP7_75t_L g3464 ( 
.A1(n_3394),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3241),
.B(n_66),
.Y(n_3465)
);

NAND2x1p5_ASAP7_75t_L g3466 ( 
.A(n_3210),
.B(n_67),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_SL g3467 ( 
.A(n_3234),
.B(n_68),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3246),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3233),
.B(n_3380),
.Y(n_3469)
);

A2O1A1Ixp33_ASAP7_75t_SL g3470 ( 
.A1(n_3395),
.A2(n_636),
.B(n_639),
.C(n_635),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3333),
.B(n_68),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3215),
.B(n_69),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_3256),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3238),
.B(n_69),
.Y(n_3474)
);

AOI22xp5_ASAP7_75t_L g3475 ( 
.A1(n_3322),
.A2(n_73),
.B1(n_70),
.B2(n_71),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3239),
.B(n_70),
.Y(n_3476)
);

AOI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_3254),
.A2(n_650),
.B(n_649),
.Y(n_3477)
);

CKINVDCx20_ASAP7_75t_R g3478 ( 
.A(n_3298),
.Y(n_3478)
);

AOI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_3251),
.A2(n_3284),
.B(n_3230),
.Y(n_3479)
);

NOR2xp67_ASAP7_75t_SL g3480 ( 
.A(n_3398),
.B(n_73),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3243),
.B(n_74),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_SL g3482 ( 
.A(n_3396),
.B(n_3247),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3303),
.A2(n_77),
.B(n_78),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3264),
.Y(n_3484)
);

INVx2_ASAP7_75t_SL g3485 ( 
.A(n_3253),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3358),
.Y(n_3486)
);

BUFx6f_ASAP7_75t_L g3487 ( 
.A(n_3304),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3272),
.B(n_77),
.Y(n_3488)
);

BUFx6f_ASAP7_75t_L g3489 ( 
.A(n_3304),
.Y(n_3489)
);

O2A1O1Ixp33_ASAP7_75t_L g3490 ( 
.A1(n_3401),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_3490)
);

O2A1O1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_3347),
.A2(n_82),
.B(n_79),
.C(n_81),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3213),
.Y(n_3492)
);

BUFx3_ASAP7_75t_L g3493 ( 
.A(n_3311),
.Y(n_3493)
);

INVx3_ASAP7_75t_L g3494 ( 
.A(n_3291),
.Y(n_3494)
);

AOI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_3305),
.A2(n_632),
.B(n_631),
.Y(n_3495)
);

INVxp67_ASAP7_75t_SL g3496 ( 
.A(n_3247),
.Y(n_3496)
);

A2O1A1Ixp33_ASAP7_75t_SL g3497 ( 
.A1(n_3336),
.A2(n_632),
.B(n_633),
.C(n_630),
.Y(n_3497)
);

CKINVDCx5p33_ASAP7_75t_R g3498 ( 
.A(n_3373),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3225),
.Y(n_3499)
);

AOI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3299),
.A2(n_85),
.B1(n_82),
.B2(n_83),
.Y(n_3500)
);

AOI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_3340),
.A2(n_86),
.B1(n_83),
.B2(n_85),
.Y(n_3501)
);

CKINVDCx16_ASAP7_75t_R g3502 ( 
.A(n_3306),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_SL g3503 ( 
.A(n_3376),
.B(n_87),
.Y(n_3503)
);

INVx3_ASAP7_75t_L g3504 ( 
.A(n_3291),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3295),
.B(n_3252),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_3286),
.B(n_87),
.Y(n_3506)
);

OAI22xp5_ASAP7_75t_L g3507 ( 
.A1(n_3329),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_3507)
);

NOR2xp33_ASAP7_75t_SL g3508 ( 
.A(n_3278),
.B(n_3405),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3296),
.A2(n_649),
.B(n_89),
.Y(n_3509)
);

AND2x4_ASAP7_75t_L g3510 ( 
.A(n_3292),
.B(n_91),
.Y(n_3510)
);

OAI21x1_ASAP7_75t_L g3511 ( 
.A1(n_3314),
.A2(n_92),
.B(n_93),
.Y(n_3511)
);

HB1xp67_ASAP7_75t_L g3512 ( 
.A(n_3416),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3242),
.B(n_3255),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3260),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3301),
.A2(n_92),
.B(n_93),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3262),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3289),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3355),
.A2(n_97),
.B1(n_94),
.B2(n_96),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3402),
.B(n_648),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3360),
.B(n_98),
.Y(n_3520)
);

INVx4_ASAP7_75t_L g3521 ( 
.A(n_3257),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3273),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3266),
.Y(n_3523)
);

NOR2x1_ASAP7_75t_L g3524 ( 
.A(n_3249),
.B(n_99),
.Y(n_3524)
);

NAND2x1p5_ASAP7_75t_L g3525 ( 
.A(n_3354),
.B(n_99),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3267),
.Y(n_3526)
);

BUFx3_ASAP7_75t_L g3527 ( 
.A(n_3257),
.Y(n_3527)
);

O2A1O1Ixp33_ASAP7_75t_L g3528 ( 
.A1(n_3406),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_3528)
);

BUFx6f_ASAP7_75t_L g3529 ( 
.A(n_3257),
.Y(n_3529)
);

OAI21xp33_ASAP7_75t_SL g3530 ( 
.A1(n_3415),
.A2(n_104),
.B(n_105),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3283),
.Y(n_3531)
);

AO32x2_ASAP7_75t_L g3532 ( 
.A1(n_3359),
.A2(n_106),
.A3(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_3532)
);

OAI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3245),
.A2(n_107),
.B(n_108),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3271),
.Y(n_3534)
);

A2O1A1Ixp33_ASAP7_75t_L g3535 ( 
.A1(n_3349),
.A2(n_3411),
.B(n_3323),
.C(n_3361),
.Y(n_3535)
);

AND2x2_ASAP7_75t_L g3536 ( 
.A(n_3293),
.B(n_109),
.Y(n_3536)
);

BUFx10_ASAP7_75t_L g3537 ( 
.A(n_3373),
.Y(n_3537)
);

NOR2xp33_ASAP7_75t_R g3538 ( 
.A(n_3240),
.B(n_109),
.Y(n_3538)
);

A2O1A1Ixp33_ASAP7_75t_L g3539 ( 
.A1(n_3331),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3285),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3407),
.B(n_110),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3294),
.B(n_648),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3297),
.Y(n_3543)
);

INVxp67_ASAP7_75t_L g3544 ( 
.A(n_3317),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3312),
.B(n_113),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3307),
.Y(n_3546)
);

BUFx6f_ASAP7_75t_L g3547 ( 
.A(n_3269),
.Y(n_3547)
);

BUFx6f_ASAP7_75t_L g3548 ( 
.A(n_3269),
.Y(n_3548)
);

OAI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3318),
.A2(n_114),
.B(n_115),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3326),
.B(n_647),
.Y(n_3550)
);

AOI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3313),
.A2(n_114),
.B(n_115),
.Y(n_3551)
);

AOI22xp33_ASAP7_75t_L g3552 ( 
.A1(n_3274),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_3552)
);

NOR2xp33_ASAP7_75t_L g3553 ( 
.A(n_3339),
.B(n_3223),
.Y(n_3553)
);

OAI21x1_ASAP7_75t_L g3554 ( 
.A1(n_3235),
.A2(n_118),
.B(n_119),
.Y(n_3554)
);

INVx4_ASAP7_75t_L g3555 ( 
.A(n_3269),
.Y(n_3555)
);

INVx3_ASAP7_75t_L g3556 ( 
.A(n_3292),
.Y(n_3556)
);

NOR2xp33_ASAP7_75t_L g3557 ( 
.A(n_3232),
.B(n_119),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3325),
.Y(n_3558)
);

HB1xp67_ASAP7_75t_L g3559 ( 
.A(n_3364),
.Y(n_3559)
);

AND2x4_ASAP7_75t_L g3560 ( 
.A(n_3371),
.B(n_120),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_SL g3561 ( 
.A(n_3290),
.B(n_3338),
.Y(n_3561)
);

A2O1A1Ixp33_ASAP7_75t_L g3562 ( 
.A1(n_3379),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3309),
.B(n_122),
.Y(n_3563)
);

O2A1O1Ixp33_ASAP7_75t_SL g3564 ( 
.A1(n_3353),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_3224),
.A2(n_124),
.B(n_126),
.Y(n_3565)
);

O2A1O1Ixp33_ASAP7_75t_L g3566 ( 
.A1(n_3404),
.A2(n_130),
.B(n_127),
.C(n_129),
.Y(n_3566)
);

NOR3xp33_ASAP7_75t_L g3567 ( 
.A(n_3316),
.B(n_127),
.C(n_129),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3276),
.B(n_647),
.Y(n_3568)
);

O2A1O1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_3319),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3227),
.A2(n_131),
.B(n_132),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3400),
.Y(n_3571)
);

BUFx2_ASAP7_75t_L g3572 ( 
.A(n_3343),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3399),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3413),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_3277),
.B(n_134),
.Y(n_3575)
);

AOI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_3219),
.A2(n_135),
.B(n_136),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3413),
.Y(n_3577)
);

O2A1O1Ixp33_ASAP7_75t_SL g3578 ( 
.A1(n_3341),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3342),
.B(n_137),
.Y(n_3579)
);

A2O1A1Ixp33_ASAP7_75t_L g3580 ( 
.A1(n_3397),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_3580)
);

AOI22xp33_ASAP7_75t_L g3581 ( 
.A1(n_3390),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_3581)
);

INVx3_ASAP7_75t_L g3582 ( 
.A(n_3354),
.Y(n_3582)
);

A2O1A1Ixp33_ASAP7_75t_SL g3583 ( 
.A1(n_3363),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_3583)
);

BUFx3_ASAP7_75t_L g3584 ( 
.A(n_3351),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3390),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3413),
.Y(n_3586)
);

NOR2xp33_ASAP7_75t_L g3587 ( 
.A(n_3352),
.B(n_144),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3344),
.B(n_145),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_SL g3589 ( 
.A(n_3250),
.B(n_146),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3327),
.A2(n_146),
.B(n_147),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3321),
.Y(n_3591)
);

NOR2xp67_ASAP7_75t_SL g3592 ( 
.A(n_3408),
.B(n_147),
.Y(n_3592)
);

HB1xp67_ASAP7_75t_L g3593 ( 
.A(n_3287),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3350),
.B(n_646),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_3263),
.A2(n_148),
.B(n_150),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_3268),
.A2(n_148),
.B(n_151),
.Y(n_3596)
);

OAI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3282),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_3597)
);

NOR2xp33_ASAP7_75t_L g3598 ( 
.A(n_3240),
.B(n_152),
.Y(n_3598)
);

NOR2xp33_ASAP7_75t_L g3599 ( 
.A(n_3366),
.B(n_154),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3357),
.B(n_643),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3280),
.A2(n_154),
.B(n_155),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3368),
.B(n_3370),
.Y(n_3602)
);

O2A1O1Ixp33_ASAP7_75t_L g3603 ( 
.A1(n_3334),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_3603)
);

O2A1O1Ixp33_ASAP7_75t_L g3604 ( 
.A1(n_3372),
.A2(n_159),
.B(n_156),
.C(n_158),
.Y(n_3604)
);

A2O1A1Ixp33_ASAP7_75t_L g3605 ( 
.A1(n_3388),
.A2(n_3392),
.B(n_3384),
.C(n_3391),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3348),
.Y(n_3606)
);

NAND3xp33_ASAP7_75t_L g3607 ( 
.A(n_3412),
.B(n_160),
.C(n_161),
.Y(n_3607)
);

NAND3xp33_ASAP7_75t_SL g3608 ( 
.A(n_3270),
.B(n_161),
.C(n_162),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_3369),
.B(n_163),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_3320),
.A2(n_163),
.B(n_164),
.Y(n_3610)
);

BUFx8_ASAP7_75t_SL g3611 ( 
.A(n_3351),
.Y(n_3611)
);

O2A1O1Ixp33_ASAP7_75t_L g3612 ( 
.A1(n_3374),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_3612)
);

NOR2xp33_ASAP7_75t_L g3613 ( 
.A(n_3377),
.B(n_168),
.Y(n_3613)
);

O2A1O1Ixp33_ASAP7_75t_L g3614 ( 
.A1(n_3386),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_3614)
);

BUFx6f_ASAP7_75t_SL g3615 ( 
.A(n_3390),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_3332),
.A2(n_169),
.B(n_171),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3348),
.Y(n_3617)
);

OAI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3308),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_3618)
);

BUFx6f_ASAP7_75t_L g3619 ( 
.A(n_3351),
.Y(n_3619)
);

NOR2xp67_ASAP7_75t_SL g3620 ( 
.A(n_3310),
.B(n_172),
.Y(n_3620)
);

AO21x2_ASAP7_75t_L g3621 ( 
.A1(n_3345),
.A2(n_174),
.B(n_175),
.Y(n_3621)
);

CKINVDCx10_ASAP7_75t_R g3622 ( 
.A(n_3365),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3214),
.A2(n_176),
.B(n_178),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3387),
.Y(n_3624)
);

AOI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_3328),
.A2(n_176),
.B(n_179),
.Y(n_3625)
);

CKINVDCx5p33_ASAP7_75t_R g3626 ( 
.A(n_3365),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3410),
.A2(n_179),
.B(n_181),
.Y(n_3627)
);

OR2x2_ASAP7_75t_L g3628 ( 
.A(n_3403),
.B(n_181),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3559),
.Y(n_3629)
);

BUFx8_ASAP7_75t_SL g3630 ( 
.A(n_3478),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3437),
.Y(n_3631)
);

AND2x4_ASAP7_75t_L g3632 ( 
.A(n_3574),
.B(n_3324),
.Y(n_3632)
);

INVx4_ASAP7_75t_L g3633 ( 
.A(n_3463),
.Y(n_3633)
);

INVxp67_ASAP7_75t_SL g3634 ( 
.A(n_3460),
.Y(n_3634)
);

AND2x4_ASAP7_75t_L g3635 ( 
.A(n_3577),
.B(n_3315),
.Y(n_3635)
);

AND2x4_ASAP7_75t_L g3636 ( 
.A(n_3586),
.B(n_3310),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3426),
.B(n_3378),
.Y(n_3637)
);

BUFx2_ASAP7_75t_L g3638 ( 
.A(n_3512),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3456),
.Y(n_3639)
);

BUFx2_ASAP7_75t_L g3640 ( 
.A(n_3593),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3486),
.Y(n_3641)
);

HB1xp67_ASAP7_75t_L g3642 ( 
.A(n_3572),
.Y(n_3642)
);

INVx4_ASAP7_75t_L g3643 ( 
.A(n_3626),
.Y(n_3643)
);

OR2x6_ASAP7_75t_L g3644 ( 
.A(n_3424),
.B(n_3389),
.Y(n_3644)
);

BUFx6f_ASAP7_75t_L g3645 ( 
.A(n_3529),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_SL g3646 ( 
.A(n_3502),
.B(n_3389),
.Y(n_3646)
);

CKINVDCx8_ASAP7_75t_R g3647 ( 
.A(n_3622),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3422),
.Y(n_3648)
);

INVx3_ASAP7_75t_L g3649 ( 
.A(n_3611),
.Y(n_3649)
);

AOI22x1_ASAP7_75t_L g3650 ( 
.A1(n_3551),
.A2(n_3389),
.B1(n_3365),
.B2(n_3390),
.Y(n_3650)
);

OR2x2_ASAP7_75t_L g3651 ( 
.A(n_3417),
.B(n_3393),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3468),
.Y(n_3652)
);

INVx2_ASAP7_75t_SL g3653 ( 
.A(n_3537),
.Y(n_3653)
);

BUFx2_ASAP7_75t_L g3654 ( 
.A(n_3428),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3484),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_3522),
.B(n_3369),
.Y(n_3656)
);

INVx5_ASAP7_75t_L g3657 ( 
.A(n_3537),
.Y(n_3657)
);

BUFx2_ASAP7_75t_L g3658 ( 
.A(n_3496),
.Y(n_3658)
);

INVx5_ASAP7_75t_L g3659 ( 
.A(n_3582),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3531),
.Y(n_3660)
);

NOR2xp67_ASAP7_75t_L g3661 ( 
.A(n_3624),
.B(n_3409),
.Y(n_3661)
);

BUFx2_ASAP7_75t_L g3662 ( 
.A(n_3494),
.Y(n_3662)
);

BUFx12f_ASAP7_75t_L g3663 ( 
.A(n_3444),
.Y(n_3663)
);

O2A1O1Ixp33_ASAP7_75t_L g3664 ( 
.A1(n_3539),
.A2(n_3383),
.B(n_184),
.C(n_182),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3431),
.B(n_182),
.Y(n_3665)
);

BUFx2_ASAP7_75t_L g3666 ( 
.A(n_3494),
.Y(n_3666)
);

INVx3_ASAP7_75t_L g3667 ( 
.A(n_3619),
.Y(n_3667)
);

OR2x2_ASAP7_75t_L g3668 ( 
.A(n_3540),
.B(n_183),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3505),
.B(n_183),
.Y(n_3669)
);

BUFx6f_ASAP7_75t_L g3670 ( 
.A(n_3529),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3591),
.B(n_184),
.Y(n_3671)
);

O2A1O1Ixp5_ASAP7_75t_L g3672 ( 
.A1(n_3449),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_3672)
);

INVx4_ASAP7_75t_L g3673 ( 
.A(n_3619),
.Y(n_3673)
);

INVx3_ASAP7_75t_L g3674 ( 
.A(n_3619),
.Y(n_3674)
);

INVx5_ASAP7_75t_L g3675 ( 
.A(n_3582),
.Y(n_3675)
);

AND2x4_ASAP7_75t_L g3676 ( 
.A(n_3543),
.B(n_186),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3546),
.Y(n_3677)
);

OAI21x1_ASAP7_75t_L g3678 ( 
.A1(n_3479),
.A2(n_187),
.B(n_189),
.Y(n_3678)
);

XNOR2xp5_ASAP7_75t_SL g3679 ( 
.A(n_3473),
.B(n_3498),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3558),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3571),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3429),
.Y(n_3682)
);

NAND2x1p5_ASAP7_75t_L g3683 ( 
.A(n_3423),
.B(n_189),
.Y(n_3683)
);

BUFx6f_ASAP7_75t_L g3684 ( 
.A(n_3529),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_3453),
.Y(n_3685)
);

BUFx4_ASAP7_75t_SL g3686 ( 
.A(n_3493),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3573),
.B(n_190),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_3441),
.B(n_191),
.Y(n_3688)
);

BUFx6f_ASAP7_75t_L g3689 ( 
.A(n_3547),
.Y(n_3689)
);

BUFx6f_ASAP7_75t_L g3690 ( 
.A(n_3547),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3421),
.B(n_191),
.Y(n_3691)
);

INVx3_ASAP7_75t_L g3692 ( 
.A(n_3521),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3492),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3499),
.Y(n_3694)
);

AOI22xp33_ASAP7_75t_SL g3695 ( 
.A1(n_3615),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_3695)
);

O2A1O1Ixp33_ASAP7_75t_L g3696 ( 
.A1(n_3562),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_3696)
);

BUFx2_ASAP7_75t_L g3697 ( 
.A(n_3504),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3488),
.B(n_640),
.Y(n_3698)
);

INVx5_ASAP7_75t_L g3699 ( 
.A(n_3463),
.Y(n_3699)
);

OR2x6_ASAP7_75t_SL g3700 ( 
.A(n_3607),
.B(n_196),
.Y(n_3700)
);

OAI22xp5_ASAP7_75t_SL g3701 ( 
.A1(n_3440),
.A2(n_201),
.B1(n_196),
.B2(n_200),
.Y(n_3701)
);

AOI22xp33_ASAP7_75t_SL g3702 ( 
.A1(n_3615),
.A2(n_204),
.B1(n_200),
.B2(n_202),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3514),
.Y(n_3703)
);

AOI21xp5_ASAP7_75t_L g3704 ( 
.A1(n_3418),
.A2(n_202),
.B(n_206),
.Y(n_3704)
);

BUFx12f_ASAP7_75t_L g3705 ( 
.A(n_3458),
.Y(n_3705)
);

BUFx3_ASAP7_75t_L g3706 ( 
.A(n_3584),
.Y(n_3706)
);

INVx3_ASAP7_75t_L g3707 ( 
.A(n_3521),
.Y(n_3707)
);

AOI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3467),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_3708)
);

INVx3_ASAP7_75t_L g3709 ( 
.A(n_3555),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3516),
.Y(n_3710)
);

AO32x2_ASAP7_75t_L g3711 ( 
.A1(n_3618),
.A2(n_211),
.A3(n_207),
.B1(n_209),
.B2(n_212),
.Y(n_3711)
);

INVx5_ASAP7_75t_L g3712 ( 
.A(n_3443),
.Y(n_3712)
);

NOR2xp33_ASAP7_75t_L g3713 ( 
.A(n_3553),
.B(n_211),
.Y(n_3713)
);

BUFx12f_ASAP7_75t_L g3714 ( 
.A(n_3485),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3455),
.B(n_640),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3602),
.B(n_212),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3549),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_3717)
);

INVx3_ASAP7_75t_L g3718 ( 
.A(n_3555),
.Y(n_3718)
);

AO22x1_ASAP7_75t_L g3719 ( 
.A1(n_3567),
.A2(n_218),
.B1(n_215),
.B2(n_216),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3523),
.Y(n_3720)
);

INVx8_ASAP7_75t_L g3721 ( 
.A(n_3547),
.Y(n_3721)
);

AOI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_3481),
.A2(n_3506),
.B1(n_3589),
.B2(n_3480),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3526),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3534),
.Y(n_3724)
);

OR2x2_ASAP7_75t_L g3725 ( 
.A(n_3469),
.B(n_218),
.Y(n_3725)
);

BUFx3_ASAP7_75t_L g3726 ( 
.A(n_3527),
.Y(n_3726)
);

INVx3_ASAP7_75t_L g3727 ( 
.A(n_3548),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3454),
.B(n_219),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3504),
.Y(n_3729)
);

INVx3_ASAP7_75t_L g3730 ( 
.A(n_3548),
.Y(n_3730)
);

OAI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3581),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_3731)
);

BUFx4f_ASAP7_75t_SL g3732 ( 
.A(n_3443),
.Y(n_3732)
);

OAI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3585),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_3733)
);

BUFx6f_ASAP7_75t_L g3734 ( 
.A(n_3548),
.Y(n_3734)
);

HB1xp67_ASAP7_75t_L g3735 ( 
.A(n_3556),
.Y(n_3735)
);

NOR2xp33_ASAP7_75t_L g3736 ( 
.A(n_3508),
.B(n_222),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3513),
.Y(n_3737)
);

AND2x6_ASAP7_75t_L g3738 ( 
.A(n_3524),
.B(n_223),
.Y(n_3738)
);

AOI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_3561),
.A2(n_224),
.B(n_225),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3556),
.Y(n_3740)
);

AND2x4_ASAP7_75t_L g3741 ( 
.A(n_3423),
.B(n_224),
.Y(n_3741)
);

AND2x4_ASAP7_75t_L g3742 ( 
.A(n_3433),
.B(n_225),
.Y(n_3742)
);

INVx3_ASAP7_75t_L g3743 ( 
.A(n_3443),
.Y(n_3743)
);

AOI21x1_ASAP7_75t_L g3744 ( 
.A1(n_3592),
.A2(n_226),
.B(n_227),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_3420),
.A2(n_226),
.B(n_228),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3533),
.A2(n_228),
.B(n_229),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3544),
.B(n_229),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_3538),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3535),
.A2(n_230),
.B(n_231),
.Y(n_3749)
);

BUFx2_ASAP7_75t_L g3750 ( 
.A(n_3433),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_SL g3751 ( 
.A(n_3450),
.B(n_230),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_SL g3752 ( 
.A1(n_3530),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_3752)
);

AO21x2_ASAP7_75t_L g3753 ( 
.A1(n_3483),
.A2(n_232),
.B(n_234),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3425),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3519),
.Y(n_3755)
);

INVx5_ASAP7_75t_L g3756 ( 
.A(n_3487),
.Y(n_3756)
);

OAI22xp33_ASAP7_75t_L g3757 ( 
.A1(n_3475),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3482),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3541),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3461),
.B(n_235),
.Y(n_3760)
);

AOI221xp5_ASAP7_75t_L g3761 ( 
.A1(n_3604),
.A2(n_239),
.B1(n_236),
.B2(n_238),
.C(n_241),
.Y(n_3761)
);

INVxp67_ASAP7_75t_L g3762 ( 
.A(n_3487),
.Y(n_3762)
);

AOI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3436),
.A2(n_242),
.B1(n_239),
.B2(n_241),
.Y(n_3763)
);

AOI22xp33_ASAP7_75t_L g3764 ( 
.A1(n_3587),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_3764)
);

OR2x6_ASAP7_75t_L g3765 ( 
.A(n_3434),
.B(n_244),
.Y(n_3765)
);

AOI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3520),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_3766)
);

INVx3_ASAP7_75t_L g3767 ( 
.A(n_3487),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3511),
.Y(n_3768)
);

BUFx2_ASAP7_75t_L g3769 ( 
.A(n_3605),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3542),
.Y(n_3770)
);

CKINVDCx5p33_ASAP7_75t_R g3771 ( 
.A(n_3489),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3545),
.Y(n_3772)
);

BUFx6f_ASAP7_75t_L g3773 ( 
.A(n_3489),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3550),
.Y(n_3774)
);

INVxp67_ASAP7_75t_L g3775 ( 
.A(n_3489),
.Y(n_3775)
);

INVx1_ASAP7_75t_SL g3776 ( 
.A(n_3563),
.Y(n_3776)
);

INVx4_ASAP7_75t_L g3777 ( 
.A(n_3560),
.Y(n_3777)
);

BUFx2_ASAP7_75t_L g3778 ( 
.A(n_3419),
.Y(n_3778)
);

INVx3_ASAP7_75t_L g3779 ( 
.A(n_3510),
.Y(n_3779)
);

HB1xp67_ASAP7_75t_L g3780 ( 
.A(n_3554),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3474),
.Y(n_3781)
);

BUFx3_ASAP7_75t_L g3782 ( 
.A(n_3510),
.Y(n_3782)
);

AND2x4_ASAP7_75t_L g3783 ( 
.A(n_3427),
.B(n_246),
.Y(n_3783)
);

OAI221xp5_ASAP7_75t_L g3784 ( 
.A1(n_3518),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.C(n_250),
.Y(n_3784)
);

AOI22xp33_ASAP7_75t_L g3785 ( 
.A1(n_3608),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_3785)
);

AND2x4_ASAP7_75t_L g3786 ( 
.A(n_3606),
.B(n_251),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3621),
.Y(n_3787)
);

INVx4_ASAP7_75t_L g3788 ( 
.A(n_3560),
.Y(n_3788)
);

AND2x4_ASAP7_75t_L g3789 ( 
.A(n_3617),
.B(n_252),
.Y(n_3789)
);

AND2x4_ASAP7_75t_L g3790 ( 
.A(n_3430),
.B(n_252),
.Y(n_3790)
);

BUFx6f_ASAP7_75t_L g3791 ( 
.A(n_3568),
.Y(n_3791)
);

INVx4_ASAP7_75t_L g3792 ( 
.A(n_3466),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3621),
.Y(n_3793)
);

BUFx3_ASAP7_75t_L g3794 ( 
.A(n_3462),
.Y(n_3794)
);

INVx5_ASAP7_75t_L g3795 ( 
.A(n_3536),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3588),
.B(n_253),
.Y(n_3796)
);

BUFx2_ASAP7_75t_SL g3797 ( 
.A(n_3609),
.Y(n_3797)
);

BUFx10_ASAP7_75t_L g3798 ( 
.A(n_3598),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3465),
.Y(n_3799)
);

BUFx6f_ASAP7_75t_L g3800 ( 
.A(n_3476),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3557),
.B(n_253),
.Y(n_3801)
);

OR2x6_ASAP7_75t_L g3802 ( 
.A(n_3610),
.B(n_254),
.Y(n_3802)
);

BUFx6f_ASAP7_75t_SL g3803 ( 
.A(n_3503),
.Y(n_3803)
);

AND2x4_ASAP7_75t_L g3804 ( 
.A(n_3432),
.B(n_255),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3472),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3532),
.Y(n_3806)
);

AOI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3452),
.A2(n_256),
.B(n_257),
.Y(n_3807)
);

NOR2x1_ASAP7_75t_L g3808 ( 
.A(n_3477),
.B(n_256),
.Y(n_3808)
);

OAI21x1_ASAP7_75t_SL g3809 ( 
.A1(n_3435),
.A2(n_257),
.B(n_258),
.Y(n_3809)
);

INVx4_ASAP7_75t_L g3810 ( 
.A(n_3525),
.Y(n_3810)
);

INVx2_ASAP7_75t_SL g3811 ( 
.A(n_3628),
.Y(n_3811)
);

OR2x2_ASAP7_75t_L g3812 ( 
.A(n_3579),
.B(n_3594),
.Y(n_3812)
);

NAND2x2_ASAP7_75t_L g3813 ( 
.A(n_3439),
.B(n_258),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3575),
.B(n_259),
.Y(n_3814)
);

OAI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3500),
.A2(n_262),
.B1(n_259),
.B2(n_260),
.Y(n_3815)
);

OAI22xp5_ASAP7_75t_L g3816 ( 
.A1(n_3552),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_3816)
);

INVx2_ASAP7_75t_SL g3817 ( 
.A(n_3600),
.Y(n_3817)
);

INVx3_ASAP7_75t_L g3818 ( 
.A(n_3620),
.Y(n_3818)
);

INVx1_ASAP7_75t_SL g3819 ( 
.A(n_3471),
.Y(n_3819)
);

AOI21x1_ASAP7_75t_L g3820 ( 
.A1(n_3616),
.A2(n_263),
.B(n_265),
.Y(n_3820)
);

CKINVDCx20_ASAP7_75t_R g3821 ( 
.A(n_3599),
.Y(n_3821)
);

CKINVDCx5p33_ASAP7_75t_R g3822 ( 
.A(n_3613),
.Y(n_3822)
);

AOI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3507),
.A2(n_3457),
.B1(n_3451),
.B2(n_3464),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3495),
.B(n_266),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3532),
.Y(n_3825)
);

INVx5_ASAP7_75t_L g3826 ( 
.A(n_3497),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_3501),
.B(n_267),
.Y(n_3827)
);

INVx5_ASAP7_75t_L g3828 ( 
.A(n_3583),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3532),
.Y(n_3829)
);

BUFx6f_ASAP7_75t_L g3830 ( 
.A(n_3564),
.Y(n_3830)
);

BUFx3_ASAP7_75t_L g3831 ( 
.A(n_3597),
.Y(n_3831)
);

BUFx6f_ASAP7_75t_L g3832 ( 
.A(n_3576),
.Y(n_3832)
);

NAND2x1p5_ASAP7_75t_L g3833 ( 
.A(n_3438),
.B(n_267),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3509),
.Y(n_3834)
);

INVx3_ASAP7_75t_SL g3835 ( 
.A(n_3578),
.Y(n_3835)
);

CKINVDCx20_ASAP7_75t_R g3836 ( 
.A(n_3517),
.Y(n_3836)
);

OAI22xp5_ASAP7_75t_SL g3837 ( 
.A1(n_3580),
.A2(n_3491),
.B1(n_3569),
.B2(n_3612),
.Y(n_3837)
);

OR2x6_ASAP7_75t_L g3838 ( 
.A(n_3515),
.B(n_268),
.Y(n_3838)
);

OAI22xp5_ASAP7_75t_L g3839 ( 
.A1(n_3447),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_3839)
);

NOR2xp33_ASAP7_75t_L g3840 ( 
.A(n_3614),
.B(n_269),
.Y(n_3840)
);

BUFx2_ASAP7_75t_L g3841 ( 
.A(n_3595),
.Y(n_3841)
);

AOI21xp33_ASAP7_75t_L g3842 ( 
.A1(n_3470),
.A2(n_270),
.B(n_271),
.Y(n_3842)
);

NOR2x1p5_ASAP7_75t_L g3843 ( 
.A(n_3490),
.B(n_271),
.Y(n_3843)
);

AOI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3627),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3625),
.B(n_272),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3601),
.Y(n_3846)
);

AOI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_3590),
.A2(n_3446),
.B1(n_3442),
.B2(n_3448),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3565),
.B(n_273),
.Y(n_3848)
);

OAI33xp33_ASAP7_75t_L g3849 ( 
.A1(n_3528),
.A2(n_276),
.A3(n_278),
.B1(n_274),
.B2(n_275),
.B3(n_277),
.Y(n_3849)
);

NOR2xp33_ASAP7_75t_L g3850 ( 
.A(n_3570),
.B(n_275),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3603),
.A2(n_277),
.B(n_279),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3566),
.Y(n_3852)
);

HB1xp67_ASAP7_75t_L g3853 ( 
.A(n_3623),
.Y(n_3853)
);

BUFx6f_ASAP7_75t_L g3854 ( 
.A(n_3596),
.Y(n_3854)
);

BUFx3_ASAP7_75t_L g3855 ( 
.A(n_3445),
.Y(n_3855)
);

INVx1_ASAP7_75t_SL g3856 ( 
.A(n_3459),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3505),
.B(n_634),
.Y(n_3857)
);

INVx3_ASAP7_75t_L g3858 ( 
.A(n_3611),
.Y(n_3858)
);

BUFx3_ASAP7_75t_L g3859 ( 
.A(n_3714),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3660),
.Y(n_3860)
);

OR2x2_ASAP7_75t_L g3861 ( 
.A(n_3629),
.B(n_279),
.Y(n_3861)
);

INVx4_ASAP7_75t_L g3862 ( 
.A(n_3699),
.Y(n_3862)
);

OAI22xp5_ASAP7_75t_L g3863 ( 
.A1(n_3823),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3863)
);

BUFx2_ASAP7_75t_L g3864 ( 
.A(n_3640),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3648),
.Y(n_3865)
);

AOI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3769),
.A2(n_280),
.B(n_282),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3680),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_3630),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3681),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3634),
.B(n_283),
.Y(n_3870)
);

OR2x6_ASAP7_75t_L g3871 ( 
.A(n_3769),
.B(n_284),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_SL g3872 ( 
.A(n_3661),
.B(n_285),
.Y(n_3872)
);

BUFx6f_ASAP7_75t_L g3873 ( 
.A(n_3645),
.Y(n_3873)
);

AND2x4_ASAP7_75t_L g3874 ( 
.A(n_3640),
.B(n_286),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3737),
.B(n_286),
.Y(n_3875)
);

OR2x2_ASAP7_75t_SL g3876 ( 
.A(n_3651),
.B(n_287),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3652),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3642),
.B(n_288),
.Y(n_3878)
);

BUFx3_ASAP7_75t_L g3879 ( 
.A(n_3705),
.Y(n_3879)
);

AOI22xp33_ASAP7_75t_L g3880 ( 
.A1(n_3837),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3746),
.A2(n_289),
.B(n_290),
.Y(n_3881)
);

AOI22xp33_ASAP7_75t_L g3882 ( 
.A1(n_3778),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_3882)
);

O2A1O1Ixp5_ASAP7_75t_L g3883 ( 
.A1(n_3719),
.A2(n_293),
.B(n_291),
.C(n_292),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3655),
.Y(n_3884)
);

INVxp67_ASAP7_75t_SL g3885 ( 
.A(n_3735),
.Y(n_3885)
);

AOI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_3847),
.A2(n_294),
.B(n_295),
.Y(n_3886)
);

CKINVDCx6p67_ASAP7_75t_R g3887 ( 
.A(n_3663),
.Y(n_3887)
);

INVx3_ASAP7_75t_L g3888 ( 
.A(n_3659),
.Y(n_3888)
);

HB1xp67_ASAP7_75t_L g3889 ( 
.A(n_3638),
.Y(n_3889)
);

A2O1A1Ixp33_ASAP7_75t_SL g3890 ( 
.A1(n_3840),
.A2(n_297),
.B(n_294),
.C(n_296),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3677),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3638),
.B(n_296),
.Y(n_3892)
);

A2O1A1Ixp33_ASAP7_75t_L g3893 ( 
.A1(n_3749),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3719),
.A2(n_298),
.B(n_299),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3795),
.B(n_300),
.Y(n_3895)
);

BUFx6f_ASAP7_75t_L g3896 ( 
.A(n_3645),
.Y(n_3896)
);

INVx3_ASAP7_75t_L g3897 ( 
.A(n_3659),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3658),
.B(n_300),
.Y(n_3898)
);

OAI22xp5_ASAP7_75t_L g3899 ( 
.A1(n_3722),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3899)
);

AND2x4_ASAP7_75t_L g3900 ( 
.A(n_3658),
.B(n_3662),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3682),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3750),
.Y(n_3902)
);

BUFx6f_ASAP7_75t_L g3903 ( 
.A(n_3670),
.Y(n_3903)
);

HB1xp67_ASAP7_75t_SL g3904 ( 
.A(n_3647),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3778),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3905)
);

INVx3_ASAP7_75t_L g3906 ( 
.A(n_3659),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3843),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_3907)
);

NAND2xp33_ASAP7_75t_L g3908 ( 
.A(n_3738),
.B(n_304),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3664),
.A2(n_306),
.B(n_308),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3694),
.Y(n_3910)
);

CKINVDCx8_ASAP7_75t_R g3911 ( 
.A(n_3748),
.Y(n_3911)
);

AND2x4_ASAP7_75t_L g3912 ( 
.A(n_3662),
.B(n_308),
.Y(n_3912)
);

A2O1A1Ixp33_ASAP7_75t_L g3913 ( 
.A1(n_3696),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_3913)
);

BUFx4f_ASAP7_75t_L g3914 ( 
.A(n_3670),
.Y(n_3914)
);

BUFx2_ASAP7_75t_L g3915 ( 
.A(n_3750),
.Y(n_3915)
);

INVxp33_ASAP7_75t_L g3916 ( 
.A(n_3791),
.Y(n_3916)
);

BUFx12f_ASAP7_75t_L g3917 ( 
.A(n_3685),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3781),
.B(n_309),
.Y(n_3918)
);

INVx3_ASAP7_75t_L g3919 ( 
.A(n_3675),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3795),
.B(n_311),
.Y(n_3920)
);

NOR2xp33_ASAP7_75t_L g3921 ( 
.A(n_3819),
.B(n_312),
.Y(n_3921)
);

BUFx3_ASAP7_75t_L g3922 ( 
.A(n_3649),
.Y(n_3922)
);

AND2x4_ASAP7_75t_L g3923 ( 
.A(n_3666),
.B(n_312),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3703),
.Y(n_3924)
);

AOI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_3839),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3925)
);

NOR2xp67_ASAP7_75t_L g3926 ( 
.A(n_3657),
.B(n_313),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3723),
.Y(n_3927)
);

INVx3_ASAP7_75t_L g3928 ( 
.A(n_3675),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_3841),
.A2(n_314),
.B(n_317),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3799),
.B(n_317),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3841),
.A2(n_318),
.B(n_319),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3637),
.B(n_318),
.Y(n_3932)
);

AND2x2_ASAP7_75t_L g3933 ( 
.A(n_3795),
.B(n_319),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_SL g3934 ( 
.A(n_3699),
.B(n_320),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3805),
.B(n_321),
.Y(n_3935)
);

AND2x4_ASAP7_75t_L g3936 ( 
.A(n_3666),
.B(n_322),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3697),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3846),
.A2(n_322),
.B(n_323),
.Y(n_3938)
);

NAND2x1p5_ASAP7_75t_L g3939 ( 
.A(n_3675),
.B(n_323),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3776),
.B(n_324),
.Y(n_3940)
);

NAND2x1p5_ASAP7_75t_L g3941 ( 
.A(n_3699),
.B(n_3712),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3770),
.B(n_325),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3772),
.B(n_325),
.Y(n_3943)
);

AOI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_3650),
.A2(n_326),
.B(n_327),
.Y(n_3944)
);

AOI222xp33_ASAP7_75t_L g3945 ( 
.A1(n_3701),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.C1(n_330),
.C2(n_331),
.Y(n_3945)
);

A2O1A1Ixp33_ASAP7_75t_L g3946 ( 
.A1(n_3850),
.A2(n_334),
.B(n_330),
.C(n_332),
.Y(n_3946)
);

AOI21xp5_ASAP7_75t_L g3947 ( 
.A1(n_3851),
.A2(n_332),
.B(n_334),
.Y(n_3947)
);

AND2x4_ASAP7_75t_L g3948 ( 
.A(n_3697),
.B(n_335),
.Y(n_3948)
);

OAI22xp5_ASAP7_75t_L g3949 ( 
.A1(n_3717),
.A2(n_338),
.B1(n_335),
.B2(n_336),
.Y(n_3949)
);

HB1xp67_ASAP7_75t_L g3950 ( 
.A(n_3635),
.Y(n_3950)
);

AND2x4_ASAP7_75t_L g3951 ( 
.A(n_3635),
.B(n_336),
.Y(n_3951)
);

OAI21x1_ASAP7_75t_L g3952 ( 
.A1(n_3678),
.A2(n_338),
.B(n_339),
.Y(n_3952)
);

AOI21xp5_ASAP7_75t_L g3953 ( 
.A1(n_3802),
.A2(n_340),
.B(n_341),
.Y(n_3953)
);

BUFx8_ASAP7_75t_L g3954 ( 
.A(n_3803),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3802),
.A2(n_340),
.B(n_341),
.Y(n_3955)
);

AND2x2_ASAP7_75t_SL g3956 ( 
.A(n_3790),
.B(n_342),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3724),
.Y(n_3957)
);

INVx2_ASAP7_75t_SL g3958 ( 
.A(n_3686),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3774),
.B(n_342),
.Y(n_3959)
);

NAND2x1p5_ASAP7_75t_L g3960 ( 
.A(n_3712),
.B(n_343),
.Y(n_3960)
);

INVx3_ASAP7_75t_SL g3961 ( 
.A(n_3771),
.Y(n_3961)
);

NOR2xp33_ASAP7_75t_L g3962 ( 
.A(n_3794),
.B(n_3791),
.Y(n_3962)
);

CKINVDCx5p33_ASAP7_75t_R g3963 ( 
.A(n_3726),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3838),
.A2(n_343),
.B(n_344),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3811),
.B(n_344),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3838),
.A2(n_345),
.B(n_346),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3763),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3657),
.B(n_347),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3755),
.B(n_348),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3759),
.B(n_348),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3631),
.Y(n_3971)
);

AND2x4_ASAP7_75t_L g3972 ( 
.A(n_3758),
.B(n_349),
.Y(n_3972)
);

NAND2x1p5_ASAP7_75t_L g3973 ( 
.A(n_3712),
.B(n_350),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3639),
.Y(n_3974)
);

OR2x2_ASAP7_75t_L g3975 ( 
.A(n_3787),
.B(n_350),
.Y(n_3975)
);

INVx2_ASAP7_75t_SL g3976 ( 
.A(n_3706),
.Y(n_3976)
);

AOI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3831),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_3977)
);

AOI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3827),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_3978)
);

BUFx12f_ASAP7_75t_L g3979 ( 
.A(n_3798),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3641),
.B(n_354),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3817),
.B(n_356),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3693),
.Y(n_3982)
);

AND2x2_ASAP7_75t_L g3983 ( 
.A(n_3777),
.B(n_356),
.Y(n_3983)
);

OR2x6_ASAP7_75t_L g3984 ( 
.A(n_3644),
.B(n_357),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3710),
.B(n_358),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3729),
.Y(n_3986)
);

INVx3_ASAP7_75t_L g3987 ( 
.A(n_3673),
.Y(n_3987)
);

NOR2xp33_ASAP7_75t_L g3988 ( 
.A(n_3822),
.B(n_358),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3834),
.A2(n_359),
.B(n_360),
.Y(n_3989)
);

INVx3_ASAP7_75t_L g3990 ( 
.A(n_3636),
.Y(n_3990)
);

INVx1_ASAP7_75t_SL g3991 ( 
.A(n_3732),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3777),
.B(n_359),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3720),
.Y(n_3993)
);

NOR2xp33_ASAP7_75t_SL g3994 ( 
.A(n_3633),
.B(n_360),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3788),
.B(n_3779),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3800),
.B(n_361),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3740),
.Y(n_3997)
);

O2A1O1Ixp33_ASAP7_75t_L g3998 ( 
.A1(n_3688),
.A2(n_363),
.B(n_361),
.C(n_362),
.Y(n_3998)
);

AND2x4_ASAP7_75t_L g3999 ( 
.A(n_3632),
.B(n_362),
.Y(n_3999)
);

INVx5_ASAP7_75t_L g4000 ( 
.A(n_3644),
.Y(n_4000)
);

CKINVDCx6p67_ASAP7_75t_R g4001 ( 
.A(n_3798),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3800),
.B(n_363),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3812),
.B(n_364),
.Y(n_4003)
);

OAI321xp33_ASAP7_75t_L g4004 ( 
.A1(n_3757),
.A2(n_365),
.A3(n_366),
.B1(n_367),
.B2(n_368),
.C(n_369),
.Y(n_4004)
);

OR2x2_ASAP7_75t_L g4005 ( 
.A(n_3793),
.B(n_365),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3654),
.Y(n_4006)
);

INVx4_ASAP7_75t_L g4007 ( 
.A(n_3657),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3654),
.Y(n_4008)
);

O2A1O1Ixp33_ASAP7_75t_L g4009 ( 
.A1(n_3751),
.A2(n_370),
.B(n_366),
.C(n_369),
.Y(n_4009)
);

AND2x4_ASAP7_75t_L g4010 ( 
.A(n_3632),
.B(n_370),
.Y(n_4010)
);

INVx2_ASAP7_75t_L g4011 ( 
.A(n_3656),
.Y(n_4011)
);

HB1xp67_ASAP7_75t_L g4012 ( 
.A(n_3780),
.Y(n_4012)
);

INVx2_ASAP7_75t_SL g4013 ( 
.A(n_3721),
.Y(n_4013)
);

BUFx6f_ASAP7_75t_L g4014 ( 
.A(n_3684),
.Y(n_4014)
);

NOR2x1_ASAP7_75t_SL g4015 ( 
.A(n_3765),
.B(n_371),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_3656),
.Y(n_4016)
);

AOI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_3672),
.A2(n_371),
.B(n_373),
.Y(n_4017)
);

INVx3_ASAP7_75t_SL g4018 ( 
.A(n_3858),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3754),
.B(n_373),
.Y(n_4019)
);

AOI22xp5_ASAP7_75t_L g4020 ( 
.A1(n_3761),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3808),
.A2(n_374),
.B(n_375),
.Y(n_4021)
);

BUFx3_ASAP7_75t_L g4022 ( 
.A(n_3643),
.Y(n_4022)
);

BUFx8_ASAP7_75t_SL g4023 ( 
.A(n_3821),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3806),
.Y(n_4024)
);

CKINVDCx5p33_ASAP7_75t_R g4025 ( 
.A(n_3773),
.Y(n_4025)
);

INVx3_ASAP7_75t_L g4026 ( 
.A(n_3636),
.Y(n_4026)
);

AND2x4_ASAP7_75t_L g4027 ( 
.A(n_3788),
.B(n_376),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3825),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3782),
.B(n_377),
.Y(n_4029)
);

INVx3_ASAP7_75t_L g4030 ( 
.A(n_3633),
.Y(n_4030)
);

AOI21xp5_ASAP7_75t_L g4031 ( 
.A1(n_3832),
.A2(n_378),
.B(n_379),
.Y(n_4031)
);

HB1xp67_ASAP7_75t_L g4032 ( 
.A(n_3853),
.Y(n_4032)
);

AOI21xp5_ASAP7_75t_L g4033 ( 
.A1(n_3832),
.A2(n_378),
.B(n_380),
.Y(n_4033)
);

O2A1O1Ixp5_ASAP7_75t_L g4034 ( 
.A1(n_3704),
.A2(n_382),
.B(n_380),
.C(n_381),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_SL g4035 ( 
.A(n_3818),
.B(n_381),
.Y(n_4035)
);

OAI22xp33_ASAP7_75t_L g4036 ( 
.A1(n_3765),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_3810),
.B(n_385),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3768),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3669),
.B(n_385),
.Y(n_4039)
);

INVx4_ASAP7_75t_L g4040 ( 
.A(n_3979),
.Y(n_4040)
);

BUFx2_ASAP7_75t_R g4041 ( 
.A(n_4023),
.Y(n_4041)
);

OAI21xp5_ASAP7_75t_SL g4042 ( 
.A1(n_3945),
.A2(n_3766),
.B(n_3702),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3865),
.Y(n_4043)
);

BUFx6f_ASAP7_75t_L g4044 ( 
.A(n_3873),
.Y(n_4044)
);

OAI22xp5_ASAP7_75t_L g4045 ( 
.A1(n_4020),
.A2(n_3913),
.B1(n_3700),
.B2(n_3835),
.Y(n_4045)
);

INVx6_ASAP7_75t_L g4046 ( 
.A(n_3954),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3908),
.A2(n_3852),
.B1(n_3790),
.B2(n_3854),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3915),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3877),
.Y(n_4049)
);

BUFx2_ASAP7_75t_L g4050 ( 
.A(n_3900),
.Y(n_4050)
);

BUFx8_ASAP7_75t_L g4051 ( 
.A(n_3879),
.Y(n_4051)
);

CKINVDCx11_ASAP7_75t_R g4052 ( 
.A(n_3911),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3884),
.Y(n_4053)
);

INVx3_ASAP7_75t_L g4054 ( 
.A(n_3900),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3864),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3891),
.Y(n_4056)
);

AOI22xp33_ASAP7_75t_L g4057 ( 
.A1(n_3886),
.A2(n_3854),
.B1(n_3855),
.B2(n_3849),
.Y(n_4057)
);

AOI22xp33_ASAP7_75t_SL g4058 ( 
.A1(n_3956),
.A2(n_3809),
.B1(n_3797),
.B2(n_3783),
.Y(n_4058)
);

BUFx4f_ASAP7_75t_L g4059 ( 
.A(n_3871),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_L g4060 ( 
.A1(n_3881),
.A2(n_3745),
.B1(n_3833),
.B2(n_3784),
.Y(n_4060)
);

BUFx2_ASAP7_75t_SL g4061 ( 
.A(n_3958),
.Y(n_4061)
);

OAI221xp5_ASAP7_75t_L g4062 ( 
.A1(n_3978),
.A2(n_3695),
.B1(n_3764),
.B2(n_3736),
.C(n_3801),
.Y(n_4062)
);

BUFx4f_ASAP7_75t_SL g4063 ( 
.A(n_3917),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_SL g4064 ( 
.A1(n_4015),
.A2(n_3809),
.B1(n_3797),
.B2(n_3783),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3902),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_4032),
.B(n_3829),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3909),
.A2(n_3826),
.B1(n_3828),
.B2(n_3753),
.Y(n_4067)
);

INVx1_ASAP7_75t_SL g4068 ( 
.A(n_4001),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3901),
.Y(n_4069)
);

AOI22xp33_ASAP7_75t_L g4070 ( 
.A1(n_3947),
.A2(n_3826),
.B1(n_3828),
.B2(n_3807),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3984),
.A2(n_3785),
.B1(n_3844),
.B2(n_3752),
.Y(n_4071)
);

BUFx4f_ASAP7_75t_L g4072 ( 
.A(n_3871),
.Y(n_4072)
);

AOI22xp33_ASAP7_75t_L g4073 ( 
.A1(n_3967),
.A2(n_3828),
.B1(n_3826),
.B2(n_3731),
.Y(n_4073)
);

AOI22xp5_ASAP7_75t_SL g4074 ( 
.A1(n_3868),
.A2(n_3738),
.B1(n_3713),
.B2(n_3836),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3910),
.Y(n_4075)
);

INVx4_ASAP7_75t_L g4076 ( 
.A(n_4007),
.Y(n_4076)
);

INVx6_ASAP7_75t_L g4077 ( 
.A(n_3954),
.Y(n_4077)
);

CKINVDCx5p33_ASAP7_75t_R g4078 ( 
.A(n_3904),
.Y(n_4078)
);

INVx6_ASAP7_75t_L g4079 ( 
.A(n_3922),
.Y(n_4079)
);

BUFx10_ASAP7_75t_L g4080 ( 
.A(n_3921),
.Y(n_4080)
);

INVx4_ASAP7_75t_L g4081 ( 
.A(n_4007),
.Y(n_4081)
);

INVx4_ASAP7_75t_L g4082 ( 
.A(n_3887),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3924),
.Y(n_4083)
);

BUFx2_ASAP7_75t_L g4084 ( 
.A(n_3889),
.Y(n_4084)
);

INVx1_ASAP7_75t_SL g4085 ( 
.A(n_3961),
.Y(n_4085)
);

INVx4_ASAP7_75t_L g4086 ( 
.A(n_4018),
.Y(n_4086)
);

INVx4_ASAP7_75t_L g4087 ( 
.A(n_3984),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3937),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3927),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3863),
.A2(n_3733),
.B1(n_3845),
.B2(n_3824),
.Y(n_4090)
);

OAI22xp5_ASAP7_75t_L g4091 ( 
.A1(n_3925),
.A2(n_3708),
.B1(n_3848),
.B2(n_3804),
.Y(n_4091)
);

BUFx3_ASAP7_75t_L g4092 ( 
.A(n_3859),
.Y(n_4092)
);

OAI22xp33_ASAP7_75t_L g4093 ( 
.A1(n_3994),
.A2(n_3830),
.B1(n_3813),
.B2(n_3856),
.Y(n_4093)
);

AOI21xp33_ASAP7_75t_L g4094 ( 
.A1(n_3890),
.A2(n_3814),
.B(n_3760),
.Y(n_4094)
);

CKINVDCx11_ASAP7_75t_R g4095 ( 
.A(n_3991),
.Y(n_4095)
);

INVx1_ASAP7_75t_SL g4096 ( 
.A(n_3963),
.Y(n_4096)
);

AOI22xp33_ASAP7_75t_L g4097 ( 
.A1(n_3899),
.A2(n_3816),
.B1(n_3815),
.B2(n_3738),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3950),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3957),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_4011),
.B(n_4016),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3860),
.Y(n_4101)
);

INVx6_ASAP7_75t_L g4102 ( 
.A(n_3873),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3867),
.Y(n_4103)
);

BUFx3_ASAP7_75t_L g4104 ( 
.A(n_4022),
.Y(n_4104)
);

INVx8_ASAP7_75t_L g4105 ( 
.A(n_4027),
.Y(n_4105)
);

BUFx8_ASAP7_75t_L g4106 ( 
.A(n_3895),
.Y(n_4106)
);

AOI22xp33_ASAP7_75t_SL g4107 ( 
.A1(n_3949),
.A2(n_3804),
.B1(n_3830),
.B2(n_3739),
.Y(n_4107)
);

CKINVDCx20_ASAP7_75t_R g4108 ( 
.A(n_4025),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_L g4109 ( 
.A1(n_3880),
.A2(n_3842),
.B1(n_3792),
.B2(n_3646),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_4006),
.Y(n_4110)
);

INVx1_ASAP7_75t_SL g4111 ( 
.A(n_3976),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3885),
.B(n_3691),
.Y(n_4112)
);

OAI22xp5_ASAP7_75t_L g4113 ( 
.A1(n_3907),
.A2(n_3683),
.B1(n_3653),
.B2(n_3676),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3894),
.A2(n_3796),
.B1(n_3698),
.B2(n_3676),
.Y(n_4114)
);

BUFx2_ASAP7_75t_SL g4115 ( 
.A(n_3926),
.Y(n_4115)
);

AOI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_4036),
.A2(n_3893),
.B1(n_3872),
.B2(n_3946),
.Y(n_4116)
);

CKINVDCx11_ASAP7_75t_R g4117 ( 
.A(n_3873),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_4008),
.Y(n_4118)
);

AOI22xp33_ASAP7_75t_L g4119 ( 
.A1(n_4017),
.A2(n_3789),
.B1(n_3786),
.B2(n_3715),
.Y(n_4119)
);

AOI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_3951),
.A2(n_3789),
.B1(n_3786),
.B2(n_3857),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_SL g4121 ( 
.A1(n_4000),
.A2(n_3742),
.B1(n_3741),
.B2(n_3711),
.Y(n_4121)
);

OAI21xp5_ASAP7_75t_SL g4122 ( 
.A1(n_3953),
.A2(n_3744),
.B(n_3820),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_SL g4123 ( 
.A1(n_4000),
.A2(n_3742),
.B1(n_3741),
.B2(n_3711),
.Y(n_4123)
);

AOI22xp33_ASAP7_75t_L g4124 ( 
.A1(n_3938),
.A2(n_3725),
.B1(n_3716),
.B2(n_3665),
.Y(n_4124)
);

BUFx8_ASAP7_75t_SL g4125 ( 
.A(n_3914),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_3929),
.A2(n_3687),
.B1(n_3747),
.B2(n_3668),
.Y(n_4126)
);

OAI22xp5_ASAP7_75t_L g4127 ( 
.A1(n_3882),
.A2(n_3744),
.B1(n_3671),
.B2(n_3728),
.Y(n_4127)
);

AOI22xp33_ASAP7_75t_L g4128 ( 
.A1(n_3931),
.A2(n_3767),
.B1(n_3743),
.B2(n_3707),
.Y(n_4128)
);

INVx3_ASAP7_75t_L g4129 ( 
.A(n_3990),
.Y(n_4129)
);

OAI22xp5_ASAP7_75t_L g4130 ( 
.A1(n_3905),
.A2(n_3762),
.B1(n_3775),
.B2(n_3820),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3869),
.Y(n_4131)
);

INVx1_ASAP7_75t_SL g4132 ( 
.A(n_3995),
.Y(n_4132)
);

OAI22xp5_ASAP7_75t_L g4133 ( 
.A1(n_3977),
.A2(n_3756),
.B1(n_3709),
.B2(n_3718),
.Y(n_4133)
);

AOI22xp33_ASAP7_75t_SL g4134 ( 
.A1(n_4000),
.A2(n_3711),
.B1(n_3756),
.B2(n_3692),
.Y(n_4134)
);

CKINVDCx11_ASAP7_75t_R g4135 ( 
.A(n_3896),
.Y(n_4135)
);

HB1xp67_ASAP7_75t_L g4136 ( 
.A(n_4012),
.Y(n_4136)
);

BUFx4f_ASAP7_75t_SL g4137 ( 
.A(n_4013),
.Y(n_4137)
);

OAI22xp5_ASAP7_75t_SL g4138 ( 
.A1(n_3876),
.A2(n_3679),
.B1(n_3756),
.B2(n_3773),
.Y(n_4138)
);

INVx6_ASAP7_75t_L g4139 ( 
.A(n_3896),
.Y(n_4139)
);

INVx5_ASAP7_75t_L g4140 ( 
.A(n_3862),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_L g4141 ( 
.A1(n_4021),
.A2(n_3674),
.B1(n_3667),
.B2(n_3727),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_3971),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3974),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3982),
.Y(n_4144)
);

BUFx10_ASAP7_75t_L g4145 ( 
.A(n_3988),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3993),
.Y(n_4146)
);

OAI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_3944),
.A2(n_3730),
.B1(n_3689),
.B2(n_3690),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_3990),
.B(n_3684),
.Y(n_4148)
);

INVx3_ASAP7_75t_L g4149 ( 
.A(n_4026),
.Y(n_4149)
);

OAI22xp5_ASAP7_75t_L g4150 ( 
.A1(n_3955),
.A2(n_3690),
.B1(n_3734),
.B2(n_3689),
.Y(n_4150)
);

NOR2xp33_ASAP7_75t_L g4151 ( 
.A(n_3916),
.B(n_3734),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4026),
.B(n_3721),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3986),
.Y(n_4153)
);

AOI22xp33_ASAP7_75t_L g4154 ( 
.A1(n_3866),
.A2(n_389),
.B1(n_386),
.B2(n_388),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4024),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4028),
.Y(n_4156)
);

CKINVDCx6p67_ASAP7_75t_R g4157 ( 
.A(n_3920),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_3962),
.B(n_389),
.Y(n_4158)
);

INVx6_ASAP7_75t_L g4159 ( 
.A(n_3896),
.Y(n_4159)
);

INVx4_ASAP7_75t_L g4160 ( 
.A(n_3898),
.Y(n_4160)
);

OAI22xp5_ASAP7_75t_L g4161 ( 
.A1(n_3964),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_4161)
);

BUFx10_ASAP7_75t_L g4162 ( 
.A(n_4027),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3997),
.Y(n_4163)
);

BUFx4f_ASAP7_75t_L g4164 ( 
.A(n_3903),
.Y(n_4164)
);

HB1xp67_ASAP7_75t_L g4165 ( 
.A(n_4038),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_3888),
.Y(n_4166)
);

INVx6_ASAP7_75t_L g4167 ( 
.A(n_3903),
.Y(n_4167)
);

CKINVDCx8_ASAP7_75t_R g4168 ( 
.A(n_3903),
.Y(n_4168)
);

OAI22xp5_ASAP7_75t_L g4169 ( 
.A1(n_3966),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_4169)
);

BUFx3_ASAP7_75t_L g4170 ( 
.A(n_4014),
.Y(n_4170)
);

INVx2_ASAP7_75t_L g4171 ( 
.A(n_3888),
.Y(n_4171)
);

AOI22xp33_ASAP7_75t_L g4172 ( 
.A1(n_3989),
.A2(n_4033),
.B1(n_4031),
.B2(n_3951),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_3897),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_L g4174 ( 
.A1(n_3999),
.A2(n_397),
.B1(n_393),
.B2(n_396),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3975),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4005),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_3999),
.A2(n_397),
.B1(n_393),
.B2(n_396),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3861),
.Y(n_4178)
);

BUFx4_ASAP7_75t_SL g4179 ( 
.A(n_3960),
.Y(n_4179)
);

OAI22xp5_ASAP7_75t_L g4180 ( 
.A1(n_3939),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_4180)
);

BUFx8_ASAP7_75t_SL g4181 ( 
.A(n_3874),
.Y(n_4181)
);

BUFx12f_ASAP7_75t_L g4182 ( 
.A(n_3940),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_SL g4183 ( 
.A1(n_3933),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_4183)
);

OAI22x1_ASAP7_75t_L g4184 ( 
.A1(n_3874),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_4184)
);

CKINVDCx20_ASAP7_75t_R g4185 ( 
.A(n_3987),
.Y(n_4185)
);

CKINVDCx11_ASAP7_75t_R g4186 ( 
.A(n_4014),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3897),
.Y(n_4187)
);

CKINVDCx11_ASAP7_75t_R g4188 ( 
.A(n_4014),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3906),
.Y(n_4189)
);

BUFx4_ASAP7_75t_R g4190 ( 
.A(n_3973),
.Y(n_4190)
);

INVx5_ASAP7_75t_L g4191 ( 
.A(n_3862),
.Y(n_4191)
);

OR2x6_ASAP7_75t_L g4192 ( 
.A(n_4061),
.B(n_3941),
.Y(n_4192)
);

INVxp67_ASAP7_75t_L g4193 ( 
.A(n_4136),
.Y(n_4193)
);

AOI22xp33_ASAP7_75t_L g4194 ( 
.A1(n_4045),
.A2(n_4035),
.B1(n_3968),
.B2(n_3934),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4155),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_4166),
.Y(n_4196)
);

BUFx3_ASAP7_75t_L g4197 ( 
.A(n_4051),
.Y(n_4197)
);

AO21x2_ASAP7_75t_L g4198 ( 
.A1(n_4187),
.A2(n_3870),
.B(n_3878),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4156),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_4121),
.A2(n_3998),
.B1(n_4009),
.B2(n_3898),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4043),
.Y(n_4201)
);

AOI22xp33_ASAP7_75t_L g4202 ( 
.A1(n_4071),
.A2(n_4037),
.B1(n_4019),
.B2(n_3932),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4171),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_SL g4204 ( 
.A(n_4086),
.B(n_4030),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4049),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_4050),
.B(n_3906),
.Y(n_4206)
);

INVx3_ASAP7_75t_L g4207 ( 
.A(n_4086),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4053),
.Y(n_4208)
);

NAND2x1p5_ASAP7_75t_L g4209 ( 
.A(n_4140),
.B(n_3919),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_4173),
.Y(n_4210)
);

INVx3_ASAP7_75t_L g4211 ( 
.A(n_4076),
.Y(n_4211)
);

HB1xp67_ASAP7_75t_L g4212 ( 
.A(n_4066),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4142),
.B(n_4003),
.Y(n_4213)
);

HB1xp67_ASAP7_75t_L g4214 ( 
.A(n_4165),
.Y(n_4214)
);

BUFx6f_ASAP7_75t_L g4215 ( 
.A(n_4046),
.Y(n_4215)
);

AOI22xp33_ASAP7_75t_L g4216 ( 
.A1(n_4097),
.A2(n_4039),
.B1(n_4010),
.B2(n_3972),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4056),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_4189),
.Y(n_4218)
);

AOI21x1_ASAP7_75t_L g4219 ( 
.A1(n_4150),
.A2(n_3918),
.B(n_3875),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4069),
.Y(n_4220)
);

NAND2x1p5_ASAP7_75t_L g4221 ( 
.A(n_4140),
.B(n_3919),
.Y(n_4221)
);

AO21x2_ASAP7_75t_L g4222 ( 
.A1(n_4122),
.A2(n_3969),
.B(n_3959),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4075),
.Y(n_4223)
);

INVx2_ASAP7_75t_R g4224 ( 
.A(n_4140),
.Y(n_4224)
);

BUFx2_ASAP7_75t_L g4225 ( 
.A(n_4084),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4083),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_4054),
.B(n_3928),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4089),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_SL g4229 ( 
.A1(n_4074),
.A2(n_3892),
.B1(n_3923),
.B2(n_3912),
.Y(n_4229)
);

AOI22xp33_ASAP7_75t_L g4230 ( 
.A1(n_4062),
.A2(n_4010),
.B1(n_3972),
.B2(n_3952),
.Y(n_4230)
);

OA21x2_ASAP7_75t_L g4231 ( 
.A1(n_4110),
.A2(n_3883),
.B(n_3970),
.Y(n_4231)
);

AO21x2_ASAP7_75t_L g4232 ( 
.A1(n_4094),
.A2(n_3981),
.B(n_3935),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4054),
.B(n_4132),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_4148),
.B(n_3928),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4099),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4098),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_4118),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_4129),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4143),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4144),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4146),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_4100),
.B(n_4030),
.Y(n_4242)
);

BUFx6f_ASAP7_75t_L g4243 ( 
.A(n_4046),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4101),
.Y(n_4244)
);

INVx3_ASAP7_75t_L g4245 ( 
.A(n_4076),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4103),
.Y(n_4246)
);

INVx2_ASAP7_75t_SL g4247 ( 
.A(n_4079),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4131),
.Y(n_4248)
);

HB1xp67_ASAP7_75t_L g4249 ( 
.A(n_4153),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4175),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4176),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4178),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_4052),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4163),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4055),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_4129),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4065),
.Y(n_4257)
);

OAI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_4067),
.A2(n_4034),
.B(n_4004),
.Y(n_4258)
);

INVx2_ASAP7_75t_SL g4259 ( 
.A(n_4079),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4048),
.B(n_3912),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4088),
.Y(n_4261)
);

BUFx4f_ASAP7_75t_SL g4262 ( 
.A(n_4051),
.Y(n_4262)
);

INVx3_ASAP7_75t_L g4263 ( 
.A(n_4081),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4112),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4149),
.Y(n_4265)
);

OAI21x1_ASAP7_75t_L g4266 ( 
.A1(n_4149),
.A2(n_3985),
.B(n_3980),
.Y(n_4266)
);

BUFx2_ASAP7_75t_L g4267 ( 
.A(n_4185),
.Y(n_4267)
);

INVxp67_ASAP7_75t_L g4268 ( 
.A(n_4115),
.Y(n_4268)
);

BUFx10_ASAP7_75t_L g4269 ( 
.A(n_4077),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4160),
.Y(n_4270)
);

AOI22xp33_ASAP7_75t_L g4271 ( 
.A1(n_4060),
.A2(n_4002),
.B1(n_3996),
.B2(n_3936),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4152),
.B(n_3923),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4160),
.Y(n_4273)
);

OR2x6_ASAP7_75t_L g4274 ( 
.A(n_4087),
.B(n_3936),
.Y(n_4274)
);

CKINVDCx20_ASAP7_75t_R g4275 ( 
.A(n_4095),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4081),
.Y(n_4276)
);

NAND2x1p5_ASAP7_75t_L g4277 ( 
.A(n_4191),
.B(n_3948),
.Y(n_4277)
);

BUFx8_ASAP7_75t_SL g4278 ( 
.A(n_4078),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4170),
.Y(n_4279)
);

HB1xp67_ASAP7_75t_L g4280 ( 
.A(n_4191),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4044),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_4044),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_4044),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4191),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4102),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4102),
.Y(n_4286)
);

AO21x1_ASAP7_75t_SL g4287 ( 
.A1(n_4047),
.A2(n_3943),
.B(n_3942),
.Y(n_4287)
);

BUFx6f_ASAP7_75t_L g4288 ( 
.A(n_4077),
.Y(n_4288)
);

INVx3_ASAP7_75t_L g4289 ( 
.A(n_4162),
.Y(n_4289)
);

BUFx2_ASAP7_75t_L g4290 ( 
.A(n_4087),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4139),
.Y(n_4291)
);

AND2x4_ASAP7_75t_L g4292 ( 
.A(n_4082),
.B(n_3948),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4139),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4159),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4134),
.B(n_3930),
.Y(n_4295)
);

HB1xp67_ASAP7_75t_L g4296 ( 
.A(n_4111),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4159),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4167),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_4162),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4167),
.Y(n_4300)
);

AND2x2_ASAP7_75t_L g4301 ( 
.A(n_4157),
.B(n_3983),
.Y(n_4301)
);

AOI22xp5_ASAP7_75t_L g4302 ( 
.A1(n_4138),
.A2(n_4042),
.B1(n_4116),
.B2(n_4072),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4151),
.Y(n_4303)
);

OAI22xp33_ASAP7_75t_L g4304 ( 
.A1(n_4059),
.A2(n_3992),
.B1(n_4029),
.B2(n_3965),
.Y(n_4304)
);

INVx2_ASAP7_75t_SL g4305 ( 
.A(n_4105),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4105),
.Y(n_4306)
);

INVx1_ASAP7_75t_SL g4307 ( 
.A(n_4190),
.Y(n_4307)
);

OAI22xp33_ASAP7_75t_L g4308 ( 
.A1(n_4059),
.A2(n_633),
.B1(n_406),
.B2(n_404),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4104),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4123),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4168),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4120),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4106),
.Y(n_4313)
);

NAND2x1p5_ASAP7_75t_L g4314 ( 
.A(n_4072),
.B(n_405),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4106),
.Y(n_4315)
);

HB1xp67_ASAP7_75t_L g4316 ( 
.A(n_4181),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4130),
.Y(n_4317)
);

CKINVDCx5p33_ASAP7_75t_R g4318 ( 
.A(n_4125),
.Y(n_4318)
);

AND2x4_ASAP7_75t_L g4319 ( 
.A(n_4082),
.B(n_405),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4127),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4068),
.B(n_407),
.Y(n_4321)
);

INVx3_ASAP7_75t_L g4322 ( 
.A(n_4040),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4092),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4158),
.Y(n_4324)
);

OR2x6_ASAP7_75t_L g4325 ( 
.A(n_4040),
.B(n_4182),
.Y(n_4325)
);

AND2x4_ASAP7_75t_L g4326 ( 
.A(n_4085),
.B(n_408),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4147),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4080),
.Y(n_4328)
);

INVx3_ASAP7_75t_L g4329 ( 
.A(n_4117),
.Y(n_4329)
);

HB1xp67_ASAP7_75t_L g4330 ( 
.A(n_4179),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4080),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4184),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4126),
.Y(n_4333)
);

BUFx4f_ASAP7_75t_SL g4334 ( 
.A(n_4108),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4135),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_4124),
.B(n_408),
.Y(n_4336)
);

OAI21x1_ASAP7_75t_L g4337 ( 
.A1(n_4128),
.A2(n_409),
.B(n_410),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4057),
.B(n_4141),
.Y(n_4338)
);

AO21x1_ASAP7_75t_L g4339 ( 
.A1(n_4310),
.A2(n_4093),
.B(n_4091),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4239),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4222),
.B(n_4232),
.Y(n_4341)
);

OR2x2_ASAP7_75t_L g4342 ( 
.A(n_4320),
.B(n_4119),
.Y(n_4342)
);

HB1xp67_ASAP7_75t_L g4343 ( 
.A(n_4214),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4192),
.B(n_4186),
.Y(n_4344)
);

OAI21x1_ASAP7_75t_L g4345 ( 
.A1(n_4209),
.A2(n_4172),
.B(n_4114),
.Y(n_4345)
);

AO21x2_ASAP7_75t_L g4346 ( 
.A1(n_4280),
.A2(n_4169),
.B(n_4161),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4218),
.Y(n_4347)
);

NAND2x1_ASAP7_75t_L g4348 ( 
.A(n_4192),
.B(n_4041),
.Y(n_4348)
);

HB1xp67_ASAP7_75t_L g4349 ( 
.A(n_4214),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4196),
.Y(n_4350)
);

OA21x2_ASAP7_75t_L g4351 ( 
.A1(n_4280),
.A2(n_4070),
.B(n_4090),
.Y(n_4351)
);

AND2x4_ASAP7_75t_L g4352 ( 
.A(n_4192),
.B(n_4096),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_4203),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4240),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4210),
.Y(n_4355)
);

OAI21xp5_ASAP7_75t_L g4356 ( 
.A1(n_4302),
.A2(n_4107),
.B(n_4073),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_4290),
.B(n_4270),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4273),
.B(n_4188),
.Y(n_4358)
);

OA21x2_ASAP7_75t_L g4359 ( 
.A1(n_4284),
.A2(n_4109),
.B(n_4154),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4225),
.Y(n_4360)
);

INVx2_ASAP7_75t_SL g4361 ( 
.A(n_4269),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4241),
.Y(n_4362)
);

OA21x2_ASAP7_75t_L g4363 ( 
.A1(n_4268),
.A2(n_4133),
.B(n_4113),
.Y(n_4363)
);

OR2x2_ASAP7_75t_L g4364 ( 
.A(n_4264),
.B(n_4058),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4195),
.Y(n_4365)
);

INVx4_ASAP7_75t_SL g4366 ( 
.A(n_4262),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4199),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4201),
.Y(n_4368)
);

BUFx6f_ASAP7_75t_L g4369 ( 
.A(n_4215),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4237),
.Y(n_4370)
);

HB1xp67_ASAP7_75t_L g4371 ( 
.A(n_4249),
.Y(n_4371)
);

OAI21x1_ASAP7_75t_L g4372 ( 
.A1(n_4209),
.A2(n_4180),
.B(n_4177),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4205),
.Y(n_4373)
);

INVx2_ASAP7_75t_SL g4374 ( 
.A(n_4269),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4208),
.Y(n_4375)
);

AOI22xp33_ASAP7_75t_L g4376 ( 
.A1(n_4333),
.A2(n_4183),
.B1(n_4064),
.B2(n_4174),
.Y(n_4376)
);

BUFx3_ASAP7_75t_L g4377 ( 
.A(n_4262),
.Y(n_4377)
);

AND2x2_ASAP7_75t_L g4378 ( 
.A(n_4206),
.B(n_4145),
.Y(n_4378)
);

NOR2x1_ASAP7_75t_L g4379 ( 
.A(n_4207),
.B(n_4063),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4233),
.B(n_4145),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4217),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4220),
.Y(n_4382)
);

INVxp67_ASAP7_75t_SL g4383 ( 
.A(n_4193),
.Y(n_4383)
);

OR2x2_ASAP7_75t_L g4384 ( 
.A(n_4317),
.B(n_409),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4223),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4226),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_4228),
.Y(n_4387)
);

AOI21x1_ASAP7_75t_L g4388 ( 
.A1(n_4330),
.A2(n_4137),
.B(n_4164),
.Y(n_4388)
);

INVx2_ASAP7_75t_SL g4389 ( 
.A(n_4329),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4234),
.B(n_410),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4235),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_4244),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4246),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4248),
.Y(n_4394)
);

INVx3_ASAP7_75t_L g4395 ( 
.A(n_4221),
.Y(n_4395)
);

OR2x6_ASAP7_75t_L g4396 ( 
.A(n_4268),
.B(n_411),
.Y(n_4396)
);

OR2x2_ASAP7_75t_L g4397 ( 
.A(n_4198),
.B(n_411),
.Y(n_4397)
);

HB1xp67_ASAP7_75t_L g4398 ( 
.A(n_4249),
.Y(n_4398)
);

AO21x2_ASAP7_75t_L g4399 ( 
.A1(n_4204),
.A2(n_413),
.B(n_414),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_4236),
.Y(n_4400)
);

INVx2_ASAP7_75t_SL g4401 ( 
.A(n_4329),
.Y(n_4401)
);

OA21x2_ASAP7_75t_L g4402 ( 
.A1(n_4338),
.A2(n_414),
.B(n_416),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4252),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_4266),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4250),
.Y(n_4405)
);

HB1xp67_ASAP7_75t_L g4406 ( 
.A(n_4193),
.Y(n_4406)
);

OR2x2_ASAP7_75t_L g4407 ( 
.A(n_4198),
.B(n_417),
.Y(n_4407)
);

OA21x2_ASAP7_75t_L g4408 ( 
.A1(n_4338),
.A2(n_417),
.B(n_418),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4251),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4254),
.Y(n_4410)
);

BUFx3_ASAP7_75t_L g4411 ( 
.A(n_4197),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4296),
.Y(n_4412)
);

BUFx3_ASAP7_75t_L g4413 ( 
.A(n_4215),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4296),
.Y(n_4414)
);

INVx2_ASAP7_75t_L g4415 ( 
.A(n_4257),
.Y(n_4415)
);

INVx2_ASAP7_75t_SL g4416 ( 
.A(n_4215),
.Y(n_4416)
);

AO21x2_ASAP7_75t_L g4417 ( 
.A1(n_4295),
.A2(n_418),
.B(n_419),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4213),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4213),
.Y(n_4419)
);

OR2x2_ASAP7_75t_L g4420 ( 
.A(n_4312),
.B(n_419),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4261),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4255),
.Y(n_4422)
);

HB1xp67_ASAP7_75t_L g4423 ( 
.A(n_4212),
.Y(n_4423)
);

AND2x4_ASAP7_75t_L g4424 ( 
.A(n_4207),
.B(n_420),
.Y(n_4424)
);

AO21x2_ASAP7_75t_L g4425 ( 
.A1(n_4295),
.A2(n_4336),
.B(n_4308),
.Y(n_4425)
);

HB1xp67_ASAP7_75t_L g4426 ( 
.A(n_4212),
.Y(n_4426)
);

OA21x2_ASAP7_75t_L g4427 ( 
.A1(n_4258),
.A2(n_421),
.B(n_422),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4231),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4231),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4299),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4238),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4289),
.Y(n_4432)
);

AO21x2_ASAP7_75t_L g4433 ( 
.A1(n_4336),
.A2(n_421),
.B(n_423),
.Y(n_4433)
);

INVx3_ASAP7_75t_L g4434 ( 
.A(n_4221),
.Y(n_4434)
);

HB1xp67_ASAP7_75t_L g4435 ( 
.A(n_4232),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4256),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4289),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4227),
.B(n_423),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_4265),
.Y(n_4439)
);

AND2x2_ASAP7_75t_L g4440 ( 
.A(n_4307),
.B(n_424),
.Y(n_4440)
);

BUFx2_ASAP7_75t_L g4441 ( 
.A(n_4330),
.Y(n_4441)
);

HB1xp67_ASAP7_75t_L g4442 ( 
.A(n_4222),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_4276),
.Y(n_4443)
);

INVx3_ASAP7_75t_L g4444 ( 
.A(n_4243),
.Y(n_4444)
);

INVx2_ASAP7_75t_L g4445 ( 
.A(n_4281),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4282),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4283),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4328),
.Y(n_4448)
);

BUFx3_ASAP7_75t_L g4449 ( 
.A(n_4243),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_4331),
.Y(n_4450)
);

OR2x2_ASAP7_75t_L g4451 ( 
.A(n_4327),
.B(n_424),
.Y(n_4451)
);

BUFx6f_ASAP7_75t_L g4452 ( 
.A(n_4243),
.Y(n_4452)
);

BUFx6f_ASAP7_75t_L g4453 ( 
.A(n_4288),
.Y(n_4453)
);

INVxp67_ASAP7_75t_L g4454 ( 
.A(n_4287),
.Y(n_4454)
);

HB1xp67_ASAP7_75t_L g4455 ( 
.A(n_4224),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4219),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4307),
.B(n_425),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4332),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_4277),
.Y(n_4459)
);

INVx3_ASAP7_75t_L g4460 ( 
.A(n_4288),
.Y(n_4460)
);

AOI21x1_ASAP7_75t_L g4461 ( 
.A1(n_4316),
.A2(n_425),
.B(n_426),
.Y(n_4461)
);

HB1xp67_ASAP7_75t_L g4462 ( 
.A(n_4224),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4211),
.Y(n_4463)
);

BUFx3_ASAP7_75t_L g4464 ( 
.A(n_4288),
.Y(n_4464)
);

INVxp67_ASAP7_75t_SL g4465 ( 
.A(n_4277),
.Y(n_4465)
);

AND2x4_ASAP7_75t_L g4466 ( 
.A(n_4211),
.B(n_427),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4245),
.Y(n_4467)
);

AND2x4_ASAP7_75t_L g4468 ( 
.A(n_4245),
.B(n_427),
.Y(n_4468)
);

INVx3_ASAP7_75t_L g4469 ( 
.A(n_4322),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4263),
.Y(n_4470)
);

AO21x1_ASAP7_75t_SL g4471 ( 
.A1(n_4316),
.A2(n_428),
.B(n_430),
.Y(n_4471)
);

OA21x2_ASAP7_75t_L g4472 ( 
.A1(n_4258),
.A2(n_428),
.B(n_430),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4263),
.Y(n_4473)
);

INVx3_ASAP7_75t_L g4474 ( 
.A(n_4322),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4324),
.Y(n_4475)
);

AO31x2_ASAP7_75t_L g4476 ( 
.A1(n_4200),
.A2(n_433),
.A3(n_431),
.B(n_432),
.Y(n_4476)
);

AOI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_4200),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4202),
.B(n_434),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4300),
.B(n_435),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_4306),
.B(n_4285),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_SL g4481 ( 
.A(n_4229),
.B(n_435),
.Y(n_4481)
);

AND2x2_ASAP7_75t_L g4482 ( 
.A(n_4286),
.B(n_436),
.Y(n_4482)
);

INVx2_ASAP7_75t_SL g4483 ( 
.A(n_4313),
.Y(n_4483)
);

INVx3_ASAP7_75t_L g4484 ( 
.A(n_4325),
.Y(n_4484)
);

BUFx2_ASAP7_75t_R g4485 ( 
.A(n_4377),
.Y(n_4485)
);

O2A1O1Ixp33_ASAP7_75t_L g4486 ( 
.A1(n_4481),
.A2(n_4308),
.B(n_4314),
.C(n_4202),
.Y(n_4486)
);

O2A1O1Ixp33_ASAP7_75t_SL g4487 ( 
.A1(n_4481),
.A2(n_4275),
.B(n_4304),
.C(n_4259),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4441),
.B(n_4344),
.Y(n_4488)
);

A2O1A1Ixp33_ASAP7_75t_L g4489 ( 
.A1(n_4477),
.A2(n_4194),
.B(n_4229),
.C(n_4337),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4389),
.B(n_4292),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4425),
.B(n_4230),
.Y(n_4491)
);

O2A1O1Ixp33_ASAP7_75t_SL g4492 ( 
.A1(n_4348),
.A2(n_4304),
.B(n_4247),
.C(n_4315),
.Y(n_4492)
);

OR2x6_ASAP7_75t_L g4493 ( 
.A(n_4379),
.B(n_4325),
.Y(n_4493)
);

O2A1O1Ixp33_ASAP7_75t_L g4494 ( 
.A1(n_4339),
.A2(n_4314),
.B(n_4194),
.C(n_4319),
.Y(n_4494)
);

AOI221xp5_ASAP7_75t_L g4495 ( 
.A1(n_4425),
.A2(n_4230),
.B1(n_4271),
.B2(n_4216),
.C(n_4326),
.Y(n_4495)
);

INVx1_ASAP7_75t_SL g4496 ( 
.A(n_4377),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4401),
.B(n_4292),
.Y(n_4497)
);

INVx1_ASAP7_75t_SL g4498 ( 
.A(n_4366),
.Y(n_4498)
);

AOI221xp5_ASAP7_75t_L g4499 ( 
.A1(n_4356),
.A2(n_4271),
.B1(n_4216),
.B2(n_4326),
.C(n_4319),
.Y(n_4499)
);

INVx3_ASAP7_75t_L g4500 ( 
.A(n_4411),
.Y(n_4500)
);

AOI22xp5_ASAP7_75t_L g4501 ( 
.A1(n_4346),
.A2(n_4454),
.B1(n_4472),
.B2(n_4427),
.Y(n_4501)
);

OR2x6_ASAP7_75t_L g4502 ( 
.A(n_4388),
.B(n_4325),
.Y(n_4502)
);

NOR2xp33_ASAP7_75t_L g4503 ( 
.A(n_4411),
.B(n_4278),
.Y(n_4503)
);

OR2x2_ASAP7_75t_L g4504 ( 
.A(n_4458),
.B(n_4274),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4484),
.B(n_4274),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4343),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4484),
.B(n_4274),
.Y(n_4507)
);

NOR2xp33_ASAP7_75t_L g4508 ( 
.A(n_4366),
.B(n_4253),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4378),
.B(n_4357),
.Y(n_4509)
);

CKINVDCx5p33_ASAP7_75t_R g4510 ( 
.A(n_4366),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4413),
.Y(n_4511)
);

CKINVDCx5p33_ASAP7_75t_R g4512 ( 
.A(n_4413),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4352),
.B(n_4291),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4343),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4352),
.B(n_4293),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_4454),
.A2(n_4311),
.B1(n_4305),
.B2(n_4294),
.Y(n_4516)
);

OR2x2_ASAP7_75t_L g4517 ( 
.A(n_4414),
.B(n_4412),
.Y(n_4517)
);

OA21x2_ASAP7_75t_L g4518 ( 
.A1(n_4341),
.A2(n_4335),
.B(n_4298),
.Y(n_4518)
);

AND2x2_ASAP7_75t_L g4519 ( 
.A(n_4352),
.B(n_4297),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4380),
.B(n_4267),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4349),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4361),
.B(n_4301),
.Y(n_4522)
);

AO32x1_ASAP7_75t_L g4523 ( 
.A1(n_4483),
.A2(n_4323),
.A3(n_4279),
.B1(n_4309),
.B2(n_4321),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_4374),
.B(n_4358),
.Y(n_4524)
);

AOI21xp5_ASAP7_75t_SL g4525 ( 
.A1(n_4427),
.A2(n_4318),
.B(n_4334),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4444),
.B(n_4272),
.Y(n_4526)
);

AND2x2_ASAP7_75t_L g4527 ( 
.A(n_4444),
.B(n_4260),
.Y(n_4527)
);

NOR2x1_ASAP7_75t_SL g4528 ( 
.A(n_4471),
.B(n_4303),
.Y(n_4528)
);

NAND3xp33_ASAP7_75t_L g4529 ( 
.A(n_4456),
.B(n_4242),
.C(n_4334),
.Y(n_4529)
);

OA21x2_ASAP7_75t_L g4530 ( 
.A1(n_4442),
.A2(n_4429),
.B(n_4428),
.Y(n_4530)
);

OAI221xp5_ASAP7_75t_SL g4531 ( 
.A1(n_4376),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.C(n_440),
.Y(n_4531)
);

OAI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_4372),
.A2(n_438),
.B(n_441),
.Y(n_4532)
);

AOI21xp33_ASAP7_75t_L g4533 ( 
.A1(n_4346),
.A2(n_441),
.B(n_442),
.Y(n_4533)
);

INVxp67_ASAP7_75t_L g4534 ( 
.A(n_4406),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4460),
.B(n_442),
.Y(n_4535)
);

OR2x2_ASAP7_75t_L g4536 ( 
.A(n_4412),
.B(n_443),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4460),
.B(n_4360),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4449),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4360),
.B(n_443),
.Y(n_4539)
);

AND2x4_ASAP7_75t_L g4540 ( 
.A(n_4469),
.B(n_629),
.Y(n_4540)
);

OR2x2_ASAP7_75t_L g4541 ( 
.A(n_4364),
.B(n_444),
.Y(n_4541)
);

OR2x6_ASAP7_75t_L g4542 ( 
.A(n_4396),
.B(n_4369),
.Y(n_4542)
);

OAI21xp5_ASAP7_75t_L g4543 ( 
.A1(n_4372),
.A2(n_4345),
.B(n_4456),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4349),
.Y(n_4544)
);

AO32x2_ASAP7_75t_L g4545 ( 
.A1(n_4416),
.A2(n_444),
.A3(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_4545)
);

AND2x4_ASAP7_75t_L g4546 ( 
.A(n_4449),
.B(n_447),
.Y(n_4546)
);

OAI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_4427),
.A2(n_448),
.B(n_449),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4480),
.B(n_449),
.Y(n_4548)
);

INVx3_ASAP7_75t_L g4549 ( 
.A(n_4369),
.Y(n_4549)
);

NOR2x1_ASAP7_75t_SL g4550 ( 
.A(n_4397),
.B(n_450),
.Y(n_4550)
);

OR2x6_ASAP7_75t_L g4551 ( 
.A(n_4396),
.B(n_450),
.Y(n_4551)
);

OR2x2_ASAP7_75t_L g4552 ( 
.A(n_4342),
.B(n_451),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4469),
.B(n_452),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4371),
.Y(n_4554)
);

NOR2xp33_ASAP7_75t_L g4555 ( 
.A(n_4464),
.B(n_453),
.Y(n_4555)
);

INVx8_ASAP7_75t_L g4556 ( 
.A(n_4396),
.Y(n_4556)
);

INVxp67_ASAP7_75t_L g4557 ( 
.A(n_4406),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4371),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4476),
.B(n_454),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4398),
.Y(n_4560)
);

INVx2_ASAP7_75t_SL g4561 ( 
.A(n_4369),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4474),
.B(n_454),
.Y(n_4562)
);

AOI22xp5_ASAP7_75t_L g4563 ( 
.A1(n_4472),
.A2(n_455),
.B1(n_456),
.B2(n_457),
.Y(n_4563)
);

AND2x2_ASAP7_75t_SL g4564 ( 
.A(n_4472),
.B(n_4351),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4478),
.A2(n_457),
.B(n_458),
.Y(n_4565)
);

AO32x2_ASAP7_75t_L g4566 ( 
.A1(n_4383),
.A2(n_459),
.A3(n_460),
.B1(n_461),
.B2(n_462),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4476),
.B(n_460),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4474),
.B(n_461),
.Y(n_4568)
);

AOI22xp5_ASAP7_75t_L g4569 ( 
.A1(n_4402),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4398),
.Y(n_4570)
);

OR2x2_ASAP7_75t_L g4571 ( 
.A(n_4351),
.B(n_463),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4375),
.Y(n_4572)
);

OR2x2_ASAP7_75t_L g4573 ( 
.A(n_4351),
.B(n_465),
.Y(n_4573)
);

BUFx2_ASAP7_75t_L g4574 ( 
.A(n_4464),
.Y(n_4574)
);

OR2x2_ASAP7_75t_L g4575 ( 
.A(n_4475),
.B(n_466),
.Y(n_4575)
);

NAND2xp33_ASAP7_75t_L g4576 ( 
.A(n_4407),
.B(n_4369),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4465),
.B(n_466),
.Y(n_4577)
);

O2A1O1Ixp33_ASAP7_75t_SL g4578 ( 
.A1(n_4442),
.A2(n_467),
.B(n_468),
.C(n_469),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4375),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4376),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.Y(n_4580)
);

OR2x2_ASAP7_75t_L g4581 ( 
.A(n_4418),
.B(n_470),
.Y(n_4581)
);

OR2x2_ASAP7_75t_L g4582 ( 
.A(n_4419),
.B(n_4430),
.Y(n_4582)
);

OR2x2_ASAP7_75t_L g4583 ( 
.A(n_4383),
.B(n_472),
.Y(n_4583)
);

NOR2xp33_ASAP7_75t_L g4584 ( 
.A(n_4452),
.B(n_474),
.Y(n_4584)
);

INVx3_ASAP7_75t_L g4585 ( 
.A(n_4452),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4465),
.B(n_474),
.Y(n_4586)
);

NOR2x1_ASAP7_75t_SL g4587 ( 
.A(n_4399),
.B(n_475),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4381),
.Y(n_4588)
);

O2A1O1Ixp33_ASAP7_75t_SL g4589 ( 
.A1(n_4435),
.A2(n_475),
.B(n_476),
.C(n_477),
.Y(n_4589)
);

A2O1A1Ixp33_ASAP7_75t_L g4590 ( 
.A1(n_4435),
.A2(n_476),
.B(n_477),
.C(n_478),
.Y(n_4590)
);

OR2x2_ASAP7_75t_L g4591 ( 
.A(n_4400),
.B(n_478),
.Y(n_4591)
);

OAI21x1_ASAP7_75t_L g4592 ( 
.A1(n_4395),
.A2(n_479),
.B(n_480),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4381),
.Y(n_4593)
);

OAI22xp5_ASAP7_75t_L g4594 ( 
.A1(n_4363),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_4594)
);

OR2x6_ASAP7_75t_L g4595 ( 
.A(n_4452),
.B(n_481),
.Y(n_4595)
);

AOI221xp5_ASAP7_75t_L g4596 ( 
.A1(n_4433),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.C(n_485),
.Y(n_4596)
);

A2O1A1Ixp33_ASAP7_75t_L g4597 ( 
.A1(n_4455),
.A2(n_482),
.B(n_483),
.C(n_484),
.Y(n_4597)
);

OAI22xp5_ASAP7_75t_L g4598 ( 
.A1(n_4363),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_4598)
);

OR2x2_ASAP7_75t_L g4599 ( 
.A(n_4400),
.B(n_486),
.Y(n_4599)
);

AND2x4_ASAP7_75t_SL g4600 ( 
.A(n_4452),
.B(n_487),
.Y(n_4600)
);

NOR2x1_ASAP7_75t_SL g4601 ( 
.A(n_4399),
.B(n_488),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4453),
.Y(n_4602)
);

AND2x4_ASAP7_75t_L g4603 ( 
.A(n_4467),
.B(n_489),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4384),
.B(n_491),
.Y(n_4604)
);

INVxp67_ASAP7_75t_L g4605 ( 
.A(n_4417),
.Y(n_4605)
);

CKINVDCx12_ASAP7_75t_R g4606 ( 
.A(n_4440),
.Y(n_4606)
);

OAI21xp5_ASAP7_75t_L g4607 ( 
.A1(n_4363),
.A2(n_492),
.B(n_494),
.Y(n_4607)
);

OR2x2_ASAP7_75t_L g4608 ( 
.A(n_4445),
.B(n_495),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4382),
.Y(n_4609)
);

BUFx3_ASAP7_75t_L g4610 ( 
.A(n_4453),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4453),
.Y(n_4611)
);

OR2x2_ASAP7_75t_L g4612 ( 
.A(n_4445),
.B(n_495),
.Y(n_4612)
);

OAI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4402),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4476),
.B(n_496),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4459),
.B(n_500),
.Y(n_4615)
);

AOI21x1_ASAP7_75t_L g4616 ( 
.A1(n_4455),
.A2(n_500),
.B(n_501),
.Y(n_4616)
);

OR2x2_ASAP7_75t_L g4617 ( 
.A(n_4446),
.B(n_501),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4382),
.Y(n_4618)
);

OR2x2_ASAP7_75t_L g4619 ( 
.A(n_4447),
.B(n_502),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4453),
.Y(n_4620)
);

AOI22xp33_ASAP7_75t_L g4621 ( 
.A1(n_4491),
.A2(n_4359),
.B1(n_4404),
.B2(n_4459),
.Y(n_4621)
);

INVx2_ASAP7_75t_SL g4622 ( 
.A(n_4556),
.Y(n_4622)
);

BUFx6f_ASAP7_75t_L g4623 ( 
.A(n_4566),
.Y(n_4623)
);

AND2x2_ASAP7_75t_L g4624 ( 
.A(n_4488),
.B(n_4395),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4506),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4574),
.Y(n_4626)
);

AND2x2_ASAP7_75t_L g4627 ( 
.A(n_4493),
.B(n_4434),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4493),
.B(n_4502),
.Y(n_4628)
);

AND2x2_ASAP7_75t_L g4629 ( 
.A(n_4502),
.B(n_4434),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4524),
.B(n_4490),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4497),
.B(n_4513),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4515),
.B(n_4467),
.Y(n_4632)
);

NOR2xp33_ASAP7_75t_L g4633 ( 
.A(n_4485),
.B(n_4457),
.Y(n_4633)
);

INVx3_ASAP7_75t_L g4634 ( 
.A(n_4556),
.Y(n_4634)
);

HB1xp67_ASAP7_75t_L g4635 ( 
.A(n_4606),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4519),
.B(n_4432),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4509),
.B(n_4437),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4514),
.Y(n_4638)
);

BUFx2_ASAP7_75t_L g4639 ( 
.A(n_4542),
.Y(n_4639)
);

INVx1_ASAP7_75t_SL g4640 ( 
.A(n_4498),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4542),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4521),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4500),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4537),
.B(n_4463),
.Y(n_4644)
);

HB1xp67_ASAP7_75t_L g4645 ( 
.A(n_4534),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4505),
.B(n_4470),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4507),
.B(n_4473),
.Y(n_4647)
);

AND2x4_ASAP7_75t_L g4648 ( 
.A(n_4610),
.B(n_4462),
.Y(n_4648)
);

INVxp67_ASAP7_75t_L g4649 ( 
.A(n_4528),
.Y(n_4649)
);

BUFx3_ASAP7_75t_L g4650 ( 
.A(n_4510),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4549),
.B(n_4431),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_L g4652 ( 
.A(n_4495),
.B(n_4476),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_4550),
.B(n_4417),
.Y(n_4653)
);

HB1xp67_ASAP7_75t_L g4654 ( 
.A(n_4557),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4530),
.Y(n_4655)
);

INVxp67_ASAP7_75t_SL g4656 ( 
.A(n_4587),
.Y(n_4656)
);

HB1xp67_ASAP7_75t_L g4657 ( 
.A(n_4530),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4544),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4585),
.B(n_4431),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4554),
.Y(n_4660)
);

HB1xp67_ASAP7_75t_L g4661 ( 
.A(n_4518),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4577),
.B(n_4448),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4496),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4561),
.Y(n_4664)
);

HB1xp67_ASAP7_75t_L g4665 ( 
.A(n_4518),
.Y(n_4665)
);

HB1xp67_ASAP7_75t_L g4666 ( 
.A(n_4558),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4564),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4572),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4511),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4538),
.B(n_4436),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4603),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4586),
.B(n_4489),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4579),
.Y(n_4673)
);

INVx2_ASAP7_75t_R g4674 ( 
.A(n_4560),
.Y(n_4674)
);

INVxp67_ASAP7_75t_SL g4675 ( 
.A(n_4601),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4588),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4593),
.Y(n_4677)
);

BUFx4f_ASAP7_75t_SL g4678 ( 
.A(n_4546),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4609),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4570),
.Y(n_4680)
);

AOI221xp5_ASAP7_75t_L g4681 ( 
.A1(n_4533),
.A2(n_4462),
.B1(n_4433),
.B2(n_4423),
.C(n_4426),
.Y(n_4681)
);

OR2x6_ASAP7_75t_L g4682 ( 
.A(n_4525),
.B(n_4424),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4602),
.B(n_4436),
.Y(n_4683)
);

INVx2_ASAP7_75t_L g4684 ( 
.A(n_4603),
.Y(n_4684)
);

INVx1_ASAP7_75t_SL g4685 ( 
.A(n_4600),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4520),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4527),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4611),
.Y(n_4688)
);

AND2x2_ASAP7_75t_L g4689 ( 
.A(n_4620),
.B(n_4522),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4608),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4618),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4517),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4582),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4591),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4526),
.B(n_4404),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4599),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4543),
.B(n_4423),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4612),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4536),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4516),
.B(n_4426),
.Y(n_4700)
);

NOR2x1p5_ASAP7_75t_L g4701 ( 
.A(n_4541),
.B(n_4451),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4566),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4566),
.Y(n_4703)
);

INVx2_ASAP7_75t_L g4704 ( 
.A(n_4540),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4616),
.Y(n_4705)
);

OR2x2_ASAP7_75t_L g4706 ( 
.A(n_4571),
.B(n_4402),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4575),
.Y(n_4707)
);

AND2x2_ASAP7_75t_L g4708 ( 
.A(n_4532),
.B(n_4370),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4501),
.B(n_4370),
.Y(n_4709)
);

AND2x2_ASAP7_75t_L g4710 ( 
.A(n_4504),
.B(n_4350),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4617),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4607),
.B(n_4350),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4512),
.B(n_4353),
.Y(n_4713)
);

AND2x4_ASAP7_75t_L g4714 ( 
.A(n_4529),
.B(n_4385),
.Y(n_4714)
);

AND2x4_ASAP7_75t_L g4715 ( 
.A(n_4605),
.B(n_4385),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4576),
.B(n_4353),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4583),
.Y(n_4717)
);

INVx2_ASAP7_75t_L g4718 ( 
.A(n_4540),
.Y(n_4718)
);

AOI221xp5_ASAP7_75t_L g4719 ( 
.A1(n_4494),
.A2(n_4450),
.B1(n_4443),
.B2(n_4409),
.C(n_4405),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4615),
.B(n_4355),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4619),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_4551),
.Y(n_4722)
);

NOR2x1_ASAP7_75t_SL g4723 ( 
.A(n_4595),
.B(n_4461),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4551),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4499),
.B(n_4408),
.Y(n_4725)
);

BUFx6f_ASAP7_75t_L g4726 ( 
.A(n_4545),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4640),
.B(n_4552),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4656),
.B(n_4565),
.Y(n_4728)
);

OA21x2_ASAP7_75t_L g4729 ( 
.A1(n_4657),
.A2(n_4573),
.B(n_4547),
.Y(n_4729)
);

OAI221xp5_ASAP7_75t_SL g4730 ( 
.A1(n_4652),
.A2(n_4486),
.B1(n_4596),
.B2(n_4569),
.C(n_4563),
.Y(n_4730)
);

AOI221xp5_ASAP7_75t_L g4731 ( 
.A1(n_4725),
.A2(n_4487),
.B1(n_4492),
.B2(n_4580),
.C(n_4531),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4675),
.B(n_4539),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4702),
.B(n_4594),
.Y(n_4733)
);

NAND3xp33_ASAP7_75t_L g4734 ( 
.A(n_4623),
.B(n_4598),
.C(n_4597),
.Y(n_4734)
);

AOI211xp5_ASAP7_75t_L g4735 ( 
.A1(n_4681),
.A2(n_4589),
.B(n_4578),
.C(n_4590),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4702),
.B(n_4584),
.Y(n_4736)
);

OAI22xp33_ASAP7_75t_L g4737 ( 
.A1(n_4726),
.A2(n_4614),
.B1(n_4559),
.B2(n_4567),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4703),
.B(n_4535),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4645),
.Y(n_4739)
);

NAND3xp33_ASAP7_75t_L g4740 ( 
.A(n_4623),
.B(n_4613),
.C(n_4408),
.Y(n_4740)
);

OAI21xp5_ASAP7_75t_SL g4741 ( 
.A1(n_4672),
.A2(n_4508),
.B(n_4503),
.Y(n_4741)
);

NAND3xp33_ASAP7_75t_L g4742 ( 
.A(n_4623),
.B(n_4408),
.C(n_4595),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4631),
.B(n_4548),
.Y(n_4743)
);

NAND3xp33_ASAP7_75t_L g4744 ( 
.A(n_4623),
.B(n_4359),
.C(n_4555),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4703),
.B(n_4581),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4626),
.B(n_4553),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4654),
.Y(n_4747)
);

AOI22xp33_ASAP7_75t_SL g4748 ( 
.A1(n_4726),
.A2(n_4359),
.B1(n_4523),
.B2(n_4424),
.Y(n_4748)
);

NAND3xp33_ASAP7_75t_L g4749 ( 
.A(n_4623),
.B(n_4604),
.C(n_4420),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4626),
.B(n_4562),
.Y(n_4750)
);

OAI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_4667),
.A2(n_4592),
.B(n_4424),
.Y(n_4751)
);

AOI21xp33_ASAP7_75t_SL g4752 ( 
.A1(n_4682),
.A2(n_4468),
.B(n_4466),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4631),
.B(n_4568),
.Y(n_4753)
);

AOI21xp5_ASAP7_75t_L g4754 ( 
.A1(n_4723),
.A2(n_4523),
.B(n_4468),
.Y(n_4754)
);

NOR3xp33_ASAP7_75t_SL g4755 ( 
.A(n_4633),
.B(n_4403),
.C(n_4410),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4726),
.B(n_4466),
.Y(n_4756)
);

AOI22xp5_ASAP7_75t_L g4757 ( 
.A1(n_4726),
.A2(n_4466),
.B1(n_4468),
.B2(n_4340),
.Y(n_4757)
);

AND2x2_ASAP7_75t_L g4758 ( 
.A(n_4630),
.B(n_4438),
.Y(n_4758)
);

OAI221xp5_ASAP7_75t_L g4759 ( 
.A1(n_4719),
.A2(n_4682),
.B1(n_4621),
.B2(n_4649),
.C(n_4726),
.Y(n_4759)
);

AOI22xp33_ASAP7_75t_SL g4760 ( 
.A1(n_4723),
.A2(n_4390),
.B1(n_4482),
.B2(n_4479),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4630),
.B(n_4354),
.Y(n_4761)
);

OAI22xp5_ASAP7_75t_L g4762 ( 
.A1(n_4682),
.A2(n_4545),
.B1(n_4362),
.B2(n_4365),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4722),
.B(n_4367),
.Y(n_4763)
);

NAND3xp33_ASAP7_75t_L g4764 ( 
.A(n_4661),
.B(n_4421),
.C(n_4394),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4722),
.B(n_4368),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4724),
.B(n_4373),
.Y(n_4766)
);

NAND3xp33_ASAP7_75t_L g4767 ( 
.A(n_4665),
.B(n_4697),
.C(n_4667),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4724),
.B(n_4391),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4686),
.B(n_4422),
.Y(n_4769)
);

OAI22xp5_ASAP7_75t_L g4770 ( 
.A1(n_4682),
.A2(n_4653),
.B1(n_4706),
.B2(n_4705),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4686),
.B(n_4663),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4663),
.B(n_4422),
.Y(n_4772)
);

AND2x2_ASAP7_75t_L g4773 ( 
.A(n_4628),
.B(n_4355),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4671),
.B(n_4386),
.Y(n_4774)
);

NOR2xp33_ASAP7_75t_L g4775 ( 
.A(n_4678),
.B(n_4650),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_4628),
.B(n_4386),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4715),
.Y(n_4777)
);

AND2x2_ASAP7_75t_L g4778 ( 
.A(n_4624),
.B(n_4387),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4624),
.B(n_4387),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_L g4780 ( 
.A(n_4671),
.B(n_4684),
.Y(n_4780)
);

OAI221xp5_ASAP7_75t_L g4781 ( 
.A1(n_4622),
.A2(n_4439),
.B1(n_4393),
.B2(n_4392),
.C(n_4415),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4684),
.B(n_4392),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4635),
.B(n_4393),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4650),
.B(n_4634),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4705),
.B(n_4415),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_SL g4786 ( 
.A(n_4634),
.B(n_4347),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4717),
.B(n_4347),
.Y(n_4787)
);

OAI22xp5_ASAP7_75t_SL g4788 ( 
.A1(n_4685),
.A2(n_4622),
.B1(n_4706),
.B2(n_4634),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4704),
.B(n_4439),
.Y(n_4789)
);

AND2x2_ASAP7_75t_L g4790 ( 
.A(n_4627),
.B(n_4545),
.Y(n_4790)
);

OR2x2_ASAP7_75t_L g4791 ( 
.A(n_4756),
.B(n_4717),
.Y(n_4791)
);

AND2x4_ASAP7_75t_L g4792 ( 
.A(n_4784),
.B(n_4643),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4780),
.Y(n_4793)
);

OR2x2_ASAP7_75t_L g4794 ( 
.A(n_4738),
.B(n_4669),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4777),
.Y(n_4795)
);

AND2x2_ASAP7_75t_L g4796 ( 
.A(n_4753),
.B(n_4627),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4735),
.B(n_4666),
.Y(n_4797)
);

AND2x2_ASAP7_75t_L g4798 ( 
.A(n_4758),
.B(n_4689),
.Y(n_4798)
);

INVxp67_ASAP7_75t_SL g4799 ( 
.A(n_4788),
.Y(n_4799)
);

INVx4_ASAP7_75t_L g4800 ( 
.A(n_4783),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4743),
.B(n_4689),
.Y(n_4801)
);

AOI221xp5_ASAP7_75t_L g4802 ( 
.A1(n_4759),
.A2(n_4697),
.B1(n_4709),
.B2(n_4700),
.C(n_4639),
.Y(n_4802)
);

OR2x2_ASAP7_75t_L g4803 ( 
.A(n_4727),
.B(n_4669),
.Y(n_4803)
);

AND2x2_ASAP7_75t_L g4804 ( 
.A(n_4775),
.B(n_4636),
.Y(n_4804)
);

AND2x4_ASAP7_75t_L g4805 ( 
.A(n_4773),
.B(n_4643),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4760),
.B(n_4636),
.Y(n_4806)
);

AO21x2_ASAP7_75t_L g4807 ( 
.A1(n_4767),
.A2(n_4655),
.B(n_4709),
.Y(n_4807)
);

NAND3xp33_ASAP7_75t_L g4808 ( 
.A(n_4744),
.B(n_4655),
.C(n_4639),
.Y(n_4808)
);

AND2x2_ASAP7_75t_L g4809 ( 
.A(n_4790),
.B(n_4632),
.Y(n_4809)
);

INVx2_ASAP7_75t_SL g4810 ( 
.A(n_4778),
.Y(n_4810)
);

BUFx2_ASAP7_75t_L g4811 ( 
.A(n_4751),
.Y(n_4811)
);

AND2x2_ASAP7_75t_L g4812 ( 
.A(n_4761),
.B(n_4632),
.Y(n_4812)
);

INVx2_ASAP7_75t_SL g4813 ( 
.A(n_4779),
.Y(n_4813)
);

OAI22xp5_ASAP7_75t_SL g4814 ( 
.A1(n_4734),
.A2(n_4641),
.B1(n_4714),
.B2(n_4718),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4771),
.Y(n_4815)
);

NAND5xp2_ASAP7_75t_L g4816 ( 
.A(n_4741),
.B(n_4731),
.C(n_4730),
.D(n_4755),
.E(n_4747),
.Y(n_4816)
);

OAI33xp33_ASAP7_75t_L g4817 ( 
.A1(n_4737),
.A2(n_4642),
.A3(n_4658),
.B1(n_4660),
.B2(n_4680),
.B3(n_4638),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4776),
.B(n_4637),
.Y(n_4818)
);

OR2x2_ASAP7_75t_L g4819 ( 
.A(n_4736),
.B(n_4704),
.Y(n_4819)
);

AND2x2_ASAP7_75t_L g4820 ( 
.A(n_4757),
.B(n_4637),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4739),
.Y(n_4821)
);

AND2x2_ASAP7_75t_L g4822 ( 
.A(n_4751),
.B(n_4713),
.Y(n_4822)
);

INVx4_ASAP7_75t_L g4823 ( 
.A(n_4729),
.Y(n_4823)
);

BUFx2_ASAP7_75t_L g4824 ( 
.A(n_4732),
.Y(n_4824)
);

OR2x2_ASAP7_75t_L g4825 ( 
.A(n_4745),
.B(n_4718),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4729),
.B(n_4699),
.Y(n_4826)
);

OR2x2_ASAP7_75t_L g4827 ( 
.A(n_4749),
.B(n_4690),
.Y(n_4827)
);

AND2x2_ASAP7_75t_L g4828 ( 
.A(n_4752),
.B(n_4713),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4785),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4785),
.Y(n_4830)
);

CKINVDCx5p33_ASAP7_75t_R g4831 ( 
.A(n_4770),
.Y(n_4831)
);

AND2x2_ASAP7_75t_L g4832 ( 
.A(n_4746),
.B(n_4629),
.Y(n_4832)
);

HB1xp67_ASAP7_75t_L g4833 ( 
.A(n_4770),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4774),
.Y(n_4834)
);

OR2x2_ASAP7_75t_L g4835 ( 
.A(n_4750),
.B(n_4690),
.Y(n_4835)
);

NOR2x1_ASAP7_75t_SL g4836 ( 
.A(n_4742),
.B(n_4629),
.Y(n_4836)
);

INVx1_ASAP7_75t_SL g4837 ( 
.A(n_4786),
.Y(n_4837)
);

BUFx2_ASAP7_75t_L g4838 ( 
.A(n_4787),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4782),
.Y(n_4839)
);

OR2x2_ASAP7_75t_L g4840 ( 
.A(n_4733),
.B(n_4687),
.Y(n_4840)
);

OAI33xp33_ASAP7_75t_L g4841 ( 
.A1(n_4762),
.A2(n_4680),
.A3(n_4660),
.B1(n_4642),
.B2(n_4658),
.B3(n_4625),
.Y(n_4841)
);

OAI321xp33_ASAP7_75t_L g4842 ( 
.A1(n_4740),
.A2(n_4700),
.A3(n_4641),
.B1(n_4674),
.B2(n_4712),
.C(n_4716),
.Y(n_4842)
);

BUFx6f_ASAP7_75t_L g4843 ( 
.A(n_4787),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4772),
.Y(n_4844)
);

O2A1O1Ixp5_ASAP7_75t_L g4845 ( 
.A1(n_4762),
.A2(n_4714),
.B(n_4648),
.C(n_4687),
.Y(n_4845)
);

INVx1_ASAP7_75t_SL g4846 ( 
.A(n_4728),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_4748),
.B(n_4692),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4754),
.B(n_4646),
.Y(n_4848)
);

INVx2_ASAP7_75t_L g4849 ( 
.A(n_4823),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4809),
.B(n_4664),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4823),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4801),
.B(n_4664),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4848),
.B(n_4701),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4828),
.B(n_4646),
.Y(n_4854)
);

HB1xp67_ASAP7_75t_L g4855 ( 
.A(n_4807),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4796),
.B(n_4647),
.Y(n_4856)
);

NOR2xp33_ASAP7_75t_L g4857 ( 
.A(n_4800),
.B(n_4707),
.Y(n_4857)
);

AND2x2_ASAP7_75t_L g4858 ( 
.A(n_4798),
.B(n_4818),
.Y(n_4858)
);

AND2x4_ASAP7_75t_L g4859 ( 
.A(n_4807),
.B(n_4648),
.Y(n_4859)
);

OR2x2_ASAP7_75t_L g4860 ( 
.A(n_4827),
.B(n_4763),
.Y(n_4860)
);

AND2x4_ASAP7_75t_L g4861 ( 
.A(n_4792),
.B(n_4648),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_4845),
.Y(n_4862)
);

OR2x2_ASAP7_75t_L g4863 ( 
.A(n_4825),
.B(n_4819),
.Y(n_4863)
);

AND2x2_ASAP7_75t_L g4864 ( 
.A(n_4804),
.B(n_4647),
.Y(n_4864)
);

AND2x4_ASAP7_75t_SL g4865 ( 
.A(n_4792),
.B(n_4694),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_4812),
.B(n_4720),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4803),
.Y(n_4867)
);

AND2x4_ASAP7_75t_L g4868 ( 
.A(n_4800),
.B(n_4688),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4791),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4794),
.Y(n_4870)
);

AND2x2_ASAP7_75t_L g4871 ( 
.A(n_4822),
.B(n_4716),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4843),
.Y(n_4872)
);

INVx3_ASAP7_75t_L g4873 ( 
.A(n_4805),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4836),
.Y(n_4874)
);

NAND3xp33_ASAP7_75t_L g4875 ( 
.A(n_4808),
.B(n_4764),
.C(n_4688),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4805),
.B(n_4806),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4843),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4837),
.B(n_4696),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4837),
.B(n_4698),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4843),
.Y(n_4880)
);

INVxp67_ASAP7_75t_L g4881 ( 
.A(n_4833),
.Y(n_4881)
);

AND2x4_ASAP7_75t_L g4882 ( 
.A(n_4808),
.B(n_4715),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4835),
.Y(n_4883)
);

OAI21xp33_ASAP7_75t_SL g4884 ( 
.A1(n_4799),
.A2(n_4674),
.B(n_4712),
.Y(n_4884)
);

OR2x2_ASAP7_75t_L g4885 ( 
.A(n_4840),
.B(n_4765),
.Y(n_4885)
);

AND2x2_ASAP7_75t_L g4886 ( 
.A(n_4820),
.B(n_4720),
.Y(n_4886)
);

INVx2_ASAP7_75t_L g4887 ( 
.A(n_4811),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_4826),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4802),
.B(n_4711),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_L g4890 ( 
.A(n_4832),
.B(n_4721),
.Y(n_4890)
);

AND2x2_ASAP7_75t_L g4891 ( 
.A(n_4824),
.B(n_4644),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4810),
.B(n_4693),
.Y(n_4892)
);

OR2x2_ASAP7_75t_L g4893 ( 
.A(n_4797),
.B(n_4766),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4861),
.B(n_4813),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4861),
.B(n_4856),
.Y(n_4895)
);

AND2x2_ASAP7_75t_L g4896 ( 
.A(n_4854),
.B(n_4846),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4871),
.B(n_4846),
.Y(n_4897)
);

AOI22xp5_ASAP7_75t_L g4898 ( 
.A1(n_4862),
.A2(n_4814),
.B1(n_4797),
.B2(n_4831),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4861),
.B(n_4795),
.Y(n_4899)
);

AND2x2_ASAP7_75t_L g4900 ( 
.A(n_4871),
.B(n_4838),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4855),
.Y(n_4901)
);

INVx2_ASAP7_75t_L g4902 ( 
.A(n_4855),
.Y(n_4902)
);

NOR2x1_ASAP7_75t_SL g4903 ( 
.A(n_4863),
.B(n_4826),
.Y(n_4903)
);

OR2x6_ASAP7_75t_L g4904 ( 
.A(n_4849),
.B(n_4851),
.Y(n_4904)
);

NAND2xp5_ASAP7_75t_L g4905 ( 
.A(n_4873),
.B(n_4847),
.Y(n_4905)
);

INVx2_ASAP7_75t_L g4906 ( 
.A(n_4859),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4859),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4873),
.B(n_4847),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_4864),
.B(n_4821),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4859),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4849),
.Y(n_4911)
);

INVx2_ASAP7_75t_L g4912 ( 
.A(n_4851),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4865),
.Y(n_4913)
);

OR2x2_ASAP7_75t_L g4914 ( 
.A(n_4850),
.B(n_4768),
.Y(n_4914)
);

OR2x2_ASAP7_75t_L g4915 ( 
.A(n_4852),
.B(n_4887),
.Y(n_4915)
);

INVx2_ASAP7_75t_L g4916 ( 
.A(n_4882),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4874),
.B(n_4793),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4886),
.B(n_4644),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4865),
.Y(n_4919)
);

INVx3_ASAP7_75t_L g4920 ( 
.A(n_4882),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_L g4921 ( 
.A(n_4881),
.B(n_4815),
.Y(n_4921)
);

INVx2_ASAP7_75t_SL g4922 ( 
.A(n_4868),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4881),
.B(n_4814),
.Y(n_4923)
);

AND2x2_ASAP7_75t_L g4924 ( 
.A(n_4874),
.B(n_4670),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4891),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4900),
.B(n_4858),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4903),
.Y(n_4927)
);

INVx2_ASAP7_75t_L g4928 ( 
.A(n_4920),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4920),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4920),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4906),
.Y(n_4931)
);

AND2x4_ASAP7_75t_L g4932 ( 
.A(n_4922),
.B(n_4868),
.Y(n_4932)
);

XNOR2xp5_ASAP7_75t_L g4933 ( 
.A(n_4898),
.B(n_4853),
.Y(n_4933)
);

INVxp67_ASAP7_75t_SL g4934 ( 
.A(n_4906),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4907),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4910),
.Y(n_4936)
);

AOI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4918),
.A2(n_4862),
.B1(n_4884),
.B2(n_4889),
.Y(n_4937)
);

AOI22xp33_ASAP7_75t_L g4938 ( 
.A1(n_4925),
.A2(n_4816),
.B1(n_4875),
.B2(n_4882),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4896),
.B(n_4866),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4922),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4916),
.Y(n_4941)
);

AND2x4_ASAP7_75t_L g4942 ( 
.A(n_4916),
.B(n_4868),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_4900),
.B(n_4887),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4897),
.Y(n_4944)
);

OR2x2_ASAP7_75t_L g4945 ( 
.A(n_4905),
.B(n_4908),
.Y(n_4945)
);

AND2x2_ASAP7_75t_L g4946 ( 
.A(n_4909),
.B(n_4876),
.Y(n_4946)
);

NAND2x1p5_ASAP7_75t_L g4947 ( 
.A(n_4913),
.B(n_4872),
.Y(n_4947)
);

NAND3xp33_ASAP7_75t_L g4948 ( 
.A(n_4919),
.B(n_4888),
.C(n_4857),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4902),
.Y(n_4949)
);

OR2x2_ASAP7_75t_L g4950 ( 
.A(n_4926),
.B(n_4923),
.Y(n_4950)
);

INVx2_ASAP7_75t_L g4951 ( 
.A(n_4932),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4932),
.Y(n_4952)
);

INVx1_ASAP7_75t_SL g4953 ( 
.A(n_4942),
.Y(n_4953)
);

XNOR2xp5_ASAP7_75t_L g4954 ( 
.A(n_4933),
.B(n_4897),
.Y(n_4954)
);

INVx2_ASAP7_75t_SL g4955 ( 
.A(n_4942),
.Y(n_4955)
);

INVx2_ASAP7_75t_L g4956 ( 
.A(n_4928),
.Y(n_4956)
);

XOR2x2_ASAP7_75t_L g4957 ( 
.A(n_4939),
.B(n_4895),
.Y(n_4957)
);

INVx4_ASAP7_75t_L g4958 ( 
.A(n_4929),
.Y(n_4958)
);

AOI22xp5_ASAP7_75t_SL g4959 ( 
.A1(n_4927),
.A2(n_4888),
.B1(n_4816),
.B2(n_4901),
.Y(n_4959)
);

XNOR2xp5_ASAP7_75t_L g4960 ( 
.A(n_4937),
.B(n_4946),
.Y(n_4960)
);

INVx1_ASAP7_75t_SL g4961 ( 
.A(n_4927),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4930),
.Y(n_4962)
);

AND2x2_ASAP7_75t_L g4963 ( 
.A(n_4944),
.B(n_4909),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4943),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4934),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4940),
.Y(n_4966)
);

INVx2_ASAP7_75t_SL g4967 ( 
.A(n_4947),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4931),
.Y(n_4968)
);

INVx2_ASAP7_75t_SL g4969 ( 
.A(n_4941),
.Y(n_4969)
);

INVx2_ASAP7_75t_L g4970 ( 
.A(n_4949),
.Y(n_4970)
);

CKINVDCx16_ASAP7_75t_R g4971 ( 
.A(n_4954),
.Y(n_4971)
);

AND2x2_ASAP7_75t_L g4972 ( 
.A(n_4963),
.B(n_4924),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4952),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4953),
.B(n_4924),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4967),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4951),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4955),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4953),
.B(n_4883),
.Y(n_4978)
);

INVx1_ASAP7_75t_SL g4979 ( 
.A(n_4961),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4957),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4958),
.Y(n_4981)
);

AND2x2_ASAP7_75t_L g4982 ( 
.A(n_4956),
.B(n_4869),
.Y(n_4982)
);

NOR2xp33_ASAP7_75t_L g4983 ( 
.A(n_4958),
.B(n_4948),
.Y(n_4983)
);

INVx2_ASAP7_75t_SL g4984 ( 
.A(n_4965),
.Y(n_4984)
);

NOR2xp33_ASAP7_75t_L g4985 ( 
.A(n_4966),
.B(n_4894),
.Y(n_4985)
);

INVxp67_ASAP7_75t_L g4986 ( 
.A(n_4974),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4974),
.Y(n_4987)
);

OR2x2_ASAP7_75t_L g4988 ( 
.A(n_4971),
.B(n_4860),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4972),
.Y(n_4989)
);

AOI22xp33_ASAP7_75t_L g4990 ( 
.A1(n_4977),
.A2(n_4817),
.B1(n_4938),
.B2(n_4841),
.Y(n_4990)
);

OAI22xp33_ASAP7_75t_L g4991 ( 
.A1(n_4979),
.A2(n_4842),
.B1(n_4961),
.B2(n_4879),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4978),
.Y(n_4992)
);

INVx2_ASAP7_75t_L g4993 ( 
.A(n_4979),
.Y(n_4993)
);

AOI22xp5_ASAP7_75t_L g4994 ( 
.A1(n_4980),
.A2(n_4960),
.B1(n_4857),
.B2(n_4867),
.Y(n_4994)
);

NAND2x1_ASAP7_75t_L g4995 ( 
.A(n_4992),
.B(n_4904),
.Y(n_4995)
);

OR2x2_ASAP7_75t_L g4996 ( 
.A(n_4988),
.B(n_4899),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4989),
.B(n_4917),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4987),
.Y(n_4998)
);

INVx1_ASAP7_75t_SL g4999 ( 
.A(n_4993),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4994),
.Y(n_5000)
);

AOI31xp33_ASAP7_75t_L g5001 ( 
.A1(n_4986),
.A2(n_4945),
.A3(n_4983),
.B(n_4959),
.Y(n_5001)
);

AO22x2_ASAP7_75t_L g5002 ( 
.A1(n_4991),
.A2(n_4902),
.B1(n_4949),
.B2(n_4970),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4990),
.Y(n_5003)
);

A2O1A1Ixp33_ASAP7_75t_L g5004 ( 
.A1(n_4990),
.A2(n_4842),
.B(n_4959),
.C(n_4983),
.Y(n_5004)
);

NOR2xp33_ASAP7_75t_SL g5005 ( 
.A(n_4988),
.B(n_4877),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4988),
.Y(n_5006)
);

INVx1_ASAP7_75t_SL g5007 ( 
.A(n_4988),
.Y(n_5007)
);

AND3x1_ASAP7_75t_L g5008 ( 
.A(n_4990),
.B(n_4985),
.C(n_4975),
.Y(n_5008)
);

OAI22xp5_ASAP7_75t_L g5009 ( 
.A1(n_5004),
.A2(n_4893),
.B1(n_4915),
.B2(n_4880),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4995),
.Y(n_5010)
);

AND2x2_ASAP7_75t_L g5011 ( 
.A(n_4997),
.B(n_4917),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4996),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_5002),
.Y(n_5013)
);

AND2x2_ASAP7_75t_L g5014 ( 
.A(n_5007),
.B(n_4870),
.Y(n_5014)
);

NOR2x1_ASAP7_75t_L g5015 ( 
.A(n_5001),
.B(n_4970),
.Y(n_5015)
);

AND2x2_ASAP7_75t_L g5016 ( 
.A(n_4999),
.B(n_4982),
.Y(n_5016)
);

INVx2_ASAP7_75t_L g5017 ( 
.A(n_5006),
.Y(n_5017)
);

INVxp67_ASAP7_75t_SL g5018 ( 
.A(n_5005),
.Y(n_5018)
);

NAND2x1_ASAP7_75t_SL g5019 ( 
.A(n_5000),
.B(n_4912),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_5002),
.Y(n_5020)
);

NOR2xp33_ASAP7_75t_L g5021 ( 
.A(n_5003),
.B(n_4976),
.Y(n_5021)
);

AND2x2_ASAP7_75t_L g5022 ( 
.A(n_5008),
.B(n_4973),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4998),
.Y(n_5023)
);

AND2x2_ASAP7_75t_L g5024 ( 
.A(n_4997),
.B(n_4964),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4997),
.B(n_4935),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4995),
.Y(n_5026)
);

AND2x2_ASAP7_75t_L g5027 ( 
.A(n_4997),
.B(n_4936),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4995),
.Y(n_5028)
);

AND2x2_ASAP7_75t_L g5029 ( 
.A(n_4997),
.B(n_4969),
.Y(n_5029)
);

OAI22xp5_ASAP7_75t_L g5030 ( 
.A1(n_5004),
.A2(n_4878),
.B1(n_4885),
.B2(n_4890),
.Y(n_5030)
);

NOR2xp33_ASAP7_75t_L g5031 ( 
.A(n_4995),
.B(n_4914),
.Y(n_5031)
);

AOI221xp5_ASAP7_75t_L g5032 ( 
.A1(n_5009),
.A2(n_4911),
.B1(n_4962),
.B2(n_4968),
.C(n_4912),
.Y(n_5032)
);

NAND4xp25_ASAP7_75t_SL g5033 ( 
.A(n_5010),
.B(n_4921),
.C(n_4950),
.D(n_4892),
.Y(n_5033)
);

AOI22xp5_ASAP7_75t_L g5034 ( 
.A1(n_5021),
.A2(n_4984),
.B1(n_4981),
.B2(n_4904),
.Y(n_5034)
);

AOI22xp5_ASAP7_75t_L g5035 ( 
.A1(n_5030),
.A2(n_4904),
.B1(n_4844),
.B2(n_4839),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_5011),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_5019),
.Y(n_5037)
);

OAI22xp5_ASAP7_75t_L g5038 ( 
.A1(n_5026),
.A2(n_4834),
.B1(n_4830),
.B2(n_4829),
.Y(n_5038)
);

OA22x2_ASAP7_75t_L g5039 ( 
.A1(n_5028),
.A2(n_4715),
.B1(n_4789),
.B2(n_4769),
.Y(n_5039)
);

INVx1_ASAP7_75t_L g5040 ( 
.A(n_5015),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_5015),
.Y(n_5041)
);

AOI221xp5_ASAP7_75t_L g5042 ( 
.A1(n_5009),
.A2(n_4781),
.B1(n_4677),
.B2(n_4676),
.C(n_4679),
.Y(n_5042)
);

OA22x2_ASAP7_75t_L g5043 ( 
.A1(n_5018),
.A2(n_4673),
.B1(n_4668),
.B2(n_4691),
.Y(n_5043)
);

A2O1A1Ixp33_ASAP7_75t_L g5044 ( 
.A1(n_5031),
.A2(n_4714),
.B(n_4683),
.C(n_4670),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_5027),
.Y(n_5045)
);

CKINVDCx5p33_ASAP7_75t_R g5046 ( 
.A(n_5014),
.Y(n_5046)
);

INVx2_ASAP7_75t_L g5047 ( 
.A(n_5029),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_5013),
.Y(n_5048)
);

OA22x2_ASAP7_75t_L g5049 ( 
.A1(n_5020),
.A2(n_4683),
.B1(n_4710),
.B2(n_4662),
.Y(n_5049)
);

AOI22xp5_ASAP7_75t_L g5050 ( 
.A1(n_5016),
.A2(n_4710),
.B1(n_4708),
.B2(n_4695),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_5025),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_5022),
.Y(n_5052)
);

INVx2_ASAP7_75t_SL g5053 ( 
.A(n_5024),
.Y(n_5053)
);

NAND4xp75_ASAP7_75t_SL g5054 ( 
.A(n_5017),
.B(n_4708),
.C(n_4695),
.D(n_4659),
.Y(n_5054)
);

AO22x2_ASAP7_75t_L g5055 ( 
.A1(n_5012),
.A2(n_4659),
.B1(n_4651),
.B2(n_504),
.Y(n_5055)
);

OAI22xp5_ASAP7_75t_L g5056 ( 
.A1(n_5023),
.A2(n_4651),
.B1(n_503),
.B2(n_504),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_5011),
.Y(n_5057)
);

NAND3xp33_ASAP7_75t_L g5058 ( 
.A(n_5032),
.B(n_502),
.C(n_503),
.Y(n_5058)
);

BUFx2_ASAP7_75t_L g5059 ( 
.A(n_5055),
.Y(n_5059)
);

OAI21xp5_ASAP7_75t_L g5060 ( 
.A1(n_5034),
.A2(n_505),
.B(n_507),
.Y(n_5060)
);

NOR3xp33_ASAP7_75t_L g5061 ( 
.A(n_5033),
.B(n_505),
.C(n_507),
.Y(n_5061)
);

OA22x2_ASAP7_75t_L g5062 ( 
.A1(n_5035),
.A2(n_508),
.B1(n_510),
.B2(n_511),
.Y(n_5062)
);

NOR3xp33_ASAP7_75t_L g5063 ( 
.A(n_5036),
.B(n_510),
.C(n_511),
.Y(n_5063)
);

AOI21xp5_ASAP7_75t_L g5064 ( 
.A1(n_5053),
.A2(n_512),
.B(n_513),
.Y(n_5064)
);

OA22x2_ASAP7_75t_L g5065 ( 
.A1(n_5050),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_5065)
);

AOI22xp5_ASAP7_75t_L g5066 ( 
.A1(n_5052),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_5044),
.B(n_517),
.Y(n_5067)
);

OAI21xp5_ASAP7_75t_L g5068 ( 
.A1(n_5057),
.A2(n_518),
.B(n_519),
.Y(n_5068)
);

OAI211xp5_ASAP7_75t_SL g5069 ( 
.A1(n_5045),
.A2(n_518),
.B(n_519),
.C(n_520),
.Y(n_5069)
);

OA22x2_ASAP7_75t_L g5070 ( 
.A1(n_5048),
.A2(n_521),
.B1(n_522),
.B2(n_523),
.Y(n_5070)
);

OAI21xp5_ASAP7_75t_L g5071 ( 
.A1(n_5038),
.A2(n_521),
.B(n_522),
.Y(n_5071)
);

AOI22xp5_ASAP7_75t_L g5072 ( 
.A1(n_5046),
.A2(n_523),
.B1(n_524),
.B2(n_525),
.Y(n_5072)
);

AO22x2_ASAP7_75t_L g5073 ( 
.A1(n_5040),
.A2(n_526),
.B1(n_527),
.B2(n_528),
.Y(n_5073)
);

NOR3x1_ASAP7_75t_L g5074 ( 
.A(n_5056),
.B(n_5041),
.C(n_5051),
.Y(n_5074)
);

OAI21xp33_ASAP7_75t_L g5075 ( 
.A1(n_5047),
.A2(n_528),
.B(n_529),
.Y(n_5075)
);

NOR3x1_ASAP7_75t_L g5076 ( 
.A(n_5055),
.B(n_529),
.C(n_530),
.Y(n_5076)
);

AOI211xp5_ASAP7_75t_L g5077 ( 
.A1(n_5037),
.A2(n_530),
.B(n_531),
.C(n_532),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_5042),
.B(n_531),
.Y(n_5078)
);

NOR3xp33_ASAP7_75t_L g5079 ( 
.A(n_5054),
.B(n_532),
.C(n_533),
.Y(n_5079)
);

AOI21xp5_ASAP7_75t_L g5080 ( 
.A1(n_5039),
.A2(n_5043),
.B(n_5049),
.Y(n_5080)
);

INVxp67_ASAP7_75t_L g5081 ( 
.A(n_5055),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_5079),
.B(n_533),
.Y(n_5082)
);

AOI21xp5_ASAP7_75t_L g5083 ( 
.A1(n_5081),
.A2(n_5059),
.B(n_5078),
.Y(n_5083)
);

NOR2x1_ASAP7_75t_L g5084 ( 
.A(n_5058),
.B(n_534),
.Y(n_5084)
);

XOR2x2_ASAP7_75t_L g5085 ( 
.A(n_5062),
.B(n_534),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_5065),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_SL g5087 ( 
.A(n_5077),
.B(n_535),
.Y(n_5087)
);

NOR2xp33_ASAP7_75t_L g5088 ( 
.A(n_5075),
.B(n_535),
.Y(n_5088)
);

NOR2xp67_ASAP7_75t_L g5089 ( 
.A(n_5064),
.B(n_536),
.Y(n_5089)
);

A2O1A1Ixp33_ASAP7_75t_L g5090 ( 
.A1(n_5080),
.A2(n_537),
.B(n_538),
.C(n_539),
.Y(n_5090)
);

AOI22xp5_ASAP7_75t_L g5091 ( 
.A1(n_5061),
.A2(n_537),
.B1(n_538),
.B2(n_539),
.Y(n_5091)
);

AOI211x1_ASAP7_75t_L g5092 ( 
.A1(n_5067),
.A2(n_540),
.B(n_542),
.C(n_543),
.Y(n_5092)
);

NOR2x1_ASAP7_75t_L g5093 ( 
.A(n_5060),
.B(n_540),
.Y(n_5093)
);

NAND3xp33_ASAP7_75t_L g5094 ( 
.A(n_5071),
.B(n_543),
.C(n_545),
.Y(n_5094)
);

NOR2xp33_ASAP7_75t_L g5095 ( 
.A(n_5069),
.B(n_545),
.Y(n_5095)
);

NOR2xp33_ASAP7_75t_L g5096 ( 
.A(n_5068),
.B(n_546),
.Y(n_5096)
);

INVx2_ASAP7_75t_L g5097 ( 
.A(n_5073),
.Y(n_5097)
);

NAND3xp33_ASAP7_75t_L g5098 ( 
.A(n_5063),
.B(n_546),
.C(n_548),
.Y(n_5098)
);

OAI221xp5_ASAP7_75t_L g5099 ( 
.A1(n_5090),
.A2(n_5066),
.B1(n_5072),
.B2(n_5070),
.C(n_5076),
.Y(n_5099)
);

NAND4xp75_ASAP7_75t_L g5100 ( 
.A(n_5083),
.B(n_5074),
.C(n_5073),
.D(n_554),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_5085),
.Y(n_5101)
);

NAND3xp33_ASAP7_75t_SL g5102 ( 
.A(n_5097),
.B(n_549),
.C(n_550),
.Y(n_5102)
);

NOR2x1p5_ASAP7_75t_L g5103 ( 
.A(n_5082),
.B(n_549),
.Y(n_5103)
);

NOR3xp33_ASAP7_75t_SL g5104 ( 
.A(n_5086),
.B(n_550),
.C(n_554),
.Y(n_5104)
);

NAND2xp5_ASAP7_75t_L g5105 ( 
.A(n_5092),
.B(n_556),
.Y(n_5105)
);

NOR2x1_ASAP7_75t_L g5106 ( 
.A(n_5098),
.B(n_556),
.Y(n_5106)
);

NOR2x1p5_ASAP7_75t_L g5107 ( 
.A(n_5094),
.B(n_557),
.Y(n_5107)
);

AOI211x1_ASAP7_75t_SL g5108 ( 
.A1(n_5089),
.A2(n_5087),
.B(n_5084),
.C(n_5093),
.Y(n_5108)
);

AOI21xp33_ASAP7_75t_SL g5109 ( 
.A1(n_5088),
.A2(n_558),
.B(n_559),
.Y(n_5109)
);

NAND4xp75_ASAP7_75t_L g5110 ( 
.A(n_5096),
.B(n_558),
.C(n_559),
.D(n_560),
.Y(n_5110)
);

INVxp33_ASAP7_75t_L g5111 ( 
.A(n_5095),
.Y(n_5111)
);

NOR2x1_ASAP7_75t_L g5112 ( 
.A(n_5091),
.B(n_560),
.Y(n_5112)
);

NOR3x1_ASAP7_75t_L g5113 ( 
.A(n_5098),
.B(n_561),
.C(n_562),
.Y(n_5113)
);

NOR3xp33_ASAP7_75t_SL g5114 ( 
.A(n_5100),
.B(n_628),
.C(n_563),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_5105),
.Y(n_5115)
);

OAI21xp33_ASAP7_75t_L g5116 ( 
.A1(n_5111),
.A2(n_562),
.B(n_563),
.Y(n_5116)
);

NOR3xp33_ASAP7_75t_L g5117 ( 
.A(n_5101),
.B(n_628),
.C(n_565),
.Y(n_5117)
);

OAI21xp5_ASAP7_75t_L g5118 ( 
.A1(n_5106),
.A2(n_564),
.B(n_565),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_5110),
.Y(n_5119)
);

OAI221xp5_ASAP7_75t_L g5120 ( 
.A1(n_5104),
.A2(n_5099),
.B1(n_5109),
.B2(n_5112),
.C(n_5102),
.Y(n_5120)
);

OAI221xp5_ASAP7_75t_L g5121 ( 
.A1(n_5108),
.A2(n_564),
.B1(n_566),
.B2(n_567),
.C(n_569),
.Y(n_5121)
);

AOI31xp33_ASAP7_75t_L g5122 ( 
.A1(n_5103),
.A2(n_567),
.A3(n_569),
.B(n_570),
.Y(n_5122)
);

O2A1O1Ixp33_ASAP7_75t_L g5123 ( 
.A1(n_5107),
.A2(n_571),
.B(n_572),
.C(n_573),
.Y(n_5123)
);

AOI22xp5_ASAP7_75t_L g5124 ( 
.A1(n_5113),
.A2(n_575),
.B1(n_576),
.B2(n_577),
.Y(n_5124)
);

OAI211xp5_ASAP7_75t_L g5125 ( 
.A1(n_5109),
.A2(n_575),
.B(n_577),
.C(n_578),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_5105),
.Y(n_5126)
);

AOI22xp5_ASAP7_75t_L g5127 ( 
.A1(n_5102),
.A2(n_579),
.B1(n_580),
.B2(n_581),
.Y(n_5127)
);

OAI21xp5_ASAP7_75t_L g5128 ( 
.A1(n_5100),
.A2(n_580),
.B(n_581),
.Y(n_5128)
);

NAND5xp2_ASAP7_75t_L g5129 ( 
.A(n_5099),
.B(n_582),
.C(n_583),
.D(n_584),
.E(n_586),
.Y(n_5129)
);

OAI31xp33_ASAP7_75t_L g5130 ( 
.A1(n_5099),
.A2(n_627),
.A3(n_583),
.B(n_584),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_5110),
.Y(n_5131)
);

INVx2_ASAP7_75t_L g5132 ( 
.A(n_5121),
.Y(n_5132)
);

INVx2_ASAP7_75t_L g5133 ( 
.A(n_5131),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_5115),
.Y(n_5134)
);

INVxp67_ASAP7_75t_L g5135 ( 
.A(n_5129),
.Y(n_5135)
);

OAI22xp5_ASAP7_75t_L g5136 ( 
.A1(n_5124),
.A2(n_582),
.B1(n_587),
.B2(n_588),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_5122),
.Y(n_5137)
);

BUFx4f_ASAP7_75t_SL g5138 ( 
.A(n_5126),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_5123),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_5114),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_5127),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_5125),
.Y(n_5142)
);

INVxp67_ASAP7_75t_SL g5143 ( 
.A(n_5117),
.Y(n_5143)
);

AOI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_5119),
.A2(n_587),
.B1(n_588),
.B2(n_589),
.Y(n_5144)
);

INVx2_ASAP7_75t_L g5145 ( 
.A(n_5120),
.Y(n_5145)
);

NOR2xp67_ASAP7_75t_L g5146 ( 
.A(n_5128),
.B(n_589),
.Y(n_5146)
);

AND2x2_ASAP7_75t_L g5147 ( 
.A(n_5118),
.B(n_590),
.Y(n_5147)
);

OR3x1_ASAP7_75t_L g5148 ( 
.A(n_5130),
.B(n_590),
.C(n_591),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_5148),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_5146),
.B(n_5116),
.Y(n_5150)
);

NAND2x1p5_ASAP7_75t_L g5151 ( 
.A(n_5137),
.B(n_627),
.Y(n_5151)
);

AND2x4_ASAP7_75t_L g5152 ( 
.A(n_5147),
.B(n_592),
.Y(n_5152)
);

AND2x2_ASAP7_75t_SL g5153 ( 
.A(n_5132),
.B(n_626),
.Y(n_5153)
);

XNOR2x1_ASAP7_75t_L g5154 ( 
.A(n_5145),
.B(n_5133),
.Y(n_5154)
);

NAND2x1p5_ASAP7_75t_L g5155 ( 
.A(n_5140),
.B(n_626),
.Y(n_5155)
);

NOR2xp67_ASAP7_75t_L g5156 ( 
.A(n_5144),
.B(n_5136),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_5140),
.Y(n_5157)
);

NOR3x1_ASAP7_75t_L g5158 ( 
.A(n_5143),
.B(n_593),
.C(n_594),
.Y(n_5158)
);

INVx2_ASAP7_75t_L g5159 ( 
.A(n_5134),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5153),
.Y(n_5160)
);

NOR3xp33_ASAP7_75t_L g5161 ( 
.A(n_5159),
.B(n_5142),
.C(n_5139),
.Y(n_5161)
);

HB1xp67_ASAP7_75t_L g5162 ( 
.A(n_5155),
.Y(n_5162)
);

NOR2x1_ASAP7_75t_L g5163 ( 
.A(n_5149),
.B(n_5141),
.Y(n_5163)
);

NAND4xp75_ASAP7_75t_L g5164 ( 
.A(n_5157),
.B(n_5138),
.C(n_5135),
.D(n_596),
.Y(n_5164)
);

OAI22xp33_ASAP7_75t_SL g5165 ( 
.A1(n_5150),
.A2(n_593),
.B1(n_595),
.B2(n_596),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_5164),
.Y(n_5166)
);

HB1xp67_ASAP7_75t_L g5167 ( 
.A(n_5162),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_5160),
.Y(n_5168)
);

OAI22x1_ASAP7_75t_L g5169 ( 
.A1(n_5167),
.A2(n_5152),
.B1(n_5151),
.B2(n_5163),
.Y(n_5169)
);

AOI21xp5_ASAP7_75t_L g5170 ( 
.A1(n_5168),
.A2(n_5154),
.B(n_5161),
.Y(n_5170)
);

OAI22x1_ASAP7_75t_L g5171 ( 
.A1(n_5169),
.A2(n_5166),
.B1(n_5158),
.B2(n_5170),
.Y(n_5171)
);

OAI211xp5_ASAP7_75t_L g5172 ( 
.A1(n_5171),
.A2(n_5156),
.B(n_5165),
.C(n_598),
.Y(n_5172)
);

XNOR2xp5_ASAP7_75t_L g5173 ( 
.A(n_5172),
.B(n_595),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_5173),
.Y(n_5174)
);

OAI22xp33_ASAP7_75t_L g5175 ( 
.A1(n_5174),
.A2(n_597),
.B1(n_598),
.B2(n_599),
.Y(n_5175)
);

OR3x1_ASAP7_75t_L g5176 ( 
.A(n_5175),
.B(n_597),
.C(n_599),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_5176),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_SL g5178 ( 
.A(n_5177),
.B(n_600),
.Y(n_5178)
);

AOI22xp5_ASAP7_75t_L g5179 ( 
.A1(n_5178),
.A2(n_600),
.B1(n_601),
.B2(n_602),
.Y(n_5179)
);

OAI22xp5_ASAP7_75t_L g5180 ( 
.A1(n_5179),
.A2(n_601),
.B1(n_602),
.B2(n_603),
.Y(n_5180)
);

OAI21xp5_ASAP7_75t_L g5181 ( 
.A1(n_5179),
.A2(n_603),
.B(n_604),
.Y(n_5181)
);

OAI221xp5_ASAP7_75t_R g5182 ( 
.A1(n_5181),
.A2(n_604),
.B1(n_605),
.B2(n_606),
.C(n_607),
.Y(n_5182)
);

AOI221xp5_ASAP7_75t_L g5183 ( 
.A1(n_5180),
.A2(n_605),
.B1(n_607),
.B2(n_608),
.C(n_609),
.Y(n_5183)
);

AOI22xp5_ASAP7_75t_L g5184 ( 
.A1(n_5183),
.A2(n_608),
.B1(n_611),
.B2(n_612),
.Y(n_5184)
);

AOI22xp33_ASAP7_75t_SL g5185 ( 
.A1(n_5182),
.A2(n_625),
.B1(n_612),
.B2(n_613),
.Y(n_5185)
);

AOI211xp5_ASAP7_75t_L g5186 ( 
.A1(n_5184),
.A2(n_5185),
.B(n_613),
.C(n_614),
.Y(n_5186)
);


endmodule