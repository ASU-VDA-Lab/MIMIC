module fake_jpeg_9617_n_19 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_19;

wire n_13;
wire n_14;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g12 ( 
.A(n_9),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_16),
.B(n_17),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_5),
.C(n_6),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_14),
.B(n_7),
.Y(n_19)
);


endmodule