module fake_ariane_3301_n_1493 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_372, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1493);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_372;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1493;

wire n_913;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_310),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_212),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_184),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_46),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_60),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_124),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_149),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_89),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_187),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_33),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_41),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_228),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_129),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_99),
.B(n_239),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_172),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_303),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_114),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_360),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_144),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_131),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_315),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_63),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_64),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_233),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_177),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_264),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_252),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_156),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_300),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_95),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_245),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_255),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_353),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_36),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_71),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_340),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_49),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_223),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_287),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_11),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_263),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_180),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_157),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_1),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_216),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_112),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_41),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_104),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_314),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_232),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_246),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_279),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_30),
.B(n_356),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_87),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_39),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_119),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_117),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_285),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_275),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_369),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_293),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_113),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_111),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_307),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_179),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_16),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_1),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_140),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_248),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_93),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_25),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_115),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_175),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_278),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_76),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_9),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_166),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_163),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_272),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_88),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_302),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_120),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_250),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_27),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_135),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_330),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_370),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_61),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_56),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_218),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_81),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_109),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_343),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_316),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_19),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_141),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_19),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_267),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_8),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_42),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_28),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_54),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_365),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_101),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_277),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_196),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_97),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_72),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_130),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_102),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_219),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_127),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_350),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_345),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_318),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_68),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_2),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_347),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_352),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_260),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_8),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_359),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_229),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_337),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_221),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_351),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_139),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_82),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_262),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_195),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_362),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_107),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_37),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_355),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_344),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_84),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_98),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_348),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_306),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_123),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_80),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_137),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_148),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_280),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_74),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_136),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_251),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_158),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_190),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_354),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_32),
.Y(n_531)
);

BUFx2_ASAP7_75t_SL g532 ( 
.A(n_284),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_294),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_193),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_301),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_357),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_51),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_55),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_339),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_204),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_25),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_147),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_269),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_329),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_194),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_268),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_375),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_170),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_103),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_253),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_308),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_358),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_327),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_165),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_27),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_336),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_67),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_146),
.Y(n_558)
);

BUFx5_ASAP7_75t_L g559 ( 
.A(n_282),
.Y(n_559)
);

NOR2xp67_ASAP7_75t_L g560 ( 
.A(n_21),
.B(n_341),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_266),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_40),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_59),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_349),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_182),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_438),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_433),
.B(n_564),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_438),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_531),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_489),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_468),
.A2(n_44),
.B(n_43),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_380),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_442),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_433),
.B(n_0),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_564),
.B(n_0),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_485),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_415),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_385),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_R g582 ( 
.A1(n_497),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_380),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_460),
.Y(n_584)
);

BUFx8_ASAP7_75t_SL g585 ( 
.A(n_377),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_386),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_523),
.B(n_3),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_428),
.B(n_4),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_409),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_428),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_485),
.Y(n_592)
);

BUFx8_ASAP7_75t_L g593 ( 
.A(n_466),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_420),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_382),
.B(n_5),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_432),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_489),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_468),
.A2(n_47),
.B(n_45),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_383),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_554),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_554),
.B(n_5),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_464),
.B(n_6),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_423),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_384),
.Y(n_605)
);

OA21x2_ASAP7_75t_L g606 ( 
.A1(n_387),
.A2(n_6),
.B(n_7),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_7),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_411),
.B(n_9),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_443),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_485),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_477),
.B(n_10),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

BUFx12f_ASAP7_75t_L g613 ( 
.A(n_444),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_524),
.Y(n_614)
);

OAI22x1_ASAP7_75t_L g615 ( 
.A1(n_480),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_479),
.B(n_12),
.Y(n_616)
);

OA21x2_ASAP7_75t_L g617 ( 
.A1(n_397),
.A2(n_13),
.B(n_14),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_401),
.A2(n_50),
.B(n_48),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_524),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_448),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_399),
.B(n_13),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_541),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_555),
.Y(n_624)
);

INVxp33_ASAP7_75t_SL g625 ( 
.A(n_481),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

OA21x2_ASAP7_75t_L g627 ( 
.A1(n_400),
.A2(n_14),
.B(n_15),
.Y(n_627)
);

BUFx8_ASAP7_75t_L g628 ( 
.A(n_467),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_471),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_533),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_501),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_506),
.Y(n_632)
);

BUFx12f_ASAP7_75t_L g633 ( 
.A(n_513),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_416),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_421),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_404),
.Y(n_636)
);

BUFx12f_ASAP7_75t_L g637 ( 
.A(n_376),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_526),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_529),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_447),
.B(n_15),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_424),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_476),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_425),
.B(n_16),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_426),
.B(n_17),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_427),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_507),
.B(n_52),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_516),
.B(n_17),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_419),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_429),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_445),
.Y(n_650)
);

INVx6_ASAP7_75t_L g651 ( 
.A(n_559),
.Y(n_651)
);

OA21x2_ASAP7_75t_L g652 ( 
.A1(n_437),
.A2(n_18),
.B(n_20),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_439),
.B(n_18),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_450),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_454),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_455),
.B(n_20),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_456),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_430),
.Y(n_658)
);

BUFx8_ASAP7_75t_SL g659 ( 
.A(n_491),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_463),
.Y(n_660)
);

OA21x2_ASAP7_75t_L g661 ( 
.A1(n_465),
.A2(n_21),
.B(n_22),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_472),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_474),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_482),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_486),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_577),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_580),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_599),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_R g669 ( 
.A(n_586),
.B(n_487),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_567),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_594),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_605),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_585),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_636),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_596),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_659),
.Y(n_676)
);

CKINVDCx16_ASAP7_75t_R g677 ( 
.A(n_632),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_637),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_639),
.B(n_410),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_601),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_648),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_623),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_625),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_613),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_567),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_631),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_633),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_650),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_650),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_629),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_629),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_573),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_639),
.B(n_458),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_586),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_597),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_R g698 ( 
.A(n_638),
.B(n_498),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_624),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_638),
.B(n_565),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_639),
.B(n_569),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_566),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_568),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_568),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_645),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_645),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_645),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_641),
.B(n_499),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_576),
.B(n_519),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_593),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_593),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_581),
.Y(n_712)
);

BUFx6f_ASAP7_75t_SL g713 ( 
.A(n_589),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_654),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_570),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_628),
.Y(n_716)
);

INVx6_ASAP7_75t_L g717 ( 
.A(n_629),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_654),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_630),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_628),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_630),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_654),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_590),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_570),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_608),
.A2(n_558),
.B1(n_553),
.B2(n_560),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_604),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_609),
.Y(n_727)
);

AOI21x1_ASAP7_75t_L g728 ( 
.A1(n_595),
.A2(n_504),
.B(n_502),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_620),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_660),
.Y(n_730)
);

INVxp33_ASAP7_75t_L g731 ( 
.A(n_630),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_570),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_584),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_634),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_635),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_R g736 ( 
.A(n_651),
.B(n_378),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_575),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_660),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_660),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_621),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_662),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_577),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_583),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_591),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_R g745 ( 
.A(n_651),
.B(n_379),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_589),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_600),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_571),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_572),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_587),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_696),
.B(n_578),
.C(n_643),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_746),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_738),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_749),
.B(n_649),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_712),
.B(n_653),
.C(n_644),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_738),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_734),
.B(n_602),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_737),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_692),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_679),
.B(n_602),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_SL g761 ( 
.A(n_684),
.B(n_532),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_748),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_735),
.B(n_640),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_702),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_677),
.B(n_572),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_692),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_666),
.B(n_640),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_666),
.B(n_647),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_709),
.B(n_647),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_742),
.B(n_603),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_742),
.B(n_603),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_705),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_746),
.B(n_655),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_701),
.B(n_657),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_700),
.B(n_607),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_669),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_712),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_L g778 ( 
.A(n_673),
.B(n_626),
.Y(n_778)
);

BUFx6f_ASAP7_75t_SL g779 ( 
.A(n_693),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_697),
.B(n_607),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_750),
.A2(n_656),
.B1(n_611),
.B2(n_616),
.Y(n_781)
);

BUFx6f_ASAP7_75t_SL g782 ( 
.A(n_719),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_736),
.B(n_611),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_736),
.B(n_616),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_706),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_745),
.B(n_662),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_745),
.B(n_664),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_733),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_701),
.B(n_713),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_707),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_743),
.B(n_665),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_744),
.B(n_663),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_728),
.A2(n_598),
.B(n_574),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_713),
.B(n_658),
.Y(n_794)
);

NAND3xp33_ASAP7_75t_L g795 ( 
.A(n_669),
.B(n_662),
.C(n_617),
.Y(n_795)
);

INVxp33_ASAP7_75t_L g796 ( 
.A(n_672),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_714),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_723),
.B(n_381),
.Y(n_798)
);

INVxp33_ASAP7_75t_L g799 ( 
.A(n_674),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_726),
.B(n_642),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_667),
.Y(n_801)
);

BUFx5_ASAP7_75t_L g802 ( 
.A(n_718),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_747),
.B(n_642),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_671),
.A2(n_606),
.B1(n_627),
.B2(n_617),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_675),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_681),
.Y(n_806)
);

INVx8_ASAP7_75t_L g807 ( 
.A(n_678),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_727),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_729),
.B(n_615),
.Y(n_809)
);

BUFx6f_ASAP7_75t_SL g810 ( 
.A(n_721),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_722),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_683),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_725),
.B(n_509),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_699),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_708),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_730),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_739),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_695),
.B(n_388),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_708),
.B(n_390),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_741),
.B(n_571),
.Y(n_820)
);

BUFx6f_ASAP7_75t_SL g821 ( 
.A(n_676),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_670),
.B(n_571),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_717),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_680),
.B(n_579),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_731),
.B(n_511),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_717),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_686),
.B(n_579),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_685),
.B(n_391),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_682),
.B(n_661),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_690),
.B(n_582),
.C(n_515),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_687),
.B(n_392),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_689),
.B(n_579),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_691),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_717),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_688),
.B(n_393),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_668),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_703),
.B(n_588),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_704),
.A2(n_514),
.B(n_549),
.C(n_535),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_694),
.B(n_394),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_715),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_724),
.B(n_588),
.Y(n_841)
);

AO22x1_ASAP7_75t_L g842 ( 
.A1(n_830),
.A2(n_710),
.B1(n_716),
.B2(n_646),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_764),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_753),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_801),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_788),
.B(n_606),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_762),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_762),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_815),
.B(n_740),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_765),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_776),
.B(n_777),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_808),
.Y(n_852)
);

AND2x4_ASAP7_75t_SL g853 ( 
.A(n_833),
.B(n_711),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_821),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_800),
.B(n_720),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_813),
.A2(n_627),
.B1(n_661),
.B2(n_652),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_762),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_752),
.B(n_698),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_754),
.B(n_646),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_819),
.A2(n_618),
.B(n_652),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_774),
.B(n_646),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_829),
.A2(n_550),
.B1(n_551),
.B2(n_547),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_773),
.A2(n_732),
.B(n_396),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_760),
.B(n_395),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_781),
.B(n_755),
.C(n_751),
.Y(n_865)
);

NOR2x1p5_ASAP7_75t_L g866 ( 
.A(n_769),
.B(n_698),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_836),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_752),
.B(n_389),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_787),
.B(n_398),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_796),
.B(n_402),
.Y(n_870)
);

NOR2x2_ASAP7_75t_L g871 ( 
.A(n_759),
.B(n_22),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_805),
.B(n_403),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_807),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_821),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_752),
.B(n_783),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_806),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_807),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_812),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_766),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_814),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_784),
.B(n_405),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_775),
.B(n_406),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_807),
.B(n_778),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_756),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_772),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_799),
.B(n_407),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_758),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_779),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_785),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_791),
.B(n_792),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_790),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_803),
.B(n_408),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_797),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_798),
.B(n_412),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_811),
.Y(n_895)
);

AND2x4_ASAP7_75t_SL g896 ( 
.A(n_794),
.B(n_748),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_816),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_817),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_779),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_823),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_795),
.A2(n_559),
.B1(n_592),
.B2(n_588),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_770),
.B(n_23),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_820),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_771),
.B(n_413),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_782),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_767),
.B(n_414),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_768),
.B(n_417),
.Y(n_907)
);

BUFx4f_ASAP7_75t_L g908 ( 
.A(n_826),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_840),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_757),
.B(n_23),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_780),
.B(n_24),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_782),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_789),
.B(n_763),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_834),
.Y(n_914)
);

OR2x6_ASAP7_75t_L g915 ( 
.A(n_809),
.B(n_592),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_786),
.B(n_418),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_802),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_822),
.Y(n_918)
);

AO22x1_ASAP7_75t_L g919 ( 
.A1(n_825),
.A2(n_431),
.B1(n_434),
.B2(n_422),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_802),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_828),
.B(n_24),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_810),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_824),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_827),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_793),
.A2(n_436),
.B(n_435),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_838),
.A2(n_818),
.B(n_839),
.C(n_835),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_802),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_804),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_810),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_802),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_832),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_802),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_761),
.B(n_440),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_837),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_841),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_831),
.A2(n_446),
.B1(n_449),
.B2(n_441),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_808),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_815),
.B(n_451),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_815),
.B(n_452),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_764),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_764),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_847),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_865),
.A2(n_459),
.B(n_461),
.C(n_457),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_890),
.B(n_462),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_849),
.B(n_469),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_938),
.A2(n_473),
.B1(n_478),
.B2(n_470),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_L g947 ( 
.A(n_870),
.B(n_484),
.C(n_483),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_852),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_873),
.B(n_26),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_939),
.A2(n_490),
.B1(n_492),
.B2(n_488),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_917),
.A2(n_494),
.B(n_493),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_866),
.B(n_495),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_912),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_937),
.Y(n_954)
);

BUFx4f_ASAP7_75t_L g955 ( 
.A(n_883),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_843),
.A2(n_500),
.B1(n_503),
.B2(n_496),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_851),
.A2(n_508),
.B1(n_510),
.B2(n_505),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_867),
.Y(n_958)
);

BUFx4f_ASAP7_75t_L g959 ( 
.A(n_883),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_894),
.A2(n_517),
.B(n_518),
.C(n_512),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_845),
.A2(n_521),
.B1(n_522),
.B2(n_520),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_850),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_847),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_886),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_877),
.B(n_854),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_858),
.B(n_525),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_926),
.A2(n_528),
.B(n_530),
.C(n_527),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_863),
.A2(n_559),
.B(n_29),
.C(n_26),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_876),
.B(n_534),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_855),
.B(n_28),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_913),
.B(n_536),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_902),
.A2(n_538),
.B(n_539),
.C(n_537),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_910),
.B(n_540),
.Y(n_973)
);

O2A1O1Ixp5_ASAP7_75t_L g974 ( 
.A1(n_881),
.A2(n_559),
.B(n_31),
.C(n_29),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_878),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_847),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_SL g977 ( 
.A(n_874),
.B(n_542),
.Y(n_977)
);

AOI221xp5_ASAP7_75t_L g978 ( 
.A1(n_902),
.A2(n_561),
.B1(n_544),
.B2(n_545),
.C(n_546),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_905),
.B(n_543),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_880),
.B(n_548),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_940),
.B(n_552),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_941),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_853),
.B(n_34),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_864),
.B(n_556),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_857),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_927),
.A2(n_557),
.B1(n_563),
.B2(n_37),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_920),
.A2(n_748),
.B(n_610),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_910),
.B(n_559),
.Y(n_988)
);

OAI21x1_ASAP7_75t_SL g989 ( 
.A1(n_859),
.A2(n_35),
.B(n_36),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_932),
.A2(n_610),
.B(n_592),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_911),
.B(n_921),
.Y(n_991)
);

NAND3xp33_ASAP7_75t_SL g992 ( 
.A(n_936),
.B(n_892),
.C(n_882),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_885),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_930),
.A2(n_612),
.B(n_610),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_897),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_912),
.Y(n_996)
);

NAND2xp33_ASAP7_75t_L g997 ( 
.A(n_861),
.B(n_559),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_889),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_862),
.B(n_38),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_929),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_898),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_860),
.A2(n_57),
.B(n_53),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_915),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_888),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_869),
.B(n_38),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_928),
.B(n_39),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_872),
.A2(n_40),
.B(n_42),
.C(n_622),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_915),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_921),
.A2(n_622),
.B(n_619),
.C(n_614),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_911),
.B(n_935),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_904),
.A2(n_622),
.B(n_619),
.C(n_614),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_R g1012 ( 
.A(n_899),
.B(n_612),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_891),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_925),
.A2(n_614),
.B(n_612),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_875),
.A2(n_619),
.B(n_62),
.C(n_65),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_922),
.B(n_58),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_895),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_964),
.B(n_903),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_1002),
.A2(n_856),
.B(n_901),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_1003),
.B(n_842),
.Y(n_1020)
);

AO21x2_ASAP7_75t_L g1021 ( 
.A1(n_1014),
.A2(n_923),
.B(n_918),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_993),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_958),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_942),
.Y(n_1024)
);

INVx3_ASAP7_75t_SL g1025 ( 
.A(n_996),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_SL g1026 ( 
.A(n_992),
.B(n_857),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_942),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_998),
.Y(n_1028)
);

OA21x2_ASAP7_75t_L g1029 ( 
.A1(n_967),
.A2(n_931),
.B(n_924),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_987),
.A2(n_846),
.B(n_848),
.Y(n_1030)
);

BUFx4f_ASAP7_75t_SL g1031 ( 
.A(n_948),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_997),
.A2(n_933),
.B(n_934),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_942),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1013),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_991),
.B(n_953),
.Y(n_1035)
);

OA21x2_ASAP7_75t_L g1036 ( 
.A1(n_968),
.A2(n_884),
.B(n_909),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_954),
.B(n_887),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_995),
.Y(n_1038)
);

AO21x2_ASAP7_75t_L g1039 ( 
.A1(n_1006),
.A2(n_1005),
.B(n_989),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1001),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_994),
.A2(n_848),
.B(n_844),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_990),
.A2(n_868),
.B(n_916),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_1015),
.A2(n_907),
.B(n_906),
.Y(n_1043)
);

AO21x2_ASAP7_75t_L g1044 ( 
.A1(n_1009),
.A2(n_893),
.B(n_900),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_1004),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_974),
.A2(n_857),
.B(n_893),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1017),
.Y(n_1047)
);

BUFx2_ASAP7_75t_SL g1048 ( 
.A(n_949),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_1010),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_963),
.Y(n_1050)
);

BUFx2_ASAP7_75t_R g1051 ( 
.A(n_973),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_963),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_999),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_963),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_1011),
.A2(n_893),
.B(n_900),
.Y(n_1055)
);

AO21x2_ASAP7_75t_L g1056 ( 
.A1(n_984),
.A2(n_900),
.B(n_879),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_951),
.A2(n_879),
.B(n_914),
.Y(n_1057)
);

OR2x6_ASAP7_75t_L g1058 ( 
.A(n_1008),
.B(n_879),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_976),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_955),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1000),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_976),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_976),
.Y(n_1063)
);

INVx6_ASAP7_75t_L g1064 ( 
.A(n_985),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_985),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_959),
.Y(n_1066)
);

BUFx2_ASAP7_75t_R g1067 ( 
.A(n_988),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_962),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_985),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1007),
.A2(n_908),
.B(n_896),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_969),
.Y(n_1071)
);

INVx3_ASAP7_75t_SL g1072 ( 
.A(n_983),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_1016),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_980),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_970),
.Y(n_1075)
);

INVxp67_ASAP7_75t_SL g1076 ( 
.A(n_975),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_944),
.B(n_919),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_981),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_943),
.A2(n_960),
.B(n_972),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_977),
.B(n_871),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_1012),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_952),
.Y(n_1082)
);

AO21x1_ASAP7_75t_L g1083 ( 
.A1(n_1077),
.A2(n_982),
.B(n_966),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1077),
.A2(n_947),
.B1(n_971),
.B2(n_957),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1022),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1023),
.B(n_979),
.Y(n_1086)
);

CKINVDCx11_ASAP7_75t_R g1087 ( 
.A(n_1025),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1023),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1028),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1080),
.B(n_978),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1034),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1040),
.Y(n_1092)
);

AO21x1_ASAP7_75t_SL g1093 ( 
.A1(n_1079),
.A2(n_945),
.B(n_986),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1031),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1031),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_1061),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1071),
.A2(n_961),
.B1(n_956),
.B2(n_950),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1047),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1040),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1045),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1074),
.A2(n_946),
.B1(n_965),
.B2(n_70),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1068),
.A2(n_66),
.B1(n_69),
.B2(n_73),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1025),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1038),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1018),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1056),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1064),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1018),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1037),
.B(n_373),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1036),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1053),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1078),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1072),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1076),
.A2(n_1075),
.B1(n_1073),
.B2(n_1049),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1076),
.A2(n_75),
.B(n_77),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1049),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1054),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_1064),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1059),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1064),
.Y(n_1120)
);

BUFx4f_ASAP7_75t_L g1121 ( 
.A(n_1060),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1048),
.B(n_78),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1061),
.B(n_371),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1036),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1024),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1021),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1032),
.A2(n_79),
.B(n_83),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1021),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1041),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1066),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1062),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1032),
.A2(n_1030),
.B(n_1046),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1079),
.A2(n_85),
.B(n_86),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1072),
.B(n_90),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1075),
.B(n_368),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1069),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_1070),
.A2(n_91),
.B(n_92),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1082),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1058),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1058),
.B(n_94),
.Y(n_1140)
);

AOI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1029),
.A2(n_1019),
.B(n_1055),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1073),
.A2(n_96),
.B1(n_100),
.B2(n_105),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_1020),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1044),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1019),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1085),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_1087),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1090),
.B(n_1020),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_SL g1149 ( 
.A(n_1100),
.B(n_1051),
.C(n_1039),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1088),
.B(n_1020),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1104),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1088),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_1094),
.B(n_1058),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_1087),
.B(n_1081),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1094),
.B(n_1035),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1100),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_R g1157 ( 
.A(n_1086),
.B(n_1035),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1089),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_R g1159 ( 
.A(n_1113),
.B(n_1029),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_R g1160 ( 
.A(n_1121),
.B(n_1095),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_R g1161 ( 
.A(n_1121),
.B(n_1081),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1130),
.B(n_1050),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_1084),
.B(n_1051),
.C(n_1039),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1130),
.B(n_1050),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1104),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_R g1166 ( 
.A(n_1122),
.B(n_1024),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1105),
.B(n_1063),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1092),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1108),
.B(n_1027),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_1143),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_1103),
.B(n_1081),
.Y(n_1171)
);

OAI222xp33_ASAP7_75t_L g1172 ( 
.A1(n_1101),
.A2(n_1081),
.B1(n_1065),
.B2(n_1063),
.C1(n_1067),
.C2(n_1052),
.Y(n_1172)
);

OR2x6_ASAP7_75t_L g1173 ( 
.A(n_1140),
.B(n_1027),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1101),
.B(n_1026),
.C(n_1067),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1092),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1116),
.B(n_1033),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1103),
.B(n_1033),
.Y(n_1177)
);

CKINVDCx16_ASAP7_75t_R g1178 ( 
.A(n_1143),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_R g1179 ( 
.A(n_1118),
.B(n_1052),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1109),
.B(n_1056),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_1115),
.A2(n_1043),
.B(n_1057),
.C(n_1042),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1091),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1096),
.B(n_1044),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_1114),
.Y(n_1184)
);

XNOR2xp5_ASAP7_75t_L g1185 ( 
.A(n_1134),
.B(n_1138),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1097),
.A2(n_116),
.B1(n_118),
.B2(n_121),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1123),
.B(n_122),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1112),
.B(n_125),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1107),
.B(n_126),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1098),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1107),
.Y(n_1191)
);

CKINVDCx16_ASAP7_75t_R g1192 ( 
.A(n_1120),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1132),
.A2(n_128),
.B(n_132),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1111),
.B(n_367),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1118),
.B(n_133),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1126),
.A2(n_1128),
.A3(n_1144),
.B(n_1137),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1083),
.A2(n_134),
.B1(n_138),
.B2(n_142),
.Y(n_1197)
);

OA21x2_ASAP7_75t_L g1198 ( 
.A1(n_1132),
.A2(n_143),
.B(n_145),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1107),
.B(n_150),
.Y(n_1199)
);

XNOR2xp5_ASAP7_75t_L g1200 ( 
.A(n_1114),
.B(n_151),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1099),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1107),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1120),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1117),
.B(n_152),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1139),
.B(n_1125),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1125),
.B(n_153),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1119),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1099),
.Y(n_1208)
);

AOI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1133),
.A2(n_154),
.B(n_155),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1125),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_1135),
.B(n_159),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1131),
.B(n_160),
.Y(n_1212)
);

CKINVDCx6p67_ASAP7_75t_R g1213 ( 
.A(n_1125),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1136),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1097),
.B(n_161),
.Y(n_1215)
);

NAND2xp33_ASAP7_75t_R g1216 ( 
.A(n_1144),
.B(n_162),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1142),
.B(n_164),
.Y(n_1217)
);

OAI33xp33_ASAP7_75t_L g1218 ( 
.A1(n_1146),
.A2(n_1093),
.A3(n_1110),
.B1(n_1124),
.B2(n_1128),
.B3(n_1126),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1150),
.B(n_1106),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1148),
.B(n_1106),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1207),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1191),
.Y(n_1222)
);

OR2x6_ASAP7_75t_SL g1223 ( 
.A(n_1176),
.B(n_1110),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1152),
.B(n_1145),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1170),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1158),
.B(n_1124),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1185),
.B(n_1145),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1167),
.B(n_1102),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1182),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1190),
.B(n_1141),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1153),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1183),
.B(n_1129),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1214),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1196),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1201),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1198),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1169),
.B(n_1129),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1184),
.B(n_167),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1208),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1168),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1175),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1178),
.B(n_1127),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1180),
.B(n_168),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1151),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1173),
.B(n_169),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1196),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1173),
.B(n_171),
.Y(n_1247)
);

AND4x1_ASAP7_75t_L g1248 ( 
.A(n_1215),
.B(n_1163),
.C(n_1149),
.D(n_1197),
.Y(n_1248)
);

INVx5_ASAP7_75t_SL g1249 ( 
.A(n_1153),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1202),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1162),
.B(n_173),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1165),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1171),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1210),
.B(n_174),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1159),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1192),
.B(n_176),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1213),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1162),
.B(n_178),
.Y(n_1258)
);

AO21x2_ASAP7_75t_L g1259 ( 
.A1(n_1181),
.A2(n_181),
.B(n_183),
.Y(n_1259)
);

NOR2x1_ASAP7_75t_L g1260 ( 
.A(n_1155),
.B(n_185),
.Y(n_1260)
);

NOR2x1_ASAP7_75t_SL g1261 ( 
.A(n_1164),
.B(n_186),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1164),
.B(n_188),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1155),
.B(n_189),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1205),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1177),
.B(n_191),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1198),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1188),
.B(n_1200),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1193),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1204),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1200),
.B(n_192),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1194),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1203),
.B(n_197),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1212),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1217),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1187),
.B(n_198),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1217),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1160),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1199),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1174),
.B(n_199),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1211),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1186),
.A2(n_200),
.B(n_201),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1189),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1147),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1179),
.B(n_1206),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1189),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1195),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1154),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1221),
.B(n_1156),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1230),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1220),
.B(n_1209),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1239),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1229),
.B(n_1161),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1219),
.B(n_1157),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1233),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1274),
.A2(n_1172),
.B(n_1166),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1235),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1239),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1226),
.Y(n_1298)
);

AND2x4_ASAP7_75t_SL g1299 ( 
.A(n_1285),
.B(n_1216),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1222),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1232),
.B(n_202),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1274),
.B(n_203),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1252),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1237),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1244),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1244),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1240),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1240),
.Y(n_1308)
);

BUFx2_ASAP7_75t_SL g1309 ( 
.A(n_1222),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1276),
.B(n_205),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1241),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1276),
.B(n_206),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1269),
.B(n_207),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1267),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1242),
.B(n_211),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1250),
.B(n_366),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1241),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1271),
.B(n_213),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1223),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1271),
.B(n_1286),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1232),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1223),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1250),
.B(n_363),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1232),
.B(n_214),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1286),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1224),
.B(n_215),
.Y(n_1326)
);

NOR2x1_ASAP7_75t_L g1327 ( 
.A(n_1287),
.B(n_217),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1273),
.B(n_220),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1234),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1278),
.B(n_1255),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1255),
.B(n_1234),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1227),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.C(n_226),
.Y(n_1332)
);

OA211x2_ASAP7_75t_L g1333 ( 
.A1(n_1284),
.A2(n_227),
.B(n_230),
.C(n_231),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1246),
.B(n_234),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_L g1335 ( 
.A(n_1280),
.B(n_235),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1246),
.B(n_236),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1278),
.B(n_237),
.Y(n_1337)
);

AOI21xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1256),
.A2(n_238),
.B(n_240),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1231),
.B(n_361),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1225),
.B(n_241),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1266),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1327),
.B(n_1280),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1289),
.B(n_1282),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1320),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1294),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1341),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1289),
.B(n_1236),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1331),
.B(n_1330),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1309),
.B(n_1283),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1331),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1300),
.B(n_1283),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1296),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1321),
.B(n_1236),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1304),
.B(n_1298),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1288),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1303),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1319),
.B(n_1264),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1329),
.Y(n_1358)
);

NOR3xp33_ASAP7_75t_L g1359 ( 
.A(n_1302),
.B(n_1218),
.C(n_1285),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1341),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1293),
.B(n_1277),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1322),
.B(n_1228),
.Y(n_1362)
);

INVxp33_ASAP7_75t_L g1363 ( 
.A(n_1315),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1290),
.B(n_1253),
.Y(n_1364)
);

AOI211x1_ASAP7_75t_SL g1365 ( 
.A1(n_1314),
.A2(n_1268),
.B(n_1272),
.C(n_1266),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1321),
.B(n_1285),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1290),
.B(n_1257),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1325),
.B(n_1243),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1292),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1297),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1315),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1291),
.Y(n_1372)
);

AOI21xp33_ASAP7_75t_L g1373 ( 
.A1(n_1295),
.A2(n_1279),
.B(n_1238),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1291),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1310),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1326),
.B(n_1236),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1375),
.B(n_1334),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1342),
.B(n_1302),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1348),
.B(n_1299),
.Y(n_1379)
);

O2A1O1Ixp5_ASAP7_75t_R g1380 ( 
.A1(n_1343),
.A2(n_1318),
.B(n_1333),
.C(n_1340),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1349),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1370),
.Y(n_1382)
);

NOR4xp25_ASAP7_75t_L g1383 ( 
.A(n_1371),
.B(n_1373),
.C(n_1369),
.D(n_1355),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1348),
.B(n_1299),
.Y(n_1384)
);

OAI32xp33_ASAP7_75t_L g1385 ( 
.A1(n_1363),
.A2(n_1312),
.A3(n_1270),
.B1(n_1326),
.B2(n_1313),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1370),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1362),
.B(n_1350),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1348),
.B(n_1257),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1358),
.B(n_1305),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1358),
.Y(n_1390)
);

OAI322xp33_ASAP7_75t_L g1391 ( 
.A1(n_1345),
.A2(n_1247),
.A3(n_1338),
.B1(n_1328),
.B2(n_1263),
.C1(n_1317),
.C2(n_1334),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1364),
.B(n_1336),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1363),
.A2(n_1258),
.B1(n_1251),
.B2(n_1335),
.Y(n_1393)
);

AOI33xp33_ASAP7_75t_L g1394 ( 
.A1(n_1352),
.A2(n_1328),
.A3(n_1332),
.B1(n_1336),
.B2(n_1339),
.B3(n_1265),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1344),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1356),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1359),
.A2(n_1218),
.B1(n_1243),
.B2(n_1275),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1379),
.B(n_1367),
.Y(n_1398)
);

NAND2xp33_ASAP7_75t_SL g1399 ( 
.A(n_1381),
.B(n_1351),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1378),
.A2(n_1342),
.B1(n_1368),
.B2(n_1357),
.Y(n_1400)
);

NAND3xp33_ASAP7_75t_L g1401 ( 
.A(n_1397),
.B(n_1347),
.C(n_1376),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1395),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1378),
.A2(n_1361),
.B1(n_1376),
.B2(n_1337),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1380),
.A2(n_1347),
.B1(n_1366),
.B2(n_1353),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1396),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1383),
.A2(n_1385),
.B(n_1394),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1377),
.A2(n_1354),
.B1(n_1324),
.B2(n_1301),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1393),
.A2(n_1366),
.B1(n_1301),
.B2(n_1324),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1387),
.A2(n_1366),
.B1(n_1353),
.B2(n_1245),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1379),
.A2(n_1260),
.B1(n_1245),
.B2(n_1316),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1389),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1390),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1405),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1402),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1406),
.B(n_1382),
.Y(n_1415)
);

NOR4xp25_ASAP7_75t_L g1416 ( 
.A(n_1400),
.B(n_1391),
.C(n_1386),
.D(n_1392),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1411),
.B(n_1365),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1404),
.B(n_1384),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1412),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1401),
.A2(n_1360),
.B1(n_1374),
.B2(n_1388),
.Y(n_1420)
);

NAND2x1_ASAP7_75t_SL g1421 ( 
.A(n_1403),
.B(n_1245),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1398),
.Y(n_1422)
);

OAI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1408),
.A2(n_1248),
.B1(n_1374),
.B2(n_1372),
.C(n_1360),
.Y(n_1423)
);

INVx4_ASAP7_75t_L g1424 ( 
.A(n_1399),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1409),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1410),
.B(n_1257),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1407),
.A2(n_1281),
.B(n_1323),
.C(n_1360),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1405),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1415),
.B(n_1374),
.Y(n_1429)
);

NOR2x1_ASAP7_75t_L g1430 ( 
.A(n_1424),
.B(n_1259),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1416),
.A2(n_1261),
.B(n_1281),
.Y(n_1431)
);

AOI211xp5_ASAP7_75t_L g1432 ( 
.A1(n_1416),
.A2(n_1257),
.B(n_1262),
.C(n_1254),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1417),
.A2(n_1372),
.B1(n_1346),
.B2(n_1259),
.C(n_1268),
.Y(n_1433)
);

AOI211xp5_ASAP7_75t_L g1434 ( 
.A1(n_1427),
.A2(n_1346),
.B(n_1311),
.C(n_1308),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1424),
.B(n_1249),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1421),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1422),
.B(n_1249),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_L g1438 ( 
.A(n_1414),
.B(n_1249),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1432),
.A2(n_1423),
.B1(n_1418),
.B2(n_1425),
.Y(n_1439)
);

AOI211xp5_ASAP7_75t_L g1440 ( 
.A1(n_1431),
.A2(n_1420),
.B(n_1426),
.C(n_1413),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_L g1441 ( 
.A(n_1435),
.B(n_1438),
.Y(n_1441)
);

AO22x2_ASAP7_75t_L g1442 ( 
.A1(n_1436),
.A2(n_1428),
.B1(n_1419),
.B2(n_1311),
.Y(n_1442)
);

NOR2x1_ASAP7_75t_L g1443 ( 
.A(n_1430),
.B(n_1306),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1429),
.Y(n_1444)
);

OAI211xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1433),
.A2(n_1308),
.B(n_1307),
.C(n_1306),
.Y(n_1445)
);

AND4x2_ASAP7_75t_L g1446 ( 
.A(n_1441),
.B(n_1434),
.C(n_1437),
.D(n_244),
.Y(n_1446)
);

NAND4xp25_ASAP7_75t_L g1447 ( 
.A(n_1440),
.B(n_1307),
.C(n_243),
.D(n_247),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1444),
.A2(n_1445),
.B(n_1443),
.C(n_1442),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1439),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1444),
.B(n_242),
.Y(n_1450)
);

AOI222xp33_ASAP7_75t_L g1451 ( 
.A1(n_1445),
.A2(n_249),
.B1(n_254),
.B2(n_256),
.C1(n_257),
.C2(n_258),
.Y(n_1451)
);

AOI31xp33_ASAP7_75t_L g1452 ( 
.A1(n_1449),
.A2(n_259),
.A3(n_261),
.B(n_265),
.Y(n_1452)
);

NOR2x1_ASAP7_75t_L g1453 ( 
.A(n_1447),
.B(n_270),
.Y(n_1453)
);

NOR4xp25_ASAP7_75t_L g1454 ( 
.A(n_1448),
.B(n_1450),
.C(n_1446),
.D(n_1451),
.Y(n_1454)
);

AO211x2_ASAP7_75t_L g1455 ( 
.A1(n_1447),
.A2(n_271),
.B(n_273),
.C(n_274),
.Y(n_1455)
);

INVxp33_ASAP7_75t_SL g1456 ( 
.A(n_1450),
.Y(n_1456)
);

NOR2x1_ASAP7_75t_L g1457 ( 
.A(n_1447),
.B(n_276),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1447),
.A2(n_281),
.B1(n_283),
.B2(n_286),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1454),
.A2(n_288),
.B(n_289),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1453),
.B(n_1457),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1458),
.B(n_1456),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1452),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1455),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1456),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1462),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1464),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1464),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1460),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1461),
.Y(n_1469)
);

NAND2xp33_ASAP7_75t_SL g1470 ( 
.A(n_1466),
.B(n_1463),
.Y(n_1470)
);

AND4x1_ASAP7_75t_L g1471 ( 
.A(n_1469),
.B(n_1459),
.C(n_291),
.D(n_292),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1467),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_L g1473 ( 
.A(n_1465),
.B(n_290),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1468),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1470),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1474),
.Y(n_1476)
);

AOI31xp33_ASAP7_75t_L g1477 ( 
.A1(n_1472),
.A2(n_298),
.A3(n_299),
.B(n_304),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1473),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1471),
.A2(n_305),
.B1(n_309),
.B2(n_311),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1476),
.B(n_312),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1478),
.A2(n_313),
.B1(n_317),
.B2(n_319),
.Y(n_1481)
);

AOI22x1_ASAP7_75t_L g1482 ( 
.A1(n_1475),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1477),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1479),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1483),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_1485)
);

XNOR2xp5_ASAP7_75t_L g1486 ( 
.A(n_1480),
.B(n_326),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1484),
.B(n_328),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1482),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1488),
.B(n_1486),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1487),
.A2(n_1481),
.B(n_333),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1490),
.A2(n_1489),
.B1(n_1485),
.B2(n_338),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1491),
.B(n_332),
.Y(n_1492)
);

AOI211xp5_ASAP7_75t_L g1493 ( 
.A1(n_1492),
.A2(n_334),
.B(n_342),
.C(n_346),
.Y(n_1493)
);


endmodule