module real_aes_7486_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_310;
wire n_119;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g427 ( .A(n_0), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_1), .A2(n_125), .B(n_129), .C(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_2), .A2(n_154), .B(n_155), .Y(n_153) );
INVx1_ASAP7_75t_L g531 ( .A(n_3), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_4), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_4), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_5), .B(n_166), .Y(n_165) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_6), .A2(n_154), .B(n_498), .Y(n_497) );
AND2x6_ASAP7_75t_L g125 ( .A(n_7), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g271 ( .A(n_8), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_9), .B(n_41), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_10), .A2(n_175), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_11), .B(n_137), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_12), .B(n_159), .Y(n_486) );
INVx1_ASAP7_75t_L g502 ( .A(n_13), .Y(n_502) );
INVx1_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
INVx1_ASAP7_75t_L g456 ( .A(n_15), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_16), .A2(n_135), .B(n_227), .C(n_229), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_17), .B(n_166), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_18), .B(n_466), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_19), .B(n_154), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_20), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_21), .A2(n_159), .B(n_236), .C(n_238), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_22), .B(n_166), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_23), .B(n_137), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_24), .A2(n_182), .B(n_229), .C(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_25), .B(n_137), .Y(n_136) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_26), .Y(n_190) );
INVx1_ASAP7_75t_L g133 ( .A(n_27), .Y(n_133) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_28), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_29), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_30), .B(n_137), .Y(n_532) );
INVx1_ASAP7_75t_L g180 ( .A(n_31), .Y(n_180) );
INVx1_ASAP7_75t_L g510 ( .A(n_32), .Y(n_510) );
INVx2_ASAP7_75t_L g123 ( .A(n_33), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_34), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_35), .A2(n_159), .B(n_160), .C(n_162), .Y(n_158) );
INVxp67_ASAP7_75t_L g181 ( .A(n_36), .Y(n_181) );
CKINVDCx14_ASAP7_75t_R g156 ( .A(n_37), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g128 ( .A1(n_38), .A2(n_129), .B(n_132), .C(n_140), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_39), .A2(n_125), .B(n_129), .C(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_40), .A2(n_70), .B1(n_722), .B2(n_723), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_40), .Y(n_722) );
INVx1_ASAP7_75t_L g509 ( .A(n_42), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_43), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_44), .A2(n_198), .B(n_269), .C(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_45), .B(n_137), .Y(n_474) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_46), .A2(n_86), .B1(n_109), .B2(n_110), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_46), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_47), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_48), .Y(n_177) );
INVx1_ASAP7_75t_L g234 ( .A(n_49), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_50), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_51), .B(n_154), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_52), .A2(n_721), .B1(n_724), .B2(n_725), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_52), .Y(n_725) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_53), .A2(n_442), .B1(n_716), .B2(n_717), .C1(n_726), .C2(n_727), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_54), .A2(n_129), .B1(n_238), .B2(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_55), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_56), .Y(n_528) );
CKINVDCx14_ASAP7_75t_R g267 ( .A(n_57), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_58), .A2(n_162), .B(n_269), .C(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_59), .Y(n_477) );
INVx1_ASAP7_75t_L g499 ( .A(n_60), .Y(n_499) );
INVx1_ASAP7_75t_L g126 ( .A(n_61), .Y(n_126) );
INVx1_ASAP7_75t_L g144 ( .A(n_62), .Y(n_144) );
INVx1_ASAP7_75t_SL g161 ( .A(n_63), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_64), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_65), .B(n_166), .Y(n_240) );
INVx1_ASAP7_75t_L g193 ( .A(n_66), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_SL g518 ( .A1(n_67), .A2(n_162), .B(n_466), .C(n_519), .Y(n_518) );
INVxp67_ASAP7_75t_L g520 ( .A(n_68), .Y(n_520) );
INVx1_ASAP7_75t_L g439 ( .A(n_69), .Y(n_439) );
INVx1_ASAP7_75t_L g723 ( .A(n_70), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_71), .A2(n_154), .B(n_266), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_72), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_73), .A2(n_154), .B(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_74), .Y(n_513) );
INVx1_ASAP7_75t_L g471 ( .A(n_75), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_76), .A2(n_175), .B(n_176), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g225 ( .A(n_78), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_79), .A2(n_125), .B(n_129), .C(n_473), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_80), .A2(n_154), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g228 ( .A(n_81), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_82), .B(n_134), .Y(n_464) );
INVx2_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g217 ( .A(n_84), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_85), .B(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_86), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_87), .A2(n_125), .B(n_129), .C(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g424 ( .A(n_88), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g711 ( .A(n_88), .Y(n_711) );
OR2x2_ASAP7_75t_L g715 ( .A(n_88), .B(n_426), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_89), .A2(n_129), .B(n_192), .C(n_200), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_90), .B(n_141), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_91), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_92), .A2(n_125), .B(n_129), .C(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g419 ( .A1(n_93), .A2(n_99), .B1(n_420), .B2(n_421), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_93), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_94), .Y(n_490) );
INVx1_ASAP7_75t_L g517 ( .A(n_95), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_96), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_97), .B(n_134), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_98), .B(n_149), .Y(n_272) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_99), .A2(n_104), .B1(n_432), .B2(n_440), .C1(n_728), .C2(n_733), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_99), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_99), .B(n_149), .Y(n_457) );
INVx2_ASAP7_75t_L g237 ( .A(n_100), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_101), .B(n_439), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_102), .A2(n_154), .B(n_516), .Y(n_515) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_423), .B(n_429), .Y(n_105) );
OAI22xp33_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_418), .B1(n_419), .B2(n_422), .Y(n_106) );
INVx1_ASAP7_75t_L g422 ( .A(n_107), .Y(n_422) );
XOR2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g712 ( .A(n_111), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_111), .A2(n_444), .B1(n_710), .B2(n_715), .Y(n_726) );
OR3x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_329), .C(n_376), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_275), .C(n_300), .Y(n_112) );
AOI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_210), .B1(n_241), .B2(n_244), .C(n_252), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_167), .B(n_203), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_116), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_116), .B(n_257), .Y(n_373) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_151), .Y(n_116) );
AND2x2_ASAP7_75t_L g243 ( .A(n_117), .B(n_209), .Y(n_243) );
AND2x2_ASAP7_75t_L g293 ( .A(n_117), .B(n_208), .Y(n_293) );
AND2x2_ASAP7_75t_L g314 ( .A(n_117), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_117), .B(n_286), .Y(n_319) );
OR2x2_ASAP7_75t_L g327 ( .A(n_117), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g399 ( .A(n_117), .B(n_187), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_117), .B(n_348), .Y(n_413) );
INVx3_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g258 ( .A(n_118), .B(n_151), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_118), .B(n_187), .Y(n_259) );
AND2x4_ASAP7_75t_L g281 ( .A(n_118), .B(n_209), .Y(n_281) );
AND2x2_ASAP7_75t_L g311 ( .A(n_118), .B(n_169), .Y(n_311) );
AND2x2_ASAP7_75t_L g320 ( .A(n_118), .B(n_310), .Y(n_320) );
AND2x2_ASAP7_75t_L g336 ( .A(n_118), .B(n_188), .Y(n_336) );
OR2x2_ASAP7_75t_L g345 ( .A(n_118), .B(n_328), .Y(n_345) );
AND2x2_ASAP7_75t_L g351 ( .A(n_118), .B(n_286), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_118), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g365 ( .A(n_118), .B(n_205), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_118), .B(n_254), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_118), .B(n_315), .Y(n_404) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_146), .Y(n_118) );
O2A1O1Ixp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_127), .B(n_128), .C(n_141), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_120), .A2(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_120), .A2(n_214), .B(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_120), .A2(n_471), .B(n_472), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_120), .A2(n_164), .B1(n_507), .B2(n_511), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_120), .A2(n_528), .B(n_529), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g120 ( .A(n_121), .B(n_125), .Y(n_120) );
AND2x4_ASAP7_75t_L g154 ( .A(n_121), .B(n_125), .Y(n_154) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g139 ( .A(n_122), .Y(n_139) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g130 ( .A(n_123), .Y(n_130) );
INVx1_ASAP7_75t_L g239 ( .A(n_123), .Y(n_239) );
INVx1_ASAP7_75t_L g131 ( .A(n_124), .Y(n_131) );
INVx3_ASAP7_75t_L g135 ( .A(n_124), .Y(n_135) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_124), .Y(n_137) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_124), .Y(n_183) );
INVx1_ASAP7_75t_L g466 ( .A(n_124), .Y(n_466) );
BUFx3_ASAP7_75t_L g140 ( .A(n_125), .Y(n_140) );
INVx4_ASAP7_75t_SL g164 ( .A(n_125), .Y(n_164) );
INVx5_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
AND2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
BUFx3_ASAP7_75t_L g199 ( .A(n_130), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B(n_136), .C(n_138), .Y(n_132) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_134), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_134), .A2(n_531), .B(n_532), .C(n_533), .Y(n_530) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_135), .B(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_135), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_135), .B(n_520), .Y(n_519) );
INVx4_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
INVx2_ASAP7_75t_L g269 ( .A(n_137), .Y(n_269) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_139), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
INVx1_ASAP7_75t_L g212 ( .A(n_141), .Y(n_212) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_141), .A2(n_265), .B(n_272), .Y(n_264) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_141), .A2(n_451), .B(n_457), .Y(n_450) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g150 ( .A(n_142), .B(n_143), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx3_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_148), .A2(n_189), .B(n_201), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_148), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_SL g467 ( .A(n_148), .B(n_468), .Y(n_467) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_149), .A2(n_515), .B(n_521), .Y(n_514) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
INVx2_ASAP7_75t_L g209 ( .A(n_151), .Y(n_209) );
AND2x2_ASAP7_75t_L g310 ( .A(n_151), .B(n_187), .Y(n_310) );
AND2x2_ASAP7_75t_L g315 ( .A(n_151), .B(n_188), .Y(n_315) );
INVx1_ASAP7_75t_L g371 ( .A(n_151), .Y(n_371) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_165), .Y(n_151) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_152), .A2(n_223), .B(n_230), .Y(n_222) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_152), .A2(n_232), .B(n_240), .Y(n_231) );
BUFx2_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_158), .C(n_164), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_157), .A2(n_164), .B(n_177), .C(n_178), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g224 ( .A1(n_157), .A2(n_164), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_157), .A2(n_164), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_157), .A2(n_164), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_157), .A2(n_164), .B(n_453), .C(n_454), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_157), .A2(n_164), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_157), .A2(n_164), .B(n_517), .C(n_518), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_159), .B(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_163), .Y(n_487) );
INVx1_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_166), .A2(n_497), .B(n_503), .Y(n_496) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g280 ( .A(n_168), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_187), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_169), .B(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g257 ( .A(n_169), .Y(n_257) );
OR2x2_ASAP7_75t_L g328 ( .A(n_169), .B(n_187), .Y(n_328) );
OR2x2_ASAP7_75t_L g389 ( .A(n_169), .B(n_296), .Y(n_389) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_174), .B(n_184), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_171), .A2(n_206), .B(n_207), .Y(n_205) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_171), .A2(n_470), .B(n_476), .Y(n_469) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_SL g460 ( .A1(n_172), .A2(n_461), .B(n_462), .Y(n_460) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_173), .A2(n_506), .B(n_512), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_173), .B(n_513), .Y(n_512) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_173), .A2(n_527), .B(n_534), .Y(n_526) );
INVx1_ASAP7_75t_L g206 ( .A(n_174), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_182), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_182), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_182), .B(n_456), .Y(n_455) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g195 ( .A(n_183), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g508 ( .A1(n_183), .A2(n_195), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g207 ( .A(n_184), .Y(n_207) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_186), .B(n_202), .Y(n_201) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_186), .A2(n_482), .B(n_489), .Y(n_481) );
AND2x2_ASAP7_75t_L g208 ( .A(n_187), .B(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g348 ( .A(n_187), .B(n_205), .Y(n_348) );
INVx2_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
BUFx2_ASAP7_75t_L g287 ( .A(n_188), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_L g216 ( .A1(n_194), .A2(n_197), .B(n_217), .C(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_197), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_197), .A2(n_474), .B(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_204), .A2(n_393), .B1(n_397), .B2(n_400), .C(n_401), .Y(n_392) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_208), .Y(n_204) );
INVx1_ASAP7_75t_SL g255 ( .A(n_205), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_205), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g387 ( .A(n_205), .B(n_243), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_208), .B(n_257), .Y(n_379) );
AND2x2_ASAP7_75t_L g286 ( .A(n_209), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_SL g290 ( .A(n_210), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_210), .B(n_296), .Y(n_326) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_221), .Y(n_210) );
AND2x2_ASAP7_75t_L g251 ( .A(n_211), .B(n_222), .Y(n_251) );
INVx4_ASAP7_75t_L g263 ( .A(n_211), .Y(n_263) );
BUFx3_ASAP7_75t_L g306 ( .A(n_211), .Y(n_306) );
AND3x2_ASAP7_75t_L g321 ( .A(n_211), .B(n_322), .C(n_323), .Y(n_321) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_219), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_212), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_212), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_212), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g403 ( .A(n_221), .B(n_317), .Y(n_403) );
AND2x2_ASAP7_75t_L g411 ( .A(n_221), .B(n_296), .Y(n_411) );
INVx1_ASAP7_75t_SL g416 ( .A(n_221), .Y(n_416) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_231), .Y(n_221) );
INVx1_ASAP7_75t_SL g274 ( .A(n_222), .Y(n_274) );
AND2x2_ASAP7_75t_L g297 ( .A(n_222), .B(n_263), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_222), .B(n_247), .Y(n_299) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_222), .Y(n_339) );
OR2x2_ASAP7_75t_L g344 ( .A(n_222), .B(n_263), .Y(n_344) );
INVx2_ASAP7_75t_L g249 ( .A(n_231), .Y(n_249) );
AND2x2_ASAP7_75t_L g284 ( .A(n_231), .B(n_264), .Y(n_284) );
OR2x2_ASAP7_75t_L g304 ( .A(n_231), .B(n_264), .Y(n_304) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_231), .Y(n_324) );
INVx2_ASAP7_75t_L g533 ( .A(n_238), .Y(n_533) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AOI21xp33_ASAP7_75t_L g374 ( .A1(n_242), .A2(n_283), .B(n_375), .Y(n_374) );
AOI322xp5_ASAP7_75t_L g410 ( .A1(n_244), .A2(n_254), .A3(n_281), .B1(n_411), .B2(n_412), .C1(n_414), .C2(n_417), .Y(n_410) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_246), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_247), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g273 ( .A(n_248), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g341 ( .A(n_249), .B(n_263), .Y(n_341) );
AND2x2_ASAP7_75t_L g408 ( .A(n_249), .B(n_264), .Y(n_408) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g349 ( .A(n_251), .B(n_303), .Y(n_349) );
AOI31xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_256), .A3(n_259), .B(n_260), .Y(n_252) );
AND2x2_ASAP7_75t_L g308 ( .A(n_254), .B(n_286), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_254), .B(n_278), .Y(n_390) );
AND2x2_ASAP7_75t_L g409 ( .A(n_254), .B(n_314), .Y(n_409) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_257), .B(n_286), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_257), .B(n_315), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_257), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_257), .B(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_258), .B(n_315), .Y(n_347) );
INVx1_ASAP7_75t_L g391 ( .A(n_258), .Y(n_391) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_273), .Y(n_261) );
INVxp67_ASAP7_75t_L g343 ( .A(n_262), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_263), .B(n_274), .Y(n_279) );
INVx1_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_263), .B(n_362), .Y(n_396) );
BUFx3_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
AND2x2_ASAP7_75t_L g322 ( .A(n_264), .B(n_274), .Y(n_322) );
INVx2_ASAP7_75t_L g362 ( .A(n_264), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_273), .B(n_395), .Y(n_394) );
AOI211xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B(n_282), .C(n_291), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_277), .A2(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_278), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_278), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g358 ( .A(n_279), .B(n_304), .Y(n_358) );
INVx3_ASAP7_75t_L g289 ( .A(n_281), .Y(n_289) );
OAI22xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_285), .B1(n_288), .B2(n_290), .Y(n_282) );
OAI21xp5_ASAP7_75t_SL g307 ( .A1(n_284), .A2(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g333 ( .A(n_284), .B(n_297), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_284), .B(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g288 ( .A(n_287), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g357 ( .A(n_287), .Y(n_357) );
OAI21xp5_ASAP7_75t_SL g301 ( .A1(n_288), .A2(n_302), .B(n_307), .Y(n_301) );
OAI22xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_294), .B1(n_298), .B2(n_299), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_293), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_296), .B(n_339), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_312), .C(n_325), .Y(n_300) );
OAI22xp5_ASAP7_75t_SL g367 ( .A1(n_302), .A2(n_368), .B1(n_372), .B2(n_373), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g372 ( .A(n_304), .B(n_305), .Y(n_372) );
AND2x2_ASAP7_75t_L g380 ( .A(n_305), .B(n_361), .Y(n_380) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_306), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_SL g388 ( .A1(n_306), .A2(n_389), .B(n_390), .C(n_391), .Y(n_388) );
OR2x2_ASAP7_75t_L g415 ( .A(n_306), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B(n_318), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_314), .A2(n_351), .B(n_352), .C(n_355), .Y(n_350) );
OAI21xp33_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_320), .B(n_321), .Y(n_318) );
AND2x2_ASAP7_75t_L g383 ( .A(n_322), .B(n_341), .Y(n_383) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
NAND3xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_350), .C(n_363), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_334), .C(n_342), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g400 ( .A(n_337), .Y(n_400) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g360 ( .A(n_339), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_339), .B(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B(n_345), .C(n_346), .Y(n_342) );
INVx2_ASAP7_75t_SL g354 ( .A(n_344), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_345), .A2(n_356), .B1(n_358), .B2(n_359), .Y(n_355) );
OAI21xp33_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_348), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
AOI211xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B(n_367), .C(n_374), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVxp33_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g417 ( .A(n_371), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_392), .C(n_405), .D(n_410), .Y(n_376) );
AOI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_381), .C(n_388), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_386), .Y(n_381) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_382), .A2(n_402), .B(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_389), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_409), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_424), .Y(n_431) );
INVx1_ASAP7_75t_SL g732 ( .A(n_424), .Y(n_732) );
BUFx2_ASAP7_75t_L g735 ( .A(n_424), .Y(n_735) );
NOR2x2_ASAP7_75t_L g727 ( .A(n_425), .B(n_711), .Y(n_727) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g710 ( .A(n_426), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_SL g730 ( .A(n_436), .B(n_438), .Y(n_730) );
OA21x2_ASAP7_75t_L g734 ( .A1(n_436), .A2(n_437), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_708), .B1(n_712), .B2(n_713), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
OR4x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_604), .C(n_663), .D(n_690), .Y(n_444) );
NAND3xp33_ASAP7_75t_SL g445 ( .A(n_446), .B(n_546), .C(n_571), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_478), .B(n_495), .C(n_522), .Y(n_446) );
AOI211xp5_ASAP7_75t_SL g694 ( .A1(n_447), .A2(n_695), .B(n_697), .C(n_700), .Y(n_694) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_458), .Y(n_447) );
INVx1_ASAP7_75t_L g569 ( .A(n_448), .Y(n_569) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g544 ( .A(n_449), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g576 ( .A(n_449), .Y(n_576) );
AND2x2_ASAP7_75t_L g631 ( .A(n_449), .B(n_600), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_449), .B(n_493), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_449), .B(n_494), .Y(n_689) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g550 ( .A(n_450), .Y(n_550) );
AND2x2_ASAP7_75t_L g593 ( .A(n_450), .B(n_469), .Y(n_593) );
AND2x2_ASAP7_75t_L g611 ( .A(n_450), .B(n_494), .Y(n_611) );
INVx4_ASAP7_75t_L g543 ( .A(n_458), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_458), .A2(n_599), .B(n_601), .Y(n_598) );
AND2x2_ASAP7_75t_L g679 ( .A(n_458), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_469), .Y(n_458) );
INVx1_ASAP7_75t_L g492 ( .A(n_459), .Y(n_492) );
AND2x2_ASAP7_75t_L g548 ( .A(n_459), .B(n_494), .Y(n_548) );
OR2x2_ASAP7_75t_L g577 ( .A(n_459), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g591 ( .A(n_459), .Y(n_591) );
INVx3_ASAP7_75t_L g600 ( .A(n_459), .Y(n_600) );
AND2x2_ASAP7_75t_L g610 ( .A(n_459), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g643 ( .A(n_459), .B(n_549), .Y(n_643) );
AND2x2_ASAP7_75t_L g667 ( .A(n_459), .B(n_623), .Y(n_667) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
INVx2_ASAP7_75t_L g494 ( .A(n_469), .Y(n_494) );
AND2x2_ASAP7_75t_L g703 ( .A(n_469), .B(n_545), .Y(n_703) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_480), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g623 ( .A(n_480), .B(n_611), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_480), .B(n_600), .Y(n_685) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g545 ( .A(n_481), .Y(n_545) );
AND2x2_ASAP7_75t_L g549 ( .A(n_481), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g590 ( .A(n_481), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_488), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_487), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_491), .B(n_586), .Y(n_608) );
INVx1_ASAP7_75t_L g647 ( .A(n_491), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_491), .B(n_574), .Y(n_691) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
AND2x2_ASAP7_75t_L g554 ( .A(n_492), .B(n_549), .Y(n_554) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_494), .B(n_545), .Y(n_578) );
INVx1_ASAP7_75t_L g657 ( .A(n_494), .Y(n_657) );
AOI322xp5_ASAP7_75t_L g681 ( .A1(n_495), .A2(n_596), .A3(n_656), .B1(n_682), .B2(n_684), .C1(n_686), .C2(n_688), .Y(n_681) );
AND2x2_ASAP7_75t_SL g495 ( .A(n_496), .B(n_504), .Y(n_495) );
AND2x2_ASAP7_75t_L g536 ( .A(n_496), .B(n_514), .Y(n_536) );
INVx1_ASAP7_75t_SL g539 ( .A(n_496), .Y(n_539) );
AND2x2_ASAP7_75t_L g541 ( .A(n_496), .B(n_505), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_496), .B(n_558), .Y(n_564) );
INVx2_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
AND2x2_ASAP7_75t_L g596 ( .A(n_496), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_558), .Y(n_634) );
BUFx2_ASAP7_75t_L g651 ( .A(n_496), .Y(n_651) );
AND2x2_ASAP7_75t_L g665 ( .A(n_496), .B(n_525), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_504), .B(n_553), .Y(n_580) );
AND2x2_ASAP7_75t_L g707 ( .A(n_504), .B(n_583), .Y(n_707) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
OR2x2_ASAP7_75t_L g552 ( .A(n_505), .B(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g558 ( .A(n_505), .Y(n_558) );
AND2x2_ASAP7_75t_L g603 ( .A(n_505), .B(n_526), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_505), .B(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_505), .Y(n_687) );
AND2x2_ASAP7_75t_L g538 ( .A(n_514), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
BUFx2_ASAP7_75t_L g566 ( .A(n_514), .Y(n_566) );
AND2x2_ASAP7_75t_L g585 ( .A(n_514), .B(n_558), .Y(n_585) );
INVx3_ASAP7_75t_L g597 ( .A(n_514), .Y(n_597) );
OR2x2_ASAP7_75t_L g607 ( .A(n_514), .B(n_558), .Y(n_607) );
AOI31xp33_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_537), .A3(n_540), .B(n_542), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_536), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_524), .B(n_559), .Y(n_570) );
OR2x2_ASAP7_75t_L g594 ( .A(n_524), .B(n_564), .Y(n_594) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_525), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g615 ( .A(n_525), .B(n_607), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_525), .B(n_597), .Y(n_625) );
AND2x2_ASAP7_75t_L g632 ( .A(n_525), .B(n_633), .Y(n_632) );
NAND2x1_ASAP7_75t_L g660 ( .A(n_525), .B(n_596), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_525), .B(n_651), .Y(n_661) );
AND2x2_ASAP7_75t_L g673 ( .A(n_525), .B(n_558), .Y(n_673) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g553 ( .A(n_526), .Y(n_553) );
INVx1_ASAP7_75t_L g619 ( .A(n_536), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_536), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_538), .B(n_614), .Y(n_648) );
AND2x4_ASAP7_75t_L g559 ( .A(n_539), .B(n_560), .Y(n_559) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g638 ( .A(n_544), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_544), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g586 ( .A(n_545), .B(n_576), .Y(n_586) );
AND2x2_ASAP7_75t_L g680 ( .A(n_545), .B(n_550), .Y(n_680) );
INVx1_ASAP7_75t_L g705 ( .A(n_545), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_551), .B1(n_554), .B2(n_555), .C(n_561), .Y(n_546) );
CKINVDCx14_ASAP7_75t_R g567 ( .A(n_547), .Y(n_567) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_548), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_551), .B(n_602), .Y(n_621) );
INVx3_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g670 ( .A(n_552), .B(n_566), .Y(n_670) );
AND2x2_ASAP7_75t_L g584 ( .A(n_553), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g614 ( .A(n_553), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_553), .B(n_597), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_553), .B(n_654), .C(n_685), .Y(n_684) );
AOI211xp5_ASAP7_75t_SL g617 ( .A1(n_554), .A2(n_618), .B(n_620), .C(n_628), .Y(n_617) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_556), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_557), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_557), .B(n_641), .Y(n_640) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g699 ( .A(n_559), .B(n_673), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_567), .B1(n_568), .B2(n_570), .Y(n_561) );
NOR2xp33_ASAP7_75t_SL g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_565), .B(n_614), .Y(n_645) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_568), .A2(n_660), .B1(n_691), .B2(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_579), .B1(n_581), .B2(n_586), .C(n_587), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_577), .A2(n_588), .B1(n_594), .B2(n_595), .C(n_598), .Y(n_587) );
INVx1_ASAP7_75t_L g630 ( .A(n_578), .Y(n_630) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_SL g602 ( .A(n_583), .Y(n_602) );
OR2x2_ASAP7_75t_L g675 ( .A(n_583), .B(n_607), .Y(n_675) );
AND2x2_ASAP7_75t_L g677 ( .A(n_583), .B(n_585), .Y(n_677) );
INVx1_ASAP7_75t_L g616 ( .A(n_586), .Y(n_616) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
AOI21xp33_ASAP7_75t_SL g646 ( .A1(n_589), .A2(n_647), .B(n_648), .Y(n_646) );
OR2x2_ASAP7_75t_L g653 ( .A(n_589), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g627 ( .A(n_590), .B(n_611), .Y(n_627) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp33_ASAP7_75t_SL g644 ( .A(n_595), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_596), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_597), .B(n_633), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_600), .A2(n_613), .B(n_615), .C(n_616), .Y(n_612) );
NAND2x1_ASAP7_75t_SL g637 ( .A(n_600), .B(n_638), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_601), .A2(n_650), .B1(n_652), .B2(n_655), .Y(n_649) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_603), .B(n_693), .Y(n_692) );
NAND5xp2_ASAP7_75t_L g604 ( .A(n_605), .B(n_617), .C(n_635), .D(n_649), .E(n_658), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_612), .Y(n_605) );
INVx1_ASAP7_75t_L g662 ( .A(n_608), .Y(n_662) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_610), .A2(n_629), .B1(n_669), .B2(n_671), .C(n_674), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_611), .B(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_614), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_614), .B(n_680), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_624), .B2(n_626), .Y(n_620) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g702 ( .A(n_631), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_639), .B1(n_643), .B2(n_644), .C(n_646), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g686 ( .A(n_641), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g693 ( .A(n_651), .Y(n_693) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_661), .B(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_666), .B(n_668), .C(n_681), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_666), .A2(n_691), .B(n_692), .C(n_694), .Y(n_690) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_670), .B(n_672), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_704), .B(n_706), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g724 ( .A(n_721), .Y(n_724) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
NAND2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
endmodule