module fake_netlist_5_1264_n_1942 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1942);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1942;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_999;
wire n_758;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g192 ( 
.A(n_56),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_64),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_68),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_177),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_17),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_34),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_34),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_78),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_127),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_73),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_33),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_59),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_33),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_31),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_4),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_142),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_36),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_87),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_35),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_159),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_90),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_121),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_4),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_0),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_58),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_110),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_151),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_104),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_84),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_24),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_5),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_158),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_77),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_147),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_18),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_44),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_115),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_108),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_52),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_162),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_89),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_106),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_141),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_128),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_21),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_86),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_120),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_83),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_51),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_79),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_45),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_19),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_43),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_100),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_98),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_143),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_61),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_118),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_136),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_66),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_59),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_102),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_80),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_116),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_18),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_186),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_81),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_9),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_173),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_146),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_138),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_49),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_145),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_139),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_67),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_119),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_17),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_7),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_144),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_168),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_71),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_0),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_135),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_19),
.Y(n_294)
);

BUFx8_ASAP7_75t_SL g295 ( 
.A(n_36),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_107),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_190),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_179),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_15),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_54),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_70),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_149),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_65),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_130),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_72),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_22),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_8),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_76),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_16),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_5),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_171),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_6),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_40),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_55),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_44),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_31),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_46),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_47),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_21),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_69),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_37),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_7),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_112),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_39),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_103),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_63),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_12),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_175),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_155),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_114),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_2),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_153),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_99),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_46),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_11),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_178),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_58),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_30),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_97),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_95),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_150),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_181),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_189),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_50),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_137),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_92),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_75),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_187),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_29),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_109),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_93),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_51),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_88),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_32),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_191),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_10),
.Y(n_358)
);

BUFx2_ASAP7_75t_SL g359 ( 
.A(n_49),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_161),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_48),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_22),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_74),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_32),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_169),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_156),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_1),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_85),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_1),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_29),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_39),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_160),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_41),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_165),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_28),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_14),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_176),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_117),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_96),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_61),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_43),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_63),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_82),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_229),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_295),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_229),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_208),
.B(n_2),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_259),
.B(n_3),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_229),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_229),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_238),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_202),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_250),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_229),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_255),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_294),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_208),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_348),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_244),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_294),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_294),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_284),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_248),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_294),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_252),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_294),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_256),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_264),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_265),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_193),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_268),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_193),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_206),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_206),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_260),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_260),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_272),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_383),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_233),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_291),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_301),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_306),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_301),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_211),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_213),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_198),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_192),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_275),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_210),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_214),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_278),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_236),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_313),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_345),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_242),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_254),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_280),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_253),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_283),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_270),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_277),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_286),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_259),
.B(n_3),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_297),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_211),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_287),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_200),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_298),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_374),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_288),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_303),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_377),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_305),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_245),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_311),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_316),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_320),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_245),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_307),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_199),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_310),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_198),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_322),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_327),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_330),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_329),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_333),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_339),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_331),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_326),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_259),
.A2(n_6),
.B(n_9),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_335),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_347),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_346),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_354),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_199),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_349),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_358),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_387),
.B(n_249),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_384),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_220),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_388),
.B(n_249),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_390),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

AND2x4_ASAP7_75t_SL g494 ( 
.A(n_463),
.B(n_205),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_464),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_220),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_387),
.B(n_267),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_423),
.B(n_267),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_445),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_471),
.A2(n_257),
.B(n_226),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_445),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_404),
.B(n_226),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_404),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_460),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_443),
.B(n_205),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_471),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_410),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_423),
.B(n_296),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_421),
.B(n_296),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_429),
.B(n_343),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_430),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_476),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_432),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_435),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_413),
.B(n_343),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_413),
.A2(n_341),
.B(n_257),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_435),
.B(n_194),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_414),
.B(n_341),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_415),
.B(n_201),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_438),
.B(n_194),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_440),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_440),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_415),
.B(n_292),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_416),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_416),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_478),
.B(n_292),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_441),
.B(n_195),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_446),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_446),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_450),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_450),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_453),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_453),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_455),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_489),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_489),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_479),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_479),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_498),
.Y(n_564)
);

NOR2x1p5_ASAP7_75t_L g565 ( 
.A(n_490),
.B(n_385),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_483),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

NOR2x1p5_ASAP7_75t_L g569 ( 
.A(n_490),
.B(n_419),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_491),
.B(n_391),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_483),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_528),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_485),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_498),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_486),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_493),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_495),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_487),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_L g585 ( 
.A(n_511),
.B(n_447),
.C(n_470),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_498),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_498),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_498),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_488),
.Y(n_590)
);

BUFx6f_ASAP7_75t_SL g591 ( 
.A(n_522),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_502),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_508),
.B(n_399),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_497),
.A2(n_398),
.B1(n_418),
.B2(n_324),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_497),
.A2(n_324),
.B1(n_362),
.B2(n_359),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_511),
.A2(n_302),
.B1(n_315),
.B2(n_300),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_504),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_520),
.B(n_403),
.Y(n_599)
);

NOR2x1p5_ASAP7_75t_L g600 ( 
.A(n_536),
.B(n_207),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_504),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_504),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_496),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_514),
.B(n_405),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_491),
.B(n_407),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_491),
.B(n_482),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_520),
.B(n_426),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_503),
.B(n_455),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_491),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_520),
.A2(n_361),
.B1(n_319),
.B2(n_241),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_502),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_530),
.A2(n_215),
.B1(n_225),
.B2(n_218),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_541),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_508),
.B(n_408),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_492),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_480),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_502),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_541),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_541),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_482),
.A2(n_478),
.B1(n_475),
.B2(n_474),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_482),
.B(n_409),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_514),
.B(n_216),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_500),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_500),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_501),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_499),
.B(n_411),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_512),
.B(n_417),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_499),
.B(n_428),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_512),
.A2(n_452),
.B1(n_472),
.B2(n_477),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_514),
.B(n_224),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_528),
.B(n_431),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_499),
.B(n_437),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_541),
.B(n_230),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_530),
.Y(n_638)
);

BUFx6f_ASAP7_75t_SL g639 ( 
.A(n_522),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_480),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_L g641 ( 
.A(n_538),
.B(n_462),
.C(n_271),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_502),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_496),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_480),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_536),
.B(n_439),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_509),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_519),
.B(n_442),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_481),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_502),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_502),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_519),
.B(n_444),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_481),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_507),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_538),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_542),
.B(n_448),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_481),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_542),
.B(n_451),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_459),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_519),
.B(n_461),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_505),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_507),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_519),
.B(n_465),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_481),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_505),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_513),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_550),
.B(n_469),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_550),
.B(n_473),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_494),
.A2(n_436),
.B1(n_449),
.B2(n_309),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_513),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_524),
.A2(n_247),
.B1(n_269),
.B2(n_274),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_503),
.B(n_475),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_507),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_494),
.B(n_205),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_509),
.Y(n_675)
);

INVxp33_ASAP7_75t_SL g676 ( 
.A(n_503),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_514),
.B(n_195),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_507),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_509),
.Y(n_679)
);

CKINVDCx6p67_ASAP7_75t_R g680 ( 
.A(n_522),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_507),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_SL g682 ( 
.A1(n_524),
.A2(n_342),
.B1(n_304),
.B2(n_281),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_515),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_494),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_515),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_494),
.B(n_285),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_507),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_527),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_553),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_527),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_527),
.Y(n_691)
);

BUFx6f_ASAP7_75t_SL g692 ( 
.A(n_522),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_507),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_527),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_522),
.B(n_392),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_553),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_531),
.B(n_285),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_553),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_549),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_531),
.B(n_285),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_549),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_553),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_484),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_534),
.B(n_239),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_553),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_553),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_534),
.B(n_276),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_614),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_606),
.A2(n_514),
.B1(n_433),
.B2(n_434),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_599),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_676),
.B(n_332),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_558),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_656),
.B(n_514),
.Y(n_715)
);

AO22x2_ASAP7_75t_L g716 ( 
.A1(n_686),
.A2(n_234),
.B1(n_237),
.B2(n_240),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_658),
.B(n_514),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_607),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_619),
.Y(n_719)
);

NOR2x1p5_ASAP7_75t_L g720 ( 
.A(n_684),
.B(n_207),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_572),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_607),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_700),
.B(n_553),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_700),
.B(n_531),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_624),
.B(n_211),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_702),
.B(n_578),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_676),
.A2(n_395),
.B1(n_393),
.B2(n_402),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_702),
.B(n_534),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_578),
.B(n_534),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_619),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_609),
.B(n_569),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_569),
.A2(n_420),
.B1(n_422),
.B2(n_350),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_609),
.B(n_534),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_567),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_558),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_677),
.A2(n_518),
.B(n_556),
.C(n_555),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_572),
.B(n_549),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_620),
.B(n_211),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_620),
.B(n_698),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_698),
.B(n_211),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_567),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_665),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_680),
.A2(n_293),
.B1(n_243),
.B2(n_251),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_629),
.B(n_510),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_562),
.B(n_510),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_623),
.B(n_211),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_562),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_559),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_563),
.B(n_566),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_563),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_559),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_566),
.B(n_510),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_628),
.B(n_211),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_638),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_571),
.B(n_510),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_L g756 ( 
.A1(n_596),
.A2(n_521),
.B1(n_556),
.B2(n_555),
.C(n_554),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_608),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_655),
.B(n_545),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_655),
.B(n_545),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_674),
.A2(n_632),
.B1(n_669),
.B2(n_684),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_571),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_573),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_573),
.B(n_510),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_672),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_575),
.B(n_539),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_672),
.B(n_545),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_631),
.B(n_211),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_636),
.B(n_217),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_575),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_634),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_576),
.B(n_539),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_576),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_577),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_577),
.B(n_539),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_624),
.B(n_217),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_580),
.B(n_539),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_595),
.B(n_246),
.C(n_235),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_580),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_591),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_583),
.B(n_539),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_583),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_590),
.B(n_527),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_703),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_634),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_703),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_590),
.B(n_527),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_586),
.A2(n_506),
.B(n_535),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_196),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_610),
.B(n_540),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_610),
.B(n_540),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_665),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_616),
.B(n_540),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_638),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_600),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_616),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_680),
.A2(n_263),
.B1(n_273),
.B2(n_325),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_570),
.B(n_506),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_667),
.B(n_196),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_560),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_637),
.B(n_217),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_695),
.A2(n_289),
.B1(n_203),
.B2(n_204),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_600),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_540),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_682),
.A2(n_521),
.B(n_554),
.C(n_525),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_621),
.B(n_540),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_625),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_625),
.B(n_626),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_626),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_637),
.B(n_217),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_682),
.A2(n_518),
.B(n_525),
.C(n_551),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_627),
.B(n_540),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_605),
.A2(n_652),
.B1(n_659),
.B2(n_648),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_627),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_560),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_668),
.B(n_660),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_630),
.B(n_540),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_613),
.B(n_622),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_663),
.B(n_197),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_630),
.B(n_546),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_674),
.B(n_334),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_706),
.B(n_709),
.C(n_641),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_637),
.B(n_217),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_637),
.B(n_217),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_613),
.B(n_523),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_624),
.A2(n_506),
.B1(n_535),
.B2(n_217),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_661),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_661),
.B(n_546),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_617),
.Y(n_829)
);

AND2x6_ASAP7_75t_SL g830 ( 
.A(n_603),
.B(n_456),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_666),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_624),
.B(n_217),
.Y(n_832)
);

BUFx6f_ASAP7_75t_SL g833 ( 
.A(n_643),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_666),
.B(n_338),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_671),
.B(n_197),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_646),
.B(n_675),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_670),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_591),
.A2(n_344),
.B1(n_363),
.B2(n_368),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_683),
.B(n_546),
.Y(n_839)
);

BUFx5_ASAP7_75t_L g840 ( 
.A(n_624),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_546),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_685),
.B(n_618),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_703),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_635),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_635),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_697),
.B(n_701),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_685),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_689),
.B(n_203),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_568),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_689),
.B(n_204),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_703),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_699),
.B(n_209),
.Y(n_852)
);

NOR2x1p5_ASAP7_75t_L g853 ( 
.A(n_643),
.B(n_212),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_561),
.B(n_546),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_561),
.B(n_546),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_568),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_561),
.B(n_546),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_585),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_579),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_604),
.A2(n_535),
.B(n_557),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_640),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_611),
.B(n_209),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_640),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_587),
.B(n_547),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_699),
.B(n_219),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_707),
.B(n_219),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_707),
.B(n_221),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_594),
.B(n_261),
.C(n_258),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_567),
.B(n_221),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_SL g870 ( 
.A1(n_597),
.A2(n_228),
.B1(n_225),
.B2(n_218),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_615),
.B(n_222),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_579),
.A2(n_364),
.B1(n_228),
.B2(n_356),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_587),
.B(n_547),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_644),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_587),
.B(n_547),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_591),
.B(n_222),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_593),
.B(n_547),
.Y(n_877)
);

AOI22x1_ASAP7_75t_L g878 ( 
.A1(n_565),
.A2(n_523),
.B1(n_551),
.B2(n_544),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_715),
.B(n_624),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_717),
.B(n_624),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_718),
.B(n_565),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_723),
.A2(n_654),
.B(n_651),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_847),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_847),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_793),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_742),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_793),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_729),
.A2(n_654),
.B(n_651),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_742),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_815),
.A2(n_642),
.B(n_593),
.C(n_681),
.Y(n_890)
);

AOI21xp33_ASAP7_75t_L g891 ( 
.A1(n_713),
.A2(n_266),
.B(n_262),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_785),
.Y(n_892)
);

OAI321xp33_ASAP7_75t_L g893 ( 
.A1(n_862),
.A2(n_456),
.A3(n_474),
.B1(n_468),
.B2(n_467),
.C(n_466),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_791),
.Y(n_894)
);

OAI21xp33_ASAP7_75t_L g895 ( 
.A1(n_713),
.A2(n_356),
.B(n_212),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_787),
.A2(n_612),
.B(n_593),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_791),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_812),
.B(n_815),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_747),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_726),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_733),
.A2(n_654),
.B(n_651),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_860),
.A2(n_633),
.B(n_612),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_817),
.A2(n_544),
.B(n_543),
.C(n_537),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_728),
.B(n_633),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_744),
.A2(n_662),
.B(n_647),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_835),
.A2(n_529),
.B(n_532),
.C(n_533),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_785),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_724),
.B(n_633),
.Y(n_908)
);

AND2x2_ASAP7_75t_SL g909 ( 
.A(n_820),
.B(n_696),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_SL g910 ( 
.A1(n_746),
.A2(n_690),
.B(n_688),
.C(n_704),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_820),
.B(n_612),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_835),
.A2(n_543),
.B(n_537),
.C(n_533),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_SL g913 ( 
.A(n_785),
.B(n_646),
.Y(n_913)
);

AOI21xp33_ASAP7_75t_L g914 ( 
.A1(n_788),
.A2(n_282),
.B(n_279),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_757),
.B(n_764),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_714),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_735),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_842),
.A2(n_741),
.B(n_734),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_712),
.B(n_639),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_750),
.B(n_633),
.Y(n_920)
);

INVx5_ASAP7_75t_L g921 ( 
.A(n_785),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_748),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_746),
.A2(n_767),
.B(n_753),
.Y(n_923)
);

NAND2x1_ASAP7_75t_L g924 ( 
.A(n_783),
.B(n_642),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_751),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_761),
.B(n_762),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_851),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_759),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_769),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_772),
.B(n_633),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_754),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_779),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_783),
.A2(n_662),
.B(n_647),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_722),
.B(n_639),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_773),
.B(n_633),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_766),
.B(n_642),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_778),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_781),
.B(n_633),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_795),
.B(n_681),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_766),
.B(n_681),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_806),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_711),
.A2(n_639),
.B1(n_692),
.B2(n_687),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_797),
.A2(n_693),
.B(n_687),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_753),
.A2(n_768),
.B(n_767),
.C(n_738),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_799),
.Y(n_945)
);

CKINVDCx10_ASAP7_75t_R g946 ( 
.A(n_833),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_770),
.B(n_692),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_843),
.A2(n_662),
.B(n_647),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_797),
.A2(n_693),
.B(n_687),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_843),
.A2(n_647),
.B(n_564),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_721),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_808),
.B(n_693),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_851),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_739),
.A2(n_771),
.B(n_765),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_737),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_788),
.A2(n_688),
.B(n_704),
.C(n_690),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_862),
.A2(n_457),
.B(n_466),
.C(n_467),
.Y(n_957)
);

AO22x1_ASAP7_75t_L g958 ( 
.A1(n_871),
.A2(n_373),
.B1(n_364),
.B2(n_367),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_814),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_813),
.B(n_564),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_731),
.A2(n_692),
.B1(n_564),
.B2(n_567),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_739),
.B(n_696),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_SL g963 ( 
.A1(n_768),
.A2(n_809),
.B(n_822),
.C(n_800),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_804),
.A2(n_457),
.B(n_468),
.C(n_367),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_710),
.B(n_548),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_738),
.A2(n_708),
.B(n_696),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_774),
.A2(n_564),
.B(n_696),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_826),
.B(n_567),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_784),
.B(n_326),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_776),
.A2(n_780),
.B(n_749),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_831),
.B(n_574),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_840),
.B(n_574),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_837),
.B(n_807),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_818),
.B(n_574),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_827),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_858),
.B(n_574),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_854),
.A2(n_708),
.B(n_574),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_824),
.B(n_821),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_818),
.B(n_719),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_730),
.B(n_548),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_798),
.B(n_589),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_798),
.B(n_589),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_797),
.A2(n_602),
.B(n_601),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_846),
.B(n_589),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_727),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_846),
.B(n_589),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_736),
.B(n_589),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_760),
.B(n_360),
.C(n_227),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_849),
.B(n_650),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_825),
.A2(n_650),
.B1(n_673),
.B2(n_678),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_855),
.A2(n_708),
.B(n_678),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_871),
.B(n_371),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_825),
.A2(n_602),
.B(n_601),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_745),
.A2(n_592),
.B(n_598),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_856),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_732),
.B(n_371),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_859),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_779),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_752),
.B(n_650),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_857),
.A2(n_708),
.B(n_678),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_840),
.B(n_650),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_829),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_755),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_844),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_763),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_848),
.A2(n_650),
.B1(n_673),
.B2(n_678),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_801),
.B(n_552),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_794),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_802),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_779),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_845),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_777),
.B(n_673),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_864),
.A2(n_673),
.B(n_678),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_870),
.B(n_552),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_873),
.A2(n_673),
.B(n_703),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_740),
.A2(n_598),
.B(n_592),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_876),
.B(n_557),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_868),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_740),
.A2(n_694),
.B(n_691),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_834),
.B(n_705),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_848),
.B(n_299),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_833),
.Y(n_1022)
);

AND2x6_ASAP7_75t_L g1023 ( 
.A(n_851),
.B(n_691),
.Y(n_1023)
);

OAI321xp33_ASAP7_75t_L g1024 ( 
.A1(n_872),
.A2(n_516),
.A3(n_517),
.B1(n_381),
.B2(n_373),
.C(n_382),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_850),
.A2(n_865),
.B(n_866),
.C(n_867),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_782),
.A2(n_694),
.B(n_705),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_850),
.B(n_308),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_L g1028 ( 
.A(n_756),
.B(n_705),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_840),
.B(n_646),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_875),
.A2(n_675),
.B(n_646),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_840),
.B(n_646),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_877),
.A2(n_675),
.B(n_646),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_852),
.A2(n_223),
.B1(n_227),
.B2(n_231),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_852),
.A2(n_223),
.B1(n_231),
.B2(n_352),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_840),
.B(n_675),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_834),
.B(n_581),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_786),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_810),
.A2(n_370),
.B(n_369),
.C(n_375),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_865),
.A2(n_867),
.B(n_866),
.C(n_869),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_830),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_861),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_720),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_716),
.A2(n_380),
.B(n_382),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_743),
.B(n_312),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_851),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_863),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_853),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_716),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_R g1049 ( 
.A(n_725),
.B(n_232),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_L g1050 ( 
.A(n_878),
.B(n_796),
.C(n_838),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_874),
.B(n_581),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_800),
.A2(n_588),
.B(n_584),
.C(n_582),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_789),
.A2(n_679),
.B(n_675),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_809),
.A2(n_588),
.B(n_582),
.C(n_649),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_716),
.A2(n_232),
.B1(n_290),
.B2(n_357),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_SL g1056 ( 
.A(n_840),
.B(n_352),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_822),
.B(n_644),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_823),
.B(n_353),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_823),
.B(n_369),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_790),
.B(n_649),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_792),
.A2(n_679),
.B(n_675),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_803),
.A2(n_664),
.B(n_657),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_805),
.A2(n_664),
.B(n_657),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_811),
.B(n_653),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_816),
.A2(n_653),
.B(n_679),
.Y(n_1065)
);

INVx8_ASAP7_75t_L g1066 ( 
.A(n_1023),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_899),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_929),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_900),
.B(n_819),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_896),
.A2(n_841),
.B(n_839),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_921),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_937),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_932),
.B(n_828),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_889),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_970),
.A2(n_832),
.B(n_775),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_941),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_887),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_978),
.A2(n_355),
.B(n_353),
.C(n_379),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_SL g1079 ( 
.A1(n_919),
.A2(n_516),
.B(n_517),
.C(n_526),
.Y(n_1079)
);

AOI21x1_ASAP7_75t_L g1080 ( 
.A1(n_879),
.A2(n_526),
.B(n_517),
.Y(n_1080)
);

OAI21xp33_ASAP7_75t_SL g1081 ( 
.A1(n_898),
.A2(n_909),
.B(n_978),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_988),
.A2(n_898),
.B1(n_1027),
.B2(n_1021),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_887),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_L g1084 ( 
.A(n_914),
.B(n_891),
.C(n_1044),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_981),
.A2(n_836),
.B(n_679),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_894),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_982),
.A2(n_836),
.B(n_679),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_L g1088 ( 
.A(n_1044),
.B(n_988),
.C(n_1021),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_900),
.B(n_516),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_892),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_932),
.B(n_526),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_903),
.A2(n_526),
.B(n_547),
.C(n_336),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_946),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_974),
.A2(n_355),
.B(n_357),
.C(n_360),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1027),
.A2(n_1025),
.B(n_1039),
.C(n_992),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_885),
.B(n_314),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_1010),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_919),
.A2(n_378),
.B(n_366),
.C(n_372),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_979),
.A2(n_366),
.B(n_365),
.C(n_378),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1022),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_902),
.A2(n_880),
.B(n_954),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_921),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_915),
.B(n_365),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_886),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_915),
.B(n_379),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_973),
.B(n_547),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_897),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1063),
.A2(n_509),
.B(n_679),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_955),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_895),
.B(n_381),
.C(n_380),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_975),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_903),
.A2(n_547),
.B(n_337),
.C(n_328),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_906),
.A2(n_340),
.B(n_318),
.C(n_321),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_906),
.A2(n_351),
.B(n_323),
.C(n_317),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_928),
.B(n_376),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_L g1116 ( 
.A1(n_890),
.A2(n_509),
.B(n_484),
.C(n_188),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_912),
.A2(n_376),
.B(n_375),
.C(n_370),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_928),
.B(n_484),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_926),
.B(n_484),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_995),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_1042),
.B(n_484),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1048),
.A2(n_509),
.B1(n_484),
.B2(n_12),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1002),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_931),
.B(n_10),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_997),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_977),
.A2(n_509),
.B(n_484),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_909),
.A2(n_185),
.B1(n_184),
.B2(n_180),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1004),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_904),
.A2(n_990),
.B(n_963),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1017),
.A2(n_509),
.B1(n_13),
.B2(n_14),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_976),
.B(n_509),
.Y(n_1131)
);

O2A1O1Ixp5_ASAP7_75t_L g1132 ( 
.A1(n_956),
.A2(n_509),
.B(n_167),
.C(n_152),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1011),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_912),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_984),
.A2(n_140),
.B1(n_132),
.B2(n_129),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_883),
.B(n_126),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1041),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_976),
.B(n_16),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_931),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_951),
.B(n_20),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1046),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_985),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_916),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_951),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_1009),
.B(n_125),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1003),
.B(n_20),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_964),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_892),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_917),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_922),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_963),
.A2(n_113),
.B(n_111),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_1047),
.B(n_123),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_986),
.A2(n_884),
.B1(n_987),
.B2(n_908),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_969),
.B(n_25),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_925),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_921),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1018),
.B(n_105),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_945),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_918),
.A2(n_94),
.B(n_91),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1050),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_911),
.A2(n_101),
.B1(n_30),
.B2(n_37),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1005),
.B(n_27),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_881),
.B(n_38),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_983),
.A2(n_38),
.B(n_40),
.Y(n_1164)
);

NAND2x1_ASAP7_75t_L g1165 ( 
.A(n_1023),
.B(n_41),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_944),
.A2(n_42),
.B(n_45),
.C(n_47),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_964),
.A2(n_42),
.B(n_48),
.C(n_52),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_959),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_965),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_965),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_905),
.A2(n_53),
.B(n_54),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1008),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_1008),
.B(n_55),
.Y(n_1173)
);

CKINVDCx6p67_ASAP7_75t_R g1174 ( 
.A(n_1040),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1037),
.B(n_56),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_SL g1176 ( 
.A(n_998),
.B(n_57),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_980),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_980),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_SL g1179 ( 
.A1(n_1012),
.A2(n_57),
.B(n_60),
.C(n_62),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1059),
.B(n_1007),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1014),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_892),
.Y(n_1182)
);

OR2x6_ASAP7_75t_SL g1183 ( 
.A(n_1055),
.B(n_60),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_882),
.A2(n_62),
.B(n_65),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_996),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_993),
.A2(n_66),
.B(n_1065),
.Y(n_1186)
);

BUFx4f_ASAP7_75t_SL g1187 ( 
.A(n_911),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1051),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_934),
.B(n_947),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1012),
.A2(n_1038),
.B(n_1058),
.C(n_957),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_991),
.A2(n_1000),
.B(n_1013),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_SL g1192 ( 
.A(n_1043),
.B(n_1024),
.C(n_934),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1028),
.A2(n_962),
.B1(n_960),
.B2(n_942),
.Y(n_1193)
);

INVxp67_ASAP7_75t_SL g1194 ( 
.A(n_892),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_939),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_907),
.B(n_953),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_998),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_952),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_958),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_907),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1036),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_957),
.B(n_1038),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_936),
.B(n_940),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_L g1204 ( 
.A(n_927),
.B(n_1045),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1026),
.A2(n_967),
.B(n_943),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_L g1206 ( 
.A(n_1033),
.B(n_1034),
.C(n_893),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_949),
.A2(n_888),
.B(n_901),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_R g1208 ( 
.A(n_927),
.B(n_1045),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_936),
.B(n_1049),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_968),
.A2(n_971),
.B(n_910),
.C(n_935),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_989),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_907),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_907),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_953),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_999),
.A2(n_1056),
.B(n_910),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1020),
.B(n_920),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_953),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_953),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1060),
.A2(n_1064),
.B(n_1062),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_930),
.A2(n_938),
.B(n_1052),
.C(n_1054),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1049),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1015),
.A2(n_994),
.B(n_972),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_972),
.A2(n_1001),
.B(n_950),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1057),
.Y(n_1224)
);

NOR4xp25_ASAP7_75t_L g1225 ( 
.A(n_1088),
.B(n_1006),
.C(n_961),
.D(n_1019),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1215),
.A2(n_923),
.B(n_966),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1084),
.A2(n_1016),
.B(n_948),
.C(n_933),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1067),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1082),
.A2(n_962),
.B1(n_1001),
.B2(n_1023),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1191),
.A2(n_924),
.B(n_1030),
.Y(n_1230)
);

INVxp67_ASAP7_75t_L g1231 ( 
.A(n_1139),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1077),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1075),
.A2(n_921),
.B(n_1031),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1068),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1070),
.A2(n_1223),
.B(n_1080),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1066),
.Y(n_1236)
);

INVx3_ASAP7_75t_SL g1237 ( 
.A(n_1100),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1205),
.A2(n_1061),
.A3(n_1053),
.B(n_1032),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1072),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1076),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1185),
.B(n_1029),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_1205),
.A2(n_1029),
.B(n_1031),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1066),
.B(n_1035),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1180),
.B(n_1023),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1201),
.B(n_1023),
.Y(n_1245)
);

AOI31xp67_ASAP7_75t_L g1246 ( 
.A1(n_1202),
.A2(n_913),
.A3(n_1035),
.B(n_1138),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1223),
.A2(n_1126),
.B(n_1207),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1207),
.A2(n_1222),
.B(n_1108),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1075),
.A2(n_1101),
.B(n_1219),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1101),
.A2(n_1219),
.B(n_1095),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1181),
.B(n_1154),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1120),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1206),
.A2(n_1110),
.B1(n_1187),
.B2(n_1199),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1144),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1129),
.A2(n_1193),
.B(n_1186),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1125),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1186),
.A2(n_1153),
.B(n_1106),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1081),
.A2(n_1114),
.B(n_1113),
.C(n_1190),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1113),
.A2(n_1114),
.B(n_1117),
.C(n_1192),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1116),
.A2(n_1220),
.B(n_1132),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1200),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1127),
.A2(n_1156),
.B(n_1071),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1210),
.A2(n_1119),
.B(n_1102),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1117),
.A2(n_1112),
.B(n_1164),
.C(n_1189),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1210),
.A2(n_1102),
.B(n_1071),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_1166),
.A2(n_1160),
.B(n_1098),
.C(n_1136),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1110),
.A2(n_1179),
.B(n_1078),
.C(n_1163),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1157),
.A2(n_1209),
.B1(n_1142),
.B2(n_1221),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1161),
.A2(n_1135),
.A3(n_1167),
.B1(n_1147),
.B2(n_1134),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1176),
.B(n_1066),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1104),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1107),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_SL g1273 ( 
.A1(n_1164),
.A2(n_1151),
.B(n_1134),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1156),
.A2(n_1085),
.B(n_1087),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1130),
.A2(n_1122),
.B1(n_1146),
.B2(n_1162),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1116),
.A2(n_1132),
.B(n_1092),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1085),
.A2(n_1216),
.B(n_1159),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1074),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1109),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1092),
.A2(n_1159),
.B(n_1198),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1086),
.Y(n_1281)
);

AO21x1_ASAP7_75t_L g1282 ( 
.A1(n_1171),
.A2(n_1112),
.B(n_1184),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1128),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1203),
.A2(n_1118),
.B(n_1131),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_SL g1285 ( 
.A(n_1197),
.B(n_1167),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_L g1286 ( 
.A(n_1175),
.B(n_1148),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1137),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1172),
.B(n_1083),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1169),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1124),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1094),
.A2(n_1195),
.B(n_1099),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1143),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1177),
.A2(n_1178),
.B1(n_1170),
.B2(n_1103),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1069),
.A2(n_1188),
.B(n_1211),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_SL g1295 ( 
.A1(n_1147),
.A2(n_1224),
.B(n_1214),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1213),
.A2(n_1089),
.B(n_1204),
.Y(n_1296)
);

AO32x2_ASAP7_75t_L g1297 ( 
.A1(n_1079),
.A2(n_1183),
.A3(n_1165),
.B1(n_1173),
.B2(n_1115),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1149),
.A2(n_1155),
.B(n_1150),
.Y(n_1298)
);

AOI221x1_ASAP7_75t_L g1299 ( 
.A1(n_1140),
.A2(n_1096),
.B1(n_1168),
.B2(n_1090),
.C(n_1212),
.Y(n_1299)
);

AO32x2_ASAP7_75t_L g1300 ( 
.A1(n_1196),
.A2(n_1194),
.A3(n_1073),
.B1(n_1152),
.B2(n_1121),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1090),
.A2(n_1218),
.B(n_1212),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1111),
.B(n_1141),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1105),
.A2(n_1152),
.B(n_1123),
.C(n_1133),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1196),
.A2(n_1091),
.B(n_1073),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1145),
.A2(n_1152),
.B1(n_1158),
.B2(n_1174),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1218),
.A2(n_1217),
.B(n_1073),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1148),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_SL g1308 ( 
.A(n_1097),
.B(n_1196),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1121),
.A2(n_1148),
.B1(n_1182),
.B2(n_1091),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1182),
.A2(n_1121),
.B(n_1208),
.Y(n_1310)
);

AOI221xp5_ASAP7_75t_L g1311 ( 
.A1(n_1093),
.A2(n_1088),
.B1(n_1084),
.B2(n_891),
.C(n_1082),
.Y(n_1311)
);

AOI221xp5_ASAP7_75t_L g1312 ( 
.A1(n_1182),
.A2(n_1088),
.B1(n_1084),
.B2(n_891),
.C(n_1082),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1186),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1088),
.A2(n_1084),
.B(n_1082),
.C(n_1095),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1191),
.A2(n_896),
.B(n_1070),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1067),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1071),
.B(n_1102),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1066),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1067),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1082),
.A2(n_1117),
.B1(n_1160),
.B2(n_1134),
.C(n_1164),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1200),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1191),
.A2(n_896),
.B(n_1070),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1139),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1066),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1205),
.A2(n_1095),
.A3(n_1207),
.B(n_1186),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1088),
.B(n_712),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1084),
.A2(n_1088),
.B1(n_1082),
.B2(n_392),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1097),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1180),
.B(n_900),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1067),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1088),
.B(n_712),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1169),
.B(n_932),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1100),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1071),
.B(n_1102),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1181),
.B(n_758),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1095),
.C(n_712),
.Y(n_1342)
);

AOI211x1_ASAP7_75t_L g1343 ( 
.A1(n_1088),
.A2(n_1180),
.B(n_1164),
.C(n_1043),
.Y(n_1343)
);

AOI221x1_ASAP7_75t_L g1344 ( 
.A1(n_1084),
.A2(n_1088),
.B1(n_1164),
.B2(n_1206),
.C(n_1095),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1082),
.A2(n_1088),
.B1(n_1180),
.B2(n_1095),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1180),
.B(n_900),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1095),
.C(n_712),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1180),
.B(n_900),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1205),
.A2(n_1095),
.A3(n_1207),
.B(n_1186),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1067),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1088),
.A2(n_674),
.B1(n_712),
.B2(n_1185),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1191),
.A2(n_896),
.B(n_1070),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1191),
.A2(n_896),
.B(n_1070),
.Y(n_1353)
);

AOI221x1_ASAP7_75t_L g1354 ( 
.A1(n_1084),
.A2(n_1088),
.B1(n_1164),
.B2(n_1206),
.C(n_1095),
.Y(n_1354)
);

BUFx10_ASAP7_75t_L g1355 ( 
.A(n_1093),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1169),
.B(n_932),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1180),
.B(n_900),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1200),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1081),
.A2(n_1129),
.B(n_1186),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1181),
.B(n_758),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1088),
.A2(n_1084),
.B(n_1082),
.C(n_1095),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1081),
.A2(n_1129),
.B(n_1186),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1097),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1144),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1067),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_SL g1366 ( 
.A1(n_1164),
.A2(n_1151),
.B(n_1134),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1067),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1205),
.A2(n_1186),
.B(n_1101),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1082),
.A2(n_1088),
.B1(n_1180),
.B2(n_1095),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1174),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1081),
.A2(n_1129),
.B(n_1186),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1180),
.B(n_900),
.Y(n_1372)
);

AO31x2_ASAP7_75t_L g1373 ( 
.A1(n_1205),
.A2(n_1095),
.A3(n_1207),
.B(n_1186),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1084),
.B(n_1088),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1067),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1083),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1144),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1180),
.B(n_928),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1081),
.A2(n_1129),
.B(n_1186),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1081),
.A2(n_1129),
.B(n_1186),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1095),
.A2(n_898),
.B(n_1193),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1075),
.A2(n_717),
.B(n_715),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1191),
.A2(n_896),
.B(n_1070),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1180),
.B(n_900),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1370),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1311),
.A2(n_1374),
.B1(n_1331),
.B2(n_1312),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1261),
.Y(n_1388)
);

INVx8_ASAP7_75t_L g1389 ( 
.A(n_1261),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1329),
.A2(n_1335),
.B1(n_1345),
.B2(n_1369),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1261),
.Y(n_1391)
);

INVx8_ASAP7_75t_L g1392 ( 
.A(n_1322),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1337),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1322),
.Y(n_1394)
);

BUFx4f_ASAP7_75t_SL g1395 ( 
.A(n_1332),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1270),
.A2(n_1285),
.B1(n_1345),
.B2(n_1275),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1377),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1359),
.A2(n_1371),
.B1(n_1381),
.B2(n_1380),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1234),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1275),
.A2(n_1273),
.B1(n_1366),
.B2(n_1308),
.Y(n_1401)
);

OAI22x1_ASAP7_75t_L g1402 ( 
.A1(n_1305),
.A2(n_1268),
.B1(n_1279),
.B2(n_1241),
.Y(n_1402)
);

OAI21xp33_ASAP7_75t_L g1403 ( 
.A1(n_1314),
.A2(n_1361),
.B(n_1264),
.Y(n_1403)
);

AND2x4_ASAP7_75t_SL g1404 ( 
.A(n_1358),
.B(n_1355),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1253),
.A2(n_1354),
.B(n_1344),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1355),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1239),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1363),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1351),
.A2(n_1251),
.B1(n_1340),
.B2(n_1360),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1321),
.A2(n_1259),
.B1(n_1290),
.B2(n_1357),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1377),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1240),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1252),
.Y(n_1413)
);

BUFx2_ASAP7_75t_SL g1414 ( 
.A(n_1358),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1348),
.A2(n_1385),
.B1(n_1372),
.B2(n_1379),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1308),
.A2(n_1362),
.B1(n_1371),
.B2(n_1381),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1359),
.A2(n_1380),
.B1(n_1362),
.B2(n_1282),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1358),
.Y(n_1418)
);

BUFx8_ASAP7_75t_L g1419 ( 
.A(n_1254),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1244),
.A2(n_1291),
.B1(n_1286),
.B2(n_1313),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1237),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1291),
.A2(n_1313),
.B1(n_1295),
.B2(n_1288),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1364),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1258),
.A2(n_1343),
.B1(n_1334),
.B2(n_1350),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1289),
.A2(n_1293),
.B1(n_1378),
.B2(n_1232),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1256),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1321),
.A2(n_1324),
.B1(n_1231),
.B2(n_1283),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1229),
.A2(n_1347),
.B1(n_1342),
.B2(n_1367),
.Y(n_1428)
);

CKINVDCx6p67_ASAP7_75t_R g1429 ( 
.A(n_1336),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1299),
.A2(n_1294),
.B1(n_1320),
.B2(n_1316),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1255),
.A2(n_1292),
.B1(n_1287),
.B2(n_1276),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1278),
.A2(n_1281),
.B1(n_1365),
.B2(n_1375),
.Y(n_1432)
);

CKINVDCx8_ASAP7_75t_R g1433 ( 
.A(n_1356),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1307),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1271),
.A2(n_1272),
.B1(n_1245),
.B2(n_1302),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1267),
.A2(n_1303),
.B(n_1260),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1382),
.A2(n_1245),
.B1(n_1310),
.B2(n_1309),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1243),
.A2(n_1276),
.B1(n_1260),
.B2(n_1309),
.Y(n_1438)
);

XOR2xp5_ASAP7_75t_L g1439 ( 
.A(n_1317),
.B(n_1338),
.Y(n_1439)
);

INVx6_ASAP7_75t_L g1440 ( 
.A(n_1243),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1266),
.A2(n_1280),
.B1(n_1298),
.B2(n_1225),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1301),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1250),
.A2(n_1257),
.B(n_1227),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1243),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1368),
.A2(n_1269),
.B1(n_1296),
.B2(n_1325),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1297),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1368),
.A2(n_1242),
.B1(n_1284),
.B2(n_1265),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1236),
.Y(n_1448)
);

BUFx12f_ASAP7_75t_L g1449 ( 
.A(n_1317),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1306),
.B(n_1349),
.Y(n_1450)
);

NAND2x1p5_ASAP7_75t_L g1451 ( 
.A(n_1236),
.B(n_1318),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1300),
.Y(n_1452)
);

BUFx2_ASAP7_75t_R g1453 ( 
.A(n_1318),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1300),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1242),
.A2(n_1325),
.B1(n_1263),
.B2(n_1277),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1300),
.Y(n_1456)
);

BUFx8_ASAP7_75t_L g1457 ( 
.A(n_1297),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1249),
.A2(n_1274),
.B1(n_1233),
.B2(n_1319),
.Y(n_1458)
);

BUFx4f_ASAP7_75t_SL g1459 ( 
.A(n_1304),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1269),
.A2(n_1262),
.B1(n_1339),
.B2(n_1383),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1225),
.A2(n_1327),
.B1(n_1376),
.B2(n_1330),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1269),
.A2(n_1326),
.B1(n_1341),
.B2(n_1338),
.Y(n_1462)
);

INVx4_ASAP7_75t_L g1463 ( 
.A(n_1246),
.Y(n_1463)
);

OAI21xp33_ASAP7_75t_L g1464 ( 
.A1(n_1226),
.A2(n_1248),
.B(n_1247),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1328),
.A2(n_1349),
.B(n_1373),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1235),
.A2(n_1230),
.B1(n_1384),
.B2(n_1315),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1238),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1349),
.B(n_1238),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_1323),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1352),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1238),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1353),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1332),
.Y(n_1473)
);

INVx6_ASAP7_75t_L g1474 ( 
.A(n_1261),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1228),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1270),
.A2(n_674),
.B1(n_1088),
.B2(n_820),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1332),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1261),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1483)
);

INVx5_ASAP7_75t_L g1484 ( 
.A(n_1261),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1228),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1487)
);

INVx8_ASAP7_75t_L g1488 ( 
.A(n_1261),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1261),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1228),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1228),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1332),
.Y(n_1493)
);

AOI21xp33_ASAP7_75t_L g1494 ( 
.A1(n_1342),
.A2(n_1088),
.B(n_1082),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1253),
.A2(n_1088),
.B1(n_1082),
.B2(n_820),
.Y(n_1496)
);

AOI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1342),
.A2(n_1088),
.B(n_1082),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1228),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1332),
.Y(n_1500)
);

CKINVDCx6p67_ASAP7_75t_R g1501 ( 
.A(n_1237),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1253),
.A2(n_1088),
.B1(n_1082),
.B2(n_820),
.Y(n_1503)
);

INVx3_ASAP7_75t_SL g1504 ( 
.A(n_1337),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1370),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1331),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1332),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1311),
.A2(n_1084),
.B1(n_1088),
.B2(n_1082),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1329),
.A2(n_1082),
.B(n_1084),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1253),
.A2(n_1088),
.B1(n_1082),
.B2(n_1331),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1261),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1270),
.A2(n_674),
.B1(n_1088),
.B2(n_820),
.Y(n_1513)
);

CKINVDCx16_ASAP7_75t_R g1514 ( 
.A(n_1355),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1261),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1228),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1254),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1450),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1465),
.B(n_1468),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1466),
.A2(n_1458),
.B(n_1455),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1397),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1398),
.B(n_1476),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1400),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1407),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1442),
.B(n_1399),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1397),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1413),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1416),
.B(n_1452),
.Y(n_1528)
);

AND2x4_ASAP7_75t_SL g1529 ( 
.A(n_1429),
.B(n_1423),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1454),
.B(n_1456),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1426),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1471),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1411),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1412),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1443),
.A2(n_1460),
.B(n_1403),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1424),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1443),
.B(n_1460),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1390),
.B(n_1417),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1411),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1424),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1467),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1419),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1472),
.B(n_1441),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1432),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1434),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1469),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1457),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1447),
.A2(n_1462),
.B(n_1464),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1440),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_1393),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1440),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1470),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1432),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1406),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1492),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1431),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1507),
.A2(n_1511),
.B1(n_1496),
.B2(n_1503),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1444),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_SL g1559 ( 
.A(n_1419),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1430),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1438),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1510),
.A2(n_1387),
.B1(n_1481),
.B2(n_1479),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1434),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1461),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1461),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1464),
.A2(n_1437),
.B(n_1420),
.Y(n_1566)
);

OR2x6_ASAP7_75t_L g1567 ( 
.A(n_1436),
.B(n_1405),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1499),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1422),
.A2(n_1436),
.B(n_1428),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1463),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1463),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1410),
.Y(n_1572)
);

AOI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1496),
.A2(n_1402),
.B(n_1415),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1517),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1410),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1427),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1449),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1445),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1451),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1457),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1405),
.B(n_1510),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1427),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1475),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1485),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1487),
.B(n_1495),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1415),
.B(n_1478),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1491),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1451),
.A2(n_1489),
.B(n_1498),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1459),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1396),
.B(n_1446),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1483),
.B(n_1505),
.Y(n_1591)
);

BUFx2_ASAP7_75t_SL g1592 ( 
.A(n_1448),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1423),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1401),
.B(n_1509),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1486),
.A2(n_1502),
.B(n_1439),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1516),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1494),
.A2(n_1497),
.B(n_1409),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1477),
.A2(n_1513),
.B1(n_1433),
.B2(n_1425),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1484),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1484),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1435),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1484),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1453),
.B(n_1482),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1408),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1391),
.Y(n_1605)
);

BUFx2_ASAP7_75t_SL g1606 ( 
.A(n_1394),
.Y(n_1606)
);

OA21x2_ASAP7_75t_L g1607 ( 
.A1(n_1473),
.A2(n_1480),
.B(n_1493),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1421),
.A2(n_1501),
.B1(n_1418),
.B2(n_1508),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1389),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1389),
.B(n_1392),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1514),
.A2(n_1500),
.B1(n_1395),
.B2(n_1506),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1414),
.B(n_1504),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1392),
.B(n_1488),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1404),
.B(n_1386),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1388),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1388),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1474),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1392),
.B(n_1488),
.Y(n_1618)
);

INVx5_ASAP7_75t_SL g1619 ( 
.A(n_1558),
.Y(n_1619)
);

BUFx8_ASAP7_75t_SL g1620 ( 
.A(n_1550),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1562),
.A2(n_1474),
.B1(n_1490),
.B2(n_1512),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1522),
.B(n_1515),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1535),
.A2(n_1512),
.B(n_1515),
.C(n_1594),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1557),
.A2(n_1594),
.B1(n_1591),
.B2(n_1581),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1569),
.A2(n_1595),
.B(n_1586),
.C(n_1588),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1534),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_SL g1627 ( 
.A(n_1554),
.B(n_1598),
.C(n_1614),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1607),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_SL g1629 ( 
.A1(n_1586),
.A2(n_1572),
.B(n_1575),
.C(n_1576),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1585),
.B(n_1521),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1577),
.Y(n_1631)
);

INVx5_ASAP7_75t_L g1632 ( 
.A(n_1537),
.Y(n_1632)
);

OAI211xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1560),
.A2(n_1561),
.B(n_1604),
.C(n_1564),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1525),
.B(n_1518),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1537),
.A2(n_1565),
.B(n_1564),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1581),
.A2(n_1538),
.B1(n_1567),
.B2(n_1597),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1533),
.B(n_1539),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1525),
.B(n_1541),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1567),
.B(n_1528),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1581),
.A2(n_1567),
.B1(n_1590),
.B2(n_1575),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1560),
.A2(n_1561),
.B1(n_1565),
.B2(n_1544),
.C(n_1572),
.Y(n_1641)
);

INVx4_ASAP7_75t_L g1642 ( 
.A(n_1577),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1574),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_SL g1644 ( 
.A(n_1554),
.B(n_1589),
.Y(n_1644)
);

AO32x2_ASAP7_75t_L g1645 ( 
.A1(n_1551),
.A2(n_1593),
.A3(n_1530),
.B1(n_1602),
.B2(n_1599),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1553),
.B(n_1519),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1569),
.A2(n_1588),
.B(n_1597),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1519),
.B(n_1579),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1545),
.B(n_1563),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1597),
.A2(n_1589),
.B1(n_1590),
.B2(n_1582),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1537),
.A2(n_1589),
.B1(n_1559),
.B2(n_1580),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1526),
.B(n_1584),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1597),
.A2(n_1573),
.B(n_1566),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1601),
.B(n_1556),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1547),
.B(n_1580),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1577),
.Y(n_1657)
);

AO21x2_ASAP7_75t_L g1658 ( 
.A1(n_1570),
.A2(n_1571),
.B(n_1548),
.Y(n_1658)
);

AO21x2_ASAP7_75t_L g1659 ( 
.A1(n_1548),
.A2(n_1520),
.B(n_1566),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1536),
.A2(n_1540),
.B(n_1556),
.C(n_1537),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_SL g1661 ( 
.A(n_1613),
.B(n_1617),
.C(n_1616),
.Y(n_1661)
);

AO21x2_ASAP7_75t_L g1662 ( 
.A1(n_1520),
.A2(n_1552),
.B(n_1546),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1536),
.A2(n_1540),
.B(n_1532),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1543),
.A2(n_1608),
.B(n_1611),
.Y(n_1664)
);

NAND2xp33_ASAP7_75t_R g1665 ( 
.A(n_1549),
.B(n_1578),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1578),
.A2(n_1549),
.B(n_1603),
.C(n_1529),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1524),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1624),
.A2(n_1558),
.B1(n_1592),
.B2(n_1542),
.Y(n_1668)
);

OAI22x1_ASAP7_75t_SL g1669 ( 
.A1(n_1642),
.A2(n_1551),
.B1(n_1593),
.B2(n_1609),
.Y(n_1669)
);

AND2x4_ASAP7_75t_SL g1670 ( 
.A(n_1661),
.B(n_1638),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1638),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1626),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1659),
.B(n_1543),
.Y(n_1673)
);

CKINVDCx14_ASAP7_75t_R g1674 ( 
.A(n_1655),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1645),
.B(n_1543),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1633),
.B(n_1605),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1645),
.B(n_1527),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1645),
.B(n_1531),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1555),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1628),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1636),
.A2(n_1558),
.B1(n_1592),
.B2(n_1542),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1663),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1663),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1643),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1667),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1648),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1653),
.B(n_1596),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1647),
.B(n_1596),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1667),
.B(n_1649),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1640),
.A2(n_1641),
.B1(n_1633),
.B2(n_1664),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1646),
.B(n_1654),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1662),
.B(n_1587),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1632),
.A2(n_1558),
.B1(n_1603),
.B2(n_1583),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1680),
.Y(n_1695)
);

AND3x1_ASAP7_75t_L g1696 ( 
.A(n_1691),
.B(n_1627),
.C(n_1644),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1681),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1681),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1658),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1683),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1675),
.B(n_1634),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1662),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1680),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1675),
.B(n_1634),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1683),
.Y(n_1705)
);

AOI31xp33_ASAP7_75t_L g1706 ( 
.A1(n_1691),
.A2(n_1665),
.A3(n_1651),
.B(n_1650),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1686),
.B(n_1635),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1684),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1686),
.B(n_1635),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1668),
.A2(n_1632),
.B1(n_1558),
.B2(n_1665),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1670),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1668),
.A2(n_1625),
.B(n_1623),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1688),
.B(n_1637),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1672),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1677),
.Y(n_1715)
);

AOI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1682),
.A2(n_1627),
.B1(n_1625),
.B2(n_1654),
.C(n_1629),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1677),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1672),
.Y(n_1718)
);

BUFx2_ASAP7_75t_SL g1719 ( 
.A(n_1677),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1688),
.B(n_1656),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1677),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1674),
.Y(n_1722)
);

OAI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1682),
.A2(n_1623),
.B(n_1629),
.C(n_1660),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1679),
.B(n_1648),
.Y(n_1724)
);

AOI21xp33_ASAP7_75t_L g1725 ( 
.A1(n_1676),
.A2(n_1630),
.B(n_1622),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1700),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1714),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1714),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1701),
.B(n_1674),
.Y(n_1729)
);

NAND2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1702),
.B(n_1632),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1725),
.B(n_1692),
.Y(n_1731)
);

NAND2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1702),
.B(n_1632),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1711),
.B(n_1671),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1725),
.B(n_1692),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1714),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1718),
.Y(n_1736)
);

OR2x6_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1660),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1713),
.B(n_1685),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1718),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1718),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1713),
.B(n_1690),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1705),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1707),
.B(n_1690),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1711),
.B(n_1671),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1701),
.B(n_1687),
.Y(n_1746)
);

AND2x4_ASAP7_75t_SL g1747 ( 
.A(n_1711),
.B(n_1661),
.Y(n_1747)
);

NAND2x1_ASAP7_75t_L g1748 ( 
.A(n_1702),
.B(n_1679),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1707),
.B(n_1693),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1695),
.Y(n_1750)
);

NAND2x1_ASAP7_75t_L g1751 ( 
.A(n_1711),
.B(n_1678),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1695),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1701),
.B(n_1687),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1709),
.B(n_1693),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1701),
.B(n_1687),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1722),
.B(n_1620),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1705),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1708),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1709),
.B(n_1689),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1708),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1720),
.B(n_1689),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1700),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1739),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1748),
.A2(n_1706),
.B(n_1712),
.C(n_1716),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1729),
.B(n_1719),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1729),
.B(n_1719),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1744),
.B(n_1703),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1739),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1726),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1740),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1740),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1742),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1742),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1733),
.B(n_1719),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1743),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1756),
.B(n_1620),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1743),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1731),
.B(n_1722),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1733),
.B(n_1704),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1734),
.B(n_1741),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1751),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1733),
.B(n_1715),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1745),
.B(n_1746),
.Y(n_1784)
);

OAI32xp33_ASAP7_75t_L g1785 ( 
.A1(n_1730),
.A2(n_1717),
.A3(n_1721),
.B1(n_1696),
.B2(n_1699),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1745),
.B(n_1715),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1757),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1745),
.B(n_1717),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1757),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1759),
.B(n_1697),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1746),
.B(n_1721),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1758),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1749),
.B(n_1697),
.Y(n_1793)
);

NAND2x1_ASAP7_75t_L g1794 ( 
.A(n_1737),
.B(n_1711),
.Y(n_1794)
);

NOR5xp2_ASAP7_75t_L g1795 ( 
.A(n_1750),
.B(n_1706),
.C(n_1710),
.D(n_1723),
.E(n_1712),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1758),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1752),
.B(n_1703),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1727),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1760),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1762),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1760),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1762),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1728),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1735),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1736),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1765),
.B(n_1737),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1798),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1765),
.B(n_1766),
.Y(n_1808)
);

NOR2xp67_ASAP7_75t_L g1809 ( 
.A(n_1782),
.B(n_1711),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1798),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1803),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1766),
.B(n_1737),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1781),
.A2(n_1737),
.B1(n_1716),
.B2(n_1710),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1788),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1780),
.B(n_1747),
.Y(n_1816)
);

INVx8_ASAP7_75t_L g1817 ( 
.A(n_1774),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1794),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1764),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1779),
.B(n_1738),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1788),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1780),
.B(n_1755),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1785),
.A2(n_1748),
.B(n_1723),
.C(n_1730),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1767),
.B(n_1749),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1763),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1774),
.B(n_1755),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1794),
.Y(n_1828)
);

AOI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1785),
.A2(n_1754),
.B(n_1696),
.C(n_1699),
.Y(n_1829)
);

NAND3xp33_ASAP7_75t_L g1830 ( 
.A(n_1795),
.B(n_1754),
.C(n_1676),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1767),
.B(n_1761),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1763),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1697),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1776),
.B(n_1612),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1768),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1797),
.B(n_1698),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1783),
.B(n_1724),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_R g1838 ( 
.A(n_1795),
.B(n_1577),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1782),
.B(n_1747),
.Y(n_1839)
);

OR2x6_ASAP7_75t_L g1840 ( 
.A(n_1783),
.B(n_1730),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1768),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1803),
.B(n_1805),
.C(n_1804),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1819),
.B(n_1732),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1808),
.B(n_1806),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1811),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1813),
.A2(n_1830),
.B1(n_1829),
.B2(n_1819),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1826),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1807),
.Y(n_1848)
);

OA22x2_ASAP7_75t_L g1849 ( 
.A1(n_1818),
.A2(n_1786),
.B1(n_1751),
.B2(n_1805),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1820),
.B(n_1786),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1834),
.B(n_1817),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1838),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1826),
.Y(n_1853)
);

OAI32xp33_ASAP7_75t_L g1854 ( 
.A1(n_1806),
.A2(n_1732),
.A3(n_1782),
.B1(n_1793),
.B2(n_1790),
.Y(n_1854)
);

CKINVDCx14_ASAP7_75t_R g1855 ( 
.A(n_1812),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1832),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1808),
.B(n_1812),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1824),
.A2(n_1732),
.B(n_1782),
.Y(n_1858)
);

OAI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1825),
.A2(n_1790),
.B(n_1793),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1817),
.A2(n_1670),
.B1(n_1673),
.B2(n_1639),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1817),
.A2(n_1804),
.B(n_1771),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1815),
.B(n_1791),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1815),
.B(n_1791),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1832),
.Y(n_1864)
);

OAI322xp33_ASAP7_75t_L g1865 ( 
.A1(n_1807),
.A2(n_1787),
.A3(n_1777),
.B1(n_1775),
.B2(n_1773),
.C1(n_1772),
.C2(n_1771),
.Y(n_1865)
);

NOR2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1821),
.B(n_1577),
.Y(n_1866)
);

OAI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1840),
.A2(n_1694),
.B1(n_1801),
.B2(n_1775),
.C(n_1799),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1827),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1848),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1848),
.Y(n_1870)
);

NOR2x1_ASAP7_75t_L g1871 ( 
.A(n_1846),
.B(n_1810),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1847),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1855),
.B(n_1851),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1855),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1865),
.A2(n_1842),
.B1(n_1810),
.B2(n_1821),
.C(n_1817),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1857),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1853),
.Y(n_1877)
);

INVx2_ASAP7_75t_SL g1878 ( 
.A(n_1857),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1852),
.A2(n_1816),
.B1(n_1839),
.B2(n_1840),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1856),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1868),
.B(n_1831),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1844),
.B(n_1814),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1868),
.B(n_1828),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1864),
.Y(n_1884)
);

NOR4xp25_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1841),
.C(n_1835),
.D(n_1828),
.Y(n_1885)
);

AOI21xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1851),
.A2(n_1849),
.B(n_1854),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1862),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1858),
.A2(n_1861),
.B(n_1843),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_SL g1889 ( 
.A(n_1874),
.B(n_1839),
.Y(n_1889)
);

AOI221x1_ASAP7_75t_SL g1890 ( 
.A1(n_1887),
.A2(n_1859),
.B1(n_1863),
.B2(n_1850),
.C(n_1835),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1871),
.B(n_1849),
.Y(n_1891)
);

OAI21xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1875),
.A2(n_1860),
.B(n_1816),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1883),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1878),
.B(n_1816),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1883),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1876),
.B(n_1866),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1869),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1882),
.B(n_1814),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1873),
.B(n_1867),
.Y(n_1899)
);

NAND4xp25_ASAP7_75t_L g1900 ( 
.A(n_1889),
.B(n_1879),
.C(n_1888),
.D(n_1886),
.Y(n_1900)
);

NOR3xp33_ASAP7_75t_L g1901 ( 
.A(n_1899),
.B(n_1888),
.C(n_1870),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1893),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1895),
.B(n_1885),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_L g1904 ( 
.A(n_1899),
.B(n_1877),
.C(n_1872),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1891),
.A2(n_1885),
.B(n_1881),
.Y(n_1905)
);

AOI222xp33_ASAP7_75t_L g1906 ( 
.A1(n_1891),
.A2(n_1884),
.B1(n_1880),
.B2(n_1841),
.C1(n_1839),
.C2(n_1809),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1892),
.B(n_1621),
.C(n_1833),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1890),
.B(n_1822),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_L g1909 ( 
.A(n_1894),
.B(n_1827),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1897),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1905),
.A2(n_1900),
.B(n_1903),
.Y(n_1911)
);

O2A1O1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1901),
.A2(n_1896),
.B(n_1898),
.C(n_1840),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_L g1913 ( 
.A(n_1906),
.B(n_1840),
.C(n_1836),
.Y(n_1913)
);

AOI211xp5_ASAP7_75t_L g1914 ( 
.A1(n_1904),
.A2(n_1836),
.B(n_1833),
.C(n_1822),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1902),
.B(n_1837),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1908),
.B(n_1823),
.Y(n_1916)
);

OAI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1911),
.A2(n_1907),
.B1(n_1909),
.B2(n_1910),
.C(n_1694),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_L g1918 ( 
.A(n_1912),
.B(n_1916),
.C(n_1913),
.Y(n_1918)
);

AOI211xp5_ASAP7_75t_SL g1919 ( 
.A1(n_1915),
.A2(n_1618),
.B(n_1823),
.C(n_1617),
.Y(n_1919)
);

NAND4xp25_ASAP7_75t_L g1920 ( 
.A(n_1914),
.B(n_1666),
.C(n_1618),
.D(n_1642),
.Y(n_1920)
);

NAND3xp33_ASAP7_75t_SL g1921 ( 
.A(n_1911),
.B(n_1666),
.C(n_1619),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1911),
.A2(n_1619),
.B1(n_1801),
.B2(n_1770),
.Y(n_1922)
);

AO22x1_ASAP7_75t_L g1923 ( 
.A1(n_1918),
.A2(n_1787),
.B1(n_1792),
.B2(n_1799),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1919),
.Y(n_1924)
);

NOR4xp75_ASAP7_75t_L g1925 ( 
.A(n_1917),
.B(n_1609),
.C(n_1652),
.D(n_1599),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1922),
.B(n_1770),
.Y(n_1926)
);

NOR2x1_ASAP7_75t_L g1927 ( 
.A(n_1921),
.B(n_1772),
.Y(n_1927)
);

AOI22x1_ASAP7_75t_L g1928 ( 
.A1(n_1924),
.A2(n_1920),
.B1(n_1802),
.B2(n_1800),
.Y(n_1928)
);

NOR3xp33_ASAP7_75t_L g1929 ( 
.A(n_1923),
.B(n_1616),
.C(n_1615),
.Y(n_1929)
);

NAND3xp33_ASAP7_75t_SL g1930 ( 
.A(n_1925),
.B(n_1619),
.C(n_1615),
.Y(n_1930)
);

OAI22x1_ASAP7_75t_L g1931 ( 
.A1(n_1928),
.A2(n_1927),
.B1(n_1926),
.B2(n_1777),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1931),
.A2(n_1930),
.B1(n_1929),
.B2(n_1610),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1932),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1932),
.A2(n_1802),
.B1(n_1800),
.B2(n_1769),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1933),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1934),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1935),
.Y(n_1937)
);

OAI21xp33_ASAP7_75t_L g1938 ( 
.A1(n_1937),
.A2(n_1936),
.B(n_1778),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1938),
.A2(n_1802),
.B1(n_1800),
.B2(n_1769),
.Y(n_1939)
);

AOI22x1_ASAP7_75t_L g1940 ( 
.A1(n_1939),
.A2(n_1606),
.B1(n_1600),
.B2(n_1602),
.Y(n_1940)
);

AOI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1940),
.A2(n_1796),
.B1(n_1792),
.B2(n_1773),
.C(n_1789),
.Y(n_1941)
);

AOI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1941),
.A2(n_1631),
.B(n_1657),
.C(n_1600),
.Y(n_1942)
);


endmodule