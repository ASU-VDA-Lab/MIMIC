module fake_jpeg_29402_n_156 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_156);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_30),
.Y(n_54)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_30),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_29),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_64),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_2),
.B(n_5),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_68),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_31),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_14),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_32),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_25),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_72),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_26),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_77),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_58),
.B(n_51),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_78),
.B1(n_84),
.B2(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_46),
.B1(n_53),
.B2(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_21),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_23),
.B1(n_19),
.B2(n_24),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_62),
.B1(n_59),
.B2(n_2),
.Y(n_95)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_23),
.B1(n_19),
.B2(n_30),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_12),
.Y(n_99)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_57),
.B1(n_62),
.B2(n_60),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_73),
.B1(n_77),
.B2(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_12),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_59),
.B(n_60),
.C(n_5),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_6),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_60),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_6),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_106),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_90),
.B1(n_94),
.B2(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_86),
.B1(n_59),
.B2(n_76),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_119),
.B(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_91),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_92),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_71),
.C(n_70),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_120),
.C(n_92),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_71),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_118),
.C(n_120),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_94),
.B(n_95),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_127),
.A2(n_122),
.B(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_128),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_117),
.B(n_115),
.C(n_107),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_103),
.C(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_129),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_140),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_108),
.A3(n_111),
.B1(n_125),
.B2(n_119),
.C1(n_112),
.C2(n_83),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_131),
.B(n_134),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_144),
.B(n_138),
.Y(n_146)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_91),
.Y(n_151)
);

AOI21x1_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_119),
.B(n_97),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_148),
.Y(n_149)
);

OAI21x1_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_97),
.B(n_10),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_139),
.C(n_143),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_151),
.B(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_153),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_7),
.C(n_13),
.Y(n_156)
);


endmodule