module real_jpeg_12131_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx4_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_52),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_2),
.A2(n_52),
.B1(n_62),
.B2(n_64),
.Y(n_168)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_5),
.A2(n_62),
.B1(n_64),
.B2(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_5),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_6),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_7),
.B(n_36),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_60),
.C(n_62),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_7),
.A2(n_27),
.B1(n_48),
.B2(n_50),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_7),
.A2(n_77),
.B1(n_113),
.B2(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_7),
.B(n_102),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_54),
.B1(n_62),
.B2(n_64),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_12),
.A2(n_38),
.B1(n_48),
.B2(n_50),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_12),
.A2(n_38),
.B1(n_62),
.B2(n_64),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_13),
.A2(n_62),
.B1(n_64),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_13),
.A2(n_48),
.B1(n_50),
.B2(n_80),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_14),
.A2(n_62),
.B1(n_64),
.B2(n_69),
.Y(n_95)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_96),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_96),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_86),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_21),
.B(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_22),
.B(n_40),
.C(n_70),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_23),
.A2(n_31),
.B(n_35),
.C(n_85),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_27),
.CON(n_23),
.SN(n_23)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_24),
.B(n_32),
.C(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_27),
.B(n_35),
.CON(n_135),
.SN(n_135)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_27),
.B(n_77),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_27),
.B(n_118),
.Y(n_178)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_29),
.A2(n_33),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_35),
.B(n_46),
.C(n_50),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_37),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_55),
.B2(n_70),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_51),
.B2(n_53),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_47),
.B1(n_51),
.B2(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_42),
.A2(n_53),
.B(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_43),
.A2(n_89),
.B1(n_102),
.B2(n_135),
.Y(n_137)
);

AND2x4_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_45),
.A2(n_48),
.B(n_135),
.C(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_50),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_48),
.B(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_65),
.B(n_67),
.Y(n_55)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_56),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_56),
.A2(n_118),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_56),
.A2(n_118),
.B1(n_140),
.B2(n_165),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_SL g60 ( 
.A(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_61),
.A2(n_121),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_61),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_64),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_71),
.A2(n_72),
.B1(n_86),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_83),
.B2(n_84),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_81),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_75),
.A2(n_116),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_75),
.A2(n_76),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_76),
.B(n_132),
.Y(n_191)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_79),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_95),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_77),
.A2(n_113),
.B1(n_168),
.B2(n_176),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.C(n_92),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_87),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_109),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_107),
.B2(n_108),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B(n_115),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_113),
.A2(n_170),
.B(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_200),
.B(n_205),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_154),
.B(n_199),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_142),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_142),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.C(n_138),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_128),
.A2(n_129),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_137),
.B(n_138),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_143),
.B(n_148),
.C(n_152),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_193),
.B(n_198),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_182),
.B(n_192),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_171),
.B(n_181),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_166),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_180),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_189),
.C(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_197),
.Y(n_198)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_204),
.Y(n_205)
);


endmodule