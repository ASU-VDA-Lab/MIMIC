module fake_jpeg_26459_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_54),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_26),
.Y(n_88)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_39),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_30),
.B1(n_17),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_22),
.B1(n_16),
.B2(n_31),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_20),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_62),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_30),
.B1(n_22),
.B2(n_17),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_73),
.B(n_25),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_30),
.B1(n_33),
.B2(n_16),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_72),
.B(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_81),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_22),
.B1(n_31),
.B2(n_33),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_16),
.B(n_33),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_79),
.B1(n_82),
.B2(n_32),
.Y(n_120)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_61),
.B1(n_43),
.B2(n_51),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_23),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_58),
.B1(n_43),
.B2(n_51),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_88),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_32),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_50),
.C(n_46),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_60),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g96 ( 
.A(n_92),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_67),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_108),
.C(n_122),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_100),
.Y(n_140)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_87),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_55),
.C(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_52),
.B1(n_26),
.B2(n_21),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_118),
.B1(n_78),
.B2(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_21),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_28),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_26),
.B(n_21),
.C(n_20),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_117),
.B(n_93),
.C(n_86),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_28),
.B1(n_27),
.B2(n_29),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_46),
.A3(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_78),
.B1(n_91),
.B2(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_29),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_46),
.C(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_128),
.B1(n_144),
.B2(n_111),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_77),
.C(n_90),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_105),
.C(n_100),
.Y(n_177)
);

OR2x4_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_90),
.Y(n_135)
);

OR2x4_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_93),
.B1(n_62),
.B2(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_86),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_145),
.Y(n_162)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_150),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_19),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_127),
.Y(n_183)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_64),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_64),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_153),
.A2(n_159),
.B(n_176),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_168),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_117),
.B1(n_120),
.B2(n_98),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_170),
.B1(n_178),
.B2(n_132),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_117),
.B1(n_102),
.B2(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_96),
.C(n_104),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_12),
.C(n_11),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_184),
.B1(n_19),
.B2(n_1),
.Y(n_201)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_174),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_132),
.B(n_94),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_10),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_110),
.B(n_116),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_123),
.C(n_24),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_107),
.B1(n_27),
.B2(n_24),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_64),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_181),
.B(n_0),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_24),
.B1(n_19),
.B2(n_2),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_24),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_144),
.B(n_146),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_186),
.A2(n_190),
.B(n_201),
.Y(n_234)
);

OAI22x1_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_137),
.B1(n_128),
.B2(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_127),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_195),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_133),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_125),
.B1(n_137),
.B2(n_136),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_168),
.B1(n_169),
.B2(n_181),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_19),
.C(n_8),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_14),
.C(n_13),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_14),
.C(n_13),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_184),
.C(n_183),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_162),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_12),
.C(n_11),
.Y(n_209)
);

NOR4xp25_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_179),
.C(n_162),
.D(n_160),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_182),
.B(n_163),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_10),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_213),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_217),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_226),
.B1(n_229),
.B2(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_227),
.B1(n_231),
.B2(n_233),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_186),
.A2(n_173),
.B1(n_155),
.B2(n_176),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_158),
.B1(n_154),
.B2(n_174),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_157),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_155),
.B1(n_160),
.B2(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_203),
.B(n_201),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_195),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_242),
.B1(n_246),
.B2(n_252),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_187),
.B1(n_191),
.B2(n_189),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_194),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_199),
.C(n_191),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_248),
.C(n_250),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_218),
.B1(n_231),
.B2(n_226),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_213),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_200),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_192),
.B1(n_196),
.B2(n_154),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_216),
.B1(n_233),
.B2(n_214),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_203),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_214),
.B1(n_234),
.B2(n_219),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_223),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_223),
.C(n_235),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_10),
.C(n_9),
.Y(n_275)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_215),
.B1(n_202),
.B2(n_234),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_245),
.B1(n_240),
.B2(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_196),
.B1(n_156),
.B2(n_174),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_247),
.A3(n_248),
.B1(n_250),
.B2(n_242),
.C1(n_244),
.C2(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_278),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_280),
.C(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_282),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_9),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_8),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_8),
.C(n_1),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_259),
.B(n_260),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_0),
.B(n_1),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_256),
.B1(n_257),
.B2(n_269),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_293),
.B(n_3),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_2),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_291),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_3),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_280),
.A2(n_3),
.B(n_4),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_291),
.B(n_284),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_301),
.B(n_281),
.Y(n_304)
);

A2O1A1O1Ixp25_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_287),
.B(n_282),
.C(n_277),
.D(n_7),
.Y(n_306)
);

OAI21x1_ASAP7_75t_SL g308 ( 
.A1(n_306),
.A2(n_302),
.B(n_299),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_305),
.B(n_300),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_307),
.B(n_5),
.Y(n_310)
);

AOI321xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_298),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_6),
.Y(n_312)
);


endmodule