module fake_ariane_1331_n_1816 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1816);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1816;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1777;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_24),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_4),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_21),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_29),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_64),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_31),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_98),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_106),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_76),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_8),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_32),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_45),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_45),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_10),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_125),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_74),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_24),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_150),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_129),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_18),
.Y(n_203)
);

BUFx8_ASAP7_75t_SL g204 ( 
.A(n_79),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_142),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_17),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_40),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_83),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_99),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_58),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_139),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_130),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_126),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_157),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_90),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_40),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_31),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_131),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_46),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_60),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_73),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_22),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_109),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_141),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_119),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_152),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_116),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_55),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_65),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_75),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_56),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_61),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_1),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_161),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_121),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_68),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_87),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_92),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_28),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_164),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_103),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_166),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_117),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_28),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_38),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_59),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_14),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_96),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_93),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_16),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_26),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_22),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_67),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_15),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_77),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_50),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_110),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_39),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_69),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_132),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_5),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_25),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_88),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_23),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_94),
.Y(n_280)
);

INVxp33_ASAP7_75t_R g281 ( 
.A(n_18),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_120),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_124),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_84),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_30),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_26),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_6),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_33),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_55),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_159),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_135),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_71),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_163),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_160),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_19),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_72),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_100),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_151),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_57),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_162),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_34),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_5),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_105),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_80),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_108),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_36),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_3),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_56),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_70),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_107),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_97),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_43),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_155),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_113),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_9),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_81),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_53),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_44),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_15),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_11),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_4),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_7),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_43),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_102),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_12),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_123),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_62),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_167),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_20),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_138),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_37),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_95),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_51),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_33),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_154),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_53),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_57),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_16),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_221),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_221),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_204),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_334),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_195),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_203),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_286),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_198),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_221),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_211),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_214),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_245),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_246),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_170),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_251),
.B(n_0),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_221),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_173),
.B(n_0),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_221),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_212),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_271),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_175),
.B(n_2),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_271),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_215),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_200),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_203),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_271),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_271),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_284),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_284),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_R g372 ( 
.A(n_189),
.B(n_111),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_259),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_282),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_259),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_206),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_284),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_251),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_284),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_284),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_176),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_176),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_208),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_226),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_229),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_243),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_288),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_181),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_279),
.B(n_6),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_309),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_279),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_249),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_273),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_253),
.Y(n_394)
);

BUFx10_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_181),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_258),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_316),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_260),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_273),
.B(n_7),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_262),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_338),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_194),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_194),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_265),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_180),
.B(n_9),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_196),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_R g408 ( 
.A(n_304),
.B(n_114),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_209),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_209),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_187),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_196),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_315),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_209),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_266),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_227),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_227),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_227),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_267),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_218),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_315),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_269),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_170),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_219),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_236),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_218),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_252),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_341),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_359),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_201),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_368),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_388),
.B(n_396),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_L g450 ( 
.A(n_372),
.B(n_192),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_370),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_256),
.C(n_239),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_356),
.A2(n_362),
.B(n_403),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_396),
.B(n_403),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_404),
.B(n_202),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_345),
.B(n_306),
.Y(n_462)
);

BUFx8_ASAP7_75t_L g463 ( 
.A(n_404),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_240),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_367),
.B(n_252),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_412),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_373),
.B(n_287),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_375),
.B(n_289),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_421),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_381),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_SL g481 ( 
.A(n_408),
.B(n_171),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_391),
.B(n_300),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_382),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_172),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_344),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_411),
.B(n_303),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_393),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_425),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_425),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_378),
.B(n_395),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_395),
.B(n_207),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_395),
.B(n_223),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_358),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_354),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_374),
.B(n_313),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_364),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_365),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_420),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_501),
.B(n_374),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_462),
.B(n_384),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_433),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_385),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

BUFx6f_ASAP7_75t_SL g514 ( 
.A(n_501),
.Y(n_514)
);

OA22x2_ASAP7_75t_L g515 ( 
.A1(n_487),
.A2(n_343),
.B1(n_321),
.B2(n_330),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_240),
.Y(n_518)
);

OAI22x1_ASAP7_75t_L g519 ( 
.A1(n_430),
.A2(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_472),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_430),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_472),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_426),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_490),
.B(n_386),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_501),
.B(n_392),
.Y(n_526)
);

NOR2x1p5_ASAP7_75t_L g527 ( 
.A(n_496),
.B(n_342),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_462),
.B(n_394),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_501),
.B(n_397),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_453),
.A2(n_346),
.B1(n_427),
.B2(n_326),
.Y(n_530)
);

CKINVDCx11_ASAP7_75t_R g531 ( 
.A(n_486),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_324),
.Y(n_532)
);

BUFx4f_ASAP7_75t_L g533 ( 
.A(n_501),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_501),
.B(n_399),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_502),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_472),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_487),
.B(n_462),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_490),
.B(n_401),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_438),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_501),
.B(n_405),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_443),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_463),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_492),
.B(n_415),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_493),
.B(n_419),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_442),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_453),
.A2(n_414),
.B1(n_418),
.B2(n_417),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_462),
.B(n_422),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_462),
.B(n_274),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_466),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_472),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_463),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_442),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_472),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_443),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_442),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_498),
.B(n_178),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_493),
.B(n_409),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_444),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_444),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_498),
.B(n_410),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_503),
.B(n_178),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_446),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_446),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_492),
.B(n_470),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_449),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_466),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_472),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_447),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_503),
.B(n_496),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_503),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_470),
.B(n_171),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_502),
.B(n_308),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_487),
.A2(n_416),
.B1(n_323),
.B2(n_337),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_463),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_491),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_496),
.A2(n_191),
.B1(n_174),
.B2(n_177),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_503),
.B(n_179),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_466),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_463),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_449),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_451),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_449),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_470),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_487),
.B(n_473),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_486),
.B(n_174),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_503),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g595 ( 
.A(n_504),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_496),
.B(n_349),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_495),
.B(n_179),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_496),
.B(n_352),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_449),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_503),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_458),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_449),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_481),
.A2(n_290),
.B1(n_339),
.B2(n_302),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_448),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_454),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_458),
.Y(n_606)
);

AOI22x1_ASAP7_75t_L g607 ( 
.A1(n_491),
.A2(n_191),
.B1(n_318),
.B2(n_335),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_466),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_448),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_503),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_448),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_460),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_183),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_494),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_504),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_473),
.B(n_177),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_454),
.Y(n_619)
);

INVx8_ASAP7_75t_L g620 ( 
.A(n_466),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_494),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_465),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_495),
.A2(n_322),
.B1(n_182),
.B2(n_193),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_481),
.A2(n_307),
.B1(n_296),
.B2(n_277),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_450),
.A2(n_448),
.B1(n_475),
.B2(n_473),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_499),
.B(n_183),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_448),
.B(n_475),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_454),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_499),
.B(n_184),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_454),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_454),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_465),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_428),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_467),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_467),
.Y(n_635)
);

AND3x4_ASAP7_75t_L g636 ( 
.A(n_504),
.B(n_281),
.C(n_190),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_459),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_468),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_475),
.B(n_230),
.Y(n_640)
);

BUFx8_ASAP7_75t_SL g641 ( 
.A(n_504),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_482),
.B(n_184),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_459),
.Y(n_643)
);

NAND2x1p5_ASAP7_75t_L g644 ( 
.A(n_456),
.B(n_235),
.Y(n_644)
);

AND2x2_ASAP7_75t_SL g645 ( 
.A(n_450),
.B(n_240),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_459),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_500),
.Y(n_647)
);

BUFx4f_ASAP7_75t_L g648 ( 
.A(n_434),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_500),
.A2(n_182),
.B1(n_197),
.B2(n_335),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_482),
.B(n_185),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_482),
.B(n_190),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_459),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_459),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_469),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_500),
.B(n_185),
.Y(n_655)
);

BUFx6f_ASAP7_75t_SL g656 ( 
.A(n_497),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_431),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_537),
.A2(n_616),
.B1(n_621),
.B2(n_591),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_657),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_537),
.A2(n_456),
.B1(n_469),
.B2(n_471),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_657),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_616),
.B(n_456),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_537),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_594),
.B(n_186),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_537),
.B(n_489),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_561),
.B(n_360),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_592),
.A2(n_497),
.B1(n_440),
.B2(n_478),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_505),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_531),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_592),
.B(n_591),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_521),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_506),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_594),
.B(n_186),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_533),
.B(n_312),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_510),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_510),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_512),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_512),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_533),
.B(n_312),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_621),
.B(n_489),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_545),
.B(n_489),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_564),
.B(n_366),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_489),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_513),
.Y(n_684)
);

OAI221xp5_ASAP7_75t_L g685 ( 
.A1(n_640),
.A2(n_197),
.B1(n_322),
.B2(n_320),
.C(n_319),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_538),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_513),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_559),
.A2(n_489),
.B(n_471),
.C(n_478),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_509),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_569),
.B(n_440),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_532),
.A2(n_332),
.B1(n_319),
.B2(n_318),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_521),
.B(n_320),
.C(n_193),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_540),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_625),
.B(n_457),
.Y(n_694)
);

INVxp33_ASAP7_75t_L g695 ( 
.A(n_535),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_592),
.B(n_457),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_592),
.B(n_474),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_509),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_550),
.B(n_474),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_524),
.B(n_476),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_604),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_604),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_618),
.A2(n_476),
.B1(n_484),
.B2(n_479),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_524),
.B(n_479),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_595),
.B(n_376),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_642),
.A2(n_484),
.B(n_480),
.C(n_461),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_533),
.B(n_314),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_532),
.B(n_627),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_535),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_578),
.B(n_461),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_593),
.B(n_383),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_539),
.B(n_480),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_540),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_539),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_620),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_578),
.B(n_387),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_618),
.A2(n_488),
.B1(n_477),
.B2(n_483),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_508),
.A2(n_314),
.B1(n_325),
.B2(n_336),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_538),
.B(n_325),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_574),
.A2(n_483),
.B(n_445),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_593),
.B(n_390),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_528),
.B(n_398),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_618),
.A2(n_488),
.B1(n_477),
.B2(n_483),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_549),
.B(n_402),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_544),
.B(n_477),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_516),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_627),
.B(n_483),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_544),
.B(n_488),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_596),
.B(n_332),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_516),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_617),
.B(n_276),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_538),
.A2(n_431),
.B(n_464),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_618),
.A2(n_455),
.B1(n_464),
.B2(n_431),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_654),
.B(n_597),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_538),
.B(n_327),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_654),
.B(n_327),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_523),
.B(n_328),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_582),
.B(n_328),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_577),
.B(n_455),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_582),
.B(n_586),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_575),
.B(n_329),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_523),
.B(n_329),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_532),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_582),
.B(n_333),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_575),
.B(n_333),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_604),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_532),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_525),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_575),
.B(n_336),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_598),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_532),
.A2(n_645),
.B1(n_647),
.B2(n_577),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_586),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_645),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_647),
.A2(n_431),
.B(n_464),
.C(n_435),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_525),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_575),
.B(n_241),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_586),
.B(n_455),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_611),
.B(n_242),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_547),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_614),
.B(n_435),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_614),
.B(n_435),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_641),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_614),
.B(n_435),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_556),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_547),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_612),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_554),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_650),
.A2(n_464),
.B(n_445),
.C(n_441),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_612),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_611),
.B(n_244),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_612),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_554),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_645),
.B(n_439),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_523),
.B(n_507),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_651),
.A2(n_248),
.B1(n_331),
.B2(n_317),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_610),
.B(n_439),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_542),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_611),
.B(n_255),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_610),
.B(n_439),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_558),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_583),
.B(n_261),
.C(n_285),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_558),
.Y(n_782)
);

BUFx12f_ASAP7_75t_L g783 ( 
.A(n_527),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_556),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_518),
.B(n_439),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_649),
.A2(n_264),
.B1(n_278),
.B2(n_283),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_651),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_518),
.B(n_441),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_515),
.A2(n_445),
.B1(n_441),
.B2(n_310),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_557),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_518),
.B(n_441),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_523),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_518),
.B(n_445),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_526),
.A2(n_529),
.B1(n_541),
.B2(n_534),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_518),
.B(n_199),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_565),
.A2(n_301),
.B(n_452),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_518),
.B(n_205),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_649),
.B(n_428),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_543),
.B(n_210),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_655),
.B(n_213),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_623),
.B(n_434),
.C(n_452),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_560),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_518),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_515),
.A2(n_466),
.B1(n_452),
.B2(n_437),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_L g805 ( 
.A(n_519),
.B(n_548),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_519),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_630),
.B(n_216),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_556),
.B(n_11),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_579),
.B(n_12),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_630),
.B(n_217),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_611),
.B(n_434),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_515),
.A2(n_466),
.B1(n_452),
.B2(n_437),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_560),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_567),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_630),
.B(n_222),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_637),
.B(n_224),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_637),
.B(n_225),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_562),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_626),
.B(n_228),
.C(n_311),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_543),
.B(n_231),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_629),
.B(n_232),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_600),
.B(n_434),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_L g823 ( 
.A(n_644),
.B(n_192),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_511),
.A2(n_272),
.B1(n_233),
.B2(n_234),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_SL g825 ( 
.A1(n_662),
.A2(n_584),
.B(n_581),
.C(n_613),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_809),
.A2(n_786),
.B1(n_670),
.B2(n_708),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_729),
.B(n_624),
.C(n_603),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_675),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_663),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_751),
.A2(n_600),
.B1(n_653),
.B2(n_514),
.Y(n_830)
);

OAI21xp33_ASAP7_75t_L g831 ( 
.A1(n_695),
.A2(n_530),
.B(n_607),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_743),
.B(n_517),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_681),
.A2(n_615),
.B(n_648),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_690),
.B(n_553),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_700),
.B(n_553),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_743),
.B(n_747),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_663),
.A2(n_676),
.B1(n_678),
.B2(n_677),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_734),
.A2(n_648),
.B(n_643),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_659),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_754),
.A2(n_644),
.B(n_643),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_704),
.B(n_580),
.Y(n_841)
);

AO22x1_ASAP7_75t_L g842 ( 
.A1(n_682),
.A2(n_636),
.B1(n_580),
.B2(n_587),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_709),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_714),
.A2(n_527),
.B1(n_656),
.B2(n_514),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_740),
.A2(n_648),
.B(n_588),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_811),
.A2(n_570),
.B(n_602),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_747),
.B(n_517),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_811),
.A2(n_570),
.B(n_602),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_686),
.B(n_517),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_712),
.B(n_653),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_661),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_684),
.A2(n_653),
.B1(n_514),
.B2(n_563),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_725),
.B(n_562),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_709),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_714),
.A2(n_656),
.B1(n_636),
.B2(n_601),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_686),
.B(n_517),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_750),
.B(n_656),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_685),
.A2(n_601),
.B(n_563),
.C(n_566),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_674),
.A2(n_707),
.B(n_679),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_728),
.B(n_710),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_696),
.B(n_566),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_669),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_671),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_774),
.B(n_636),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_784),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_670),
.B(n_568),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_787),
.B(n_695),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_739),
.B(n_568),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_687),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_674),
.A2(n_652),
.B(n_646),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_686),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_668),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_658),
.B(n_573),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_693),
.Y(n_875)
);

NOR2x1p5_ASAP7_75t_SL g876 ( 
.A(n_668),
.B(n_567),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_716),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_792),
.B(n_573),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_672),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_731),
.B(n_576),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_727),
.B(n_576),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_727),
.B(n_581),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_784),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_708),
.B(n_517),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_679),
.A2(n_652),
.B(n_646),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_707),
.A2(n_590),
.B(n_605),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_665),
.B(n_589),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_760),
.A2(n_590),
.B(n_605),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_761),
.A2(n_619),
.B(n_628),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_763),
.A2(n_619),
.B(n_628),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_708),
.B(n_552),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_701),
.B(n_552),
.Y(n_892)
);

AO21x1_ASAP7_75t_L g893 ( 
.A1(n_823),
.A2(n_639),
.B(n_638),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_669),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_713),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_757),
.A2(n_599),
.B(n_631),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_722),
.A2(n_639),
.B1(n_638),
.B2(n_635),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_777),
.A2(n_635),
.B1(n_634),
.B2(n_589),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_666),
.B(n_606),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_823),
.A2(n_599),
.B(n_631),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_665),
.B(n_606),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_L g902 ( 
.A1(n_718),
.A2(n_607),
.B(n_632),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_790),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_818),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_720),
.A2(n_522),
.B(n_536),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_701),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_705),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_732),
.A2(n_634),
.B(n_632),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_706),
.A2(n_660),
.B(n_781),
.C(n_775),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_724),
.A2(n_609),
.B1(n_622),
.B2(n_613),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_719),
.A2(n_555),
.B(n_522),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_711),
.B(n_622),
.C(n_609),
.Y(n_912)
);

AOI21x1_ASAP7_75t_L g913 ( 
.A1(n_773),
.A2(n_522),
.B(n_520),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_672),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_665),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_667),
.B(n_587),
.Y(n_916)
);

CKINVDCx11_ASAP7_75t_R g917 ( 
.A(n_783),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_719),
.A2(n_536),
.B(n_555),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_697),
.A2(n_520),
.B1(n_536),
.B2(n_546),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_735),
.A2(n_546),
.B(n_555),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_703),
.B(n_587),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_735),
.A2(n_520),
.B(n_546),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_699),
.B(n_552),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_792),
.B(n_552),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_683),
.B(n_552),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_721),
.B(n_572),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_694),
.B(n_572),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_680),
.B(n_572),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_741),
.A2(n_572),
.B(n_633),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_741),
.A2(n_572),
.B(n_633),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_L g931 ( 
.A(n_752),
.B(n_633),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_737),
.B(n_428),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_745),
.A2(n_633),
.B(n_620),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_702),
.B(n_633),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_702),
.B(n_620),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_784),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_808),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_689),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_742),
.B(n_428),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_746),
.B(n_620),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_785),
.A2(n_428),
.B(n_429),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_746),
.B(n_13),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_701),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_691),
.A2(n_13),
.B(n_14),
.C(n_17),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_801),
.A2(n_466),
.B(n_608),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_769),
.B(n_620),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_762),
.B(n_19),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_788),
.A2(n_428),
.B(n_429),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_715),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_745),
.A2(n_237),
.B(n_305),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_749),
.A2(n_726),
.B(n_698),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_SL g952 ( 
.A1(n_749),
.A2(n_21),
.B(n_23),
.C(n_27),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_726),
.A2(n_292),
.B(n_247),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_730),
.A2(n_293),
.B(n_250),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_692),
.B(n_428),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_730),
.A2(n_294),
.B(n_254),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_800),
.A2(n_434),
.B(n_452),
.C(n_437),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_736),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_771),
.B(n_701),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_738),
.A2(n_27),
.B(n_30),
.C(n_34),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_766),
.B(n_263),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_748),
.A2(n_298),
.B(n_257),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_748),
.A2(n_299),
.B(n_268),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_766),
.B(n_270),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_783),
.B(n_428),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_688),
.A2(n_466),
.B(n_585),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_755),
.A2(n_280),
.B(n_291),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_753),
.B(n_275),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_808),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_808),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_752),
.B(n_295),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_768),
.A2(n_802),
.B(n_780),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_798),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_755),
.A2(n_608),
.B(n_585),
.Y(n_974)
);

NOR2xp67_ASAP7_75t_L g975 ( 
.A(n_794),
.B(n_608),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_752),
.B(n_717),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_L g977 ( 
.A(n_821),
.B(n_297),
.C(n_36),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_715),
.B(n_437),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_759),
.A2(n_608),
.B(n_585),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_723),
.B(n_35),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_715),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_744),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_798),
.B(n_39),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_765),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_789),
.B(n_41),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_767),
.A2(n_437),
.B1(n_434),
.B2(n_436),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_SL g987 ( 
.A1(n_756),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_772),
.A2(n_608),
.B(n_585),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_805),
.A2(n_466),
.B1(n_434),
.B2(n_437),
.Y(n_989)
);

AND2x2_ASAP7_75t_SL g990 ( 
.A(n_799),
.B(n_240),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_782),
.B(n_436),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_806),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_664),
.B(n_42),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_782),
.B(n_436),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_664),
.B(n_46),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_673),
.B(n_47),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_813),
.A2(n_814),
.B(n_822),
.Y(n_997)
);

AOI21x1_ASAP7_75t_L g998 ( 
.A1(n_913),
.A2(n_893),
.B(n_859),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_828),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_863),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_899),
.B(n_820),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_869),
.Y(n_1002)
);

NOR3xp33_ASAP7_75t_SL g1003 ( 
.A(n_862),
.B(n_807),
.C(n_810),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_860),
.B(n_673),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_907),
.B(n_854),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_912),
.A2(n_819),
.B(n_817),
.C(n_816),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_880),
.A2(n_778),
.B(n_756),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_875),
.Y(n_1008)
);

BUFx12f_ASAP7_75t_L g1009 ( 
.A(n_917),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_912),
.B(n_779),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_853),
.A2(n_778),
.B(n_758),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_895),
.Y(n_1012)
);

INVx6_ASAP7_75t_L g1013 ( 
.A(n_965),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_843),
.B(n_803),
.Y(n_1014)
);

CKINVDCx14_ASAP7_75t_R g1015 ( 
.A(n_894),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_867),
.B(n_804),
.Y(n_1016)
);

AO22x1_ASAP7_75t_L g1017 ( 
.A1(n_977),
.A2(n_764),
.B1(n_803),
.B2(n_795),
.Y(n_1017)
);

OAI22x1_ASAP7_75t_L g1018 ( 
.A1(n_855),
.A2(n_822),
.B1(n_758),
.B2(n_770),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_996),
.A2(n_770),
.B(n_815),
.C(n_776),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_996),
.A2(n_796),
.B(n_733),
.C(n_791),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_861),
.A2(n_812),
.B1(n_824),
.B2(n_793),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_937),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_827),
.A2(n_797),
.B(n_436),
.C(n_434),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_857),
.B(n_585),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_915),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_881),
.A2(n_436),
.B1(n_437),
.B2(n_452),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_877),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_871),
.A2(n_240),
.B(n_551),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_903),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_864),
.B(n_429),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_969),
.B(n_970),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_857),
.B(n_571),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_926),
.B(n_47),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_864),
.B(n_48),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_871),
.A2(n_571),
.B(n_551),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_882),
.A2(n_868),
.B1(n_909),
.B2(n_866),
.Y(n_1036)
);

AO21x1_ASAP7_75t_L g1037 ( 
.A1(n_983),
.A2(n_192),
.B(n_238),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_931),
.A2(n_571),
.B(n_551),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_826),
.B(n_48),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_990),
.A2(n_571),
.B1(n_551),
.B2(n_429),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_904),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_943),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_943),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_SL g1044 ( 
.A(n_990),
.B(n_571),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_909),
.A2(n_436),
.B1(n_452),
.B2(n_429),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_878),
.A2(n_436),
.B(n_429),
.C(n_571),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_908),
.A2(n_551),
.B(n_429),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_826),
.B(n_429),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_947),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_SL g1050 ( 
.A1(n_849),
.A2(n_856),
.B(n_978),
.C(n_850),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_965),
.B(n_551),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_833),
.A2(n_49),
.B(n_52),
.C(n_54),
.Y(n_1052)
);

AOI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_993),
.A2(n_52),
.B(n_54),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_900),
.A2(n_118),
.B(n_66),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_834),
.B(n_238),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_923),
.A2(n_122),
.B(n_78),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_965),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_943),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_897),
.A2(n_58),
.B1(n_238),
.B2(n_192),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_840),
.A2(n_238),
.B(n_192),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_958),
.B(n_238),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_992),
.B(n_82),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_838),
.A2(n_85),
.B(n_89),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_831),
.B(n_104),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_865),
.B(n_133),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_829),
.B(n_192),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_884),
.B(n_136),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_829),
.B(n_192),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_943),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_SL g1070 ( 
.A(n_906),
.B(n_192),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_928),
.A2(n_140),
.B(n_147),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_910),
.A2(n_158),
.B1(n_238),
.B2(n_874),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_942),
.B(n_238),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_902),
.A2(n_238),
.B(n_995),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_SL g1075 ( 
.A1(n_960),
.A2(n_982),
.B(n_858),
.C(n_878),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_925),
.A2(n_845),
.B(n_825),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_906),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_887),
.A2(n_901),
.B1(n_837),
.B2(n_898),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_SL g1079 ( 
.A1(n_985),
.A2(n_942),
.B1(n_980),
.B2(n_844),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_955),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_865),
.B(n_936),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_884),
.B(n_891),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_842),
.B(n_973),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_896),
.A2(n_889),
.B(n_888),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_890),
.A2(n_927),
.B(n_978),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_929),
.A2(n_930),
.B(n_852),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_959),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_972),
.A2(n_885),
.B(n_886),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_865),
.Y(n_1089)
);

OAI22x1_ASAP7_75t_L g1090 ( 
.A1(n_891),
.A2(n_989),
.B1(n_836),
.B2(n_959),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_872),
.Y(n_1091)
);

BUFx8_ASAP7_75t_L g1092 ( 
.A(n_865),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_961),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_870),
.A2(n_848),
.B(n_846),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_835),
.A2(n_841),
.B1(n_976),
.B2(n_973),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_944),
.A2(n_924),
.B(n_876),
.C(n_975),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_936),
.Y(n_1097)
);

INVx5_ASAP7_75t_L g1098 ( 
.A(n_936),
.Y(n_1098)
);

AO22x1_ASAP7_75t_L g1099 ( 
.A1(n_873),
.A2(n_883),
.B1(n_936),
.B2(n_968),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_981),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_879),
.B(n_914),
.Y(n_1101)
);

OAI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_921),
.A2(n_916),
.B1(n_964),
.B2(n_830),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_911),
.A2(n_922),
.B(n_918),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_938),
.B(n_984),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_981),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_924),
.A2(n_951),
.B(n_934),
.C(n_997),
.Y(n_1106)
);

HAxp5_ASAP7_75t_L g1107 ( 
.A(n_987),
.B(n_952),
.CON(n_1107),
.SN(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_839),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_932),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_981),
.B(n_934),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_873),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_957),
.A2(n_939),
.B(n_933),
.C(n_832),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_981),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_883),
.B(n_949),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_892),
.Y(n_1115)
);

INVx6_ASAP7_75t_L g1116 ( 
.A(n_836),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_832),
.A2(n_847),
.B1(n_851),
.B2(n_892),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_SL g1118 ( 
.A(n_950),
.B(n_971),
.C(n_963),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_847),
.B(n_940),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_949),
.B(n_935),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_952),
.A2(n_987),
.B(n_957),
.C(n_919),
.Y(n_1121)
);

BUFx4f_ASAP7_75t_L g1122 ( 
.A(n_946),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_991),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_994),
.B(n_962),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_994),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_986),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_966),
.B(n_954),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_953),
.B(n_956),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_967),
.B(n_920),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_941),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_945),
.B(n_979),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_SL g1132 ( 
.A(n_988),
.B(n_905),
.C(n_948),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_974),
.A2(n_861),
.B1(n_882),
.B2(n_881),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_907),
.B(n_682),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_915),
.B(n_708),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_907),
.B(n_709),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_915),
.B(n_708),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_894),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_863),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_912),
.A2(n_545),
.B(n_496),
.C(n_564),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_L g1141 ( 
.A(n_907),
.B(n_750),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1009),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_SL g1143 ( 
.A1(n_1129),
.A2(n_1059),
.B(n_1053),
.C(n_1128),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1134),
.B(n_1005),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1072),
.A2(n_1007),
.B(n_1019),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1088),
.A2(n_1085),
.B(n_1084),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1141),
.B(n_1004),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1036),
.A2(n_1133),
.B(n_1076),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1094),
.A2(n_1086),
.B(n_1060),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_SL g1150 ( 
.A(n_1034),
.B(n_1140),
.C(n_1001),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1036),
.A2(n_1133),
.B(n_1044),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_1103),
.A2(n_1074),
.B(n_1023),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1044),
.A2(n_1045),
.B(n_1072),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1138),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1092),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1000),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1139),
.B(n_1016),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1045),
.A2(n_1050),
.B(n_1078),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1078),
.A2(n_1106),
.B(n_1010),
.Y(n_1159)
);

INVx3_ASAP7_75t_SL g1160 ( 
.A(n_1136),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_1113),
.B(n_1098),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1027),
.B(n_1022),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1037),
.A2(n_1102),
.B(n_998),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_999),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1015),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1130),
.A2(n_1132),
.B(n_1112),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1011),
.A2(n_1006),
.B(n_1026),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1093),
.B(n_1002),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1131),
.A2(n_1063),
.B(n_1047),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1026),
.A2(n_1118),
.B(n_1120),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1126),
.A2(n_1079),
.B1(n_1049),
.B2(n_1082),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1029),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1120),
.A2(n_1096),
.B(n_1046),
.Y(n_1174)
);

AOI211x1_ASAP7_75t_L g1175 ( 
.A1(n_1053),
.A2(n_1041),
.B(n_1033),
.C(n_1014),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1075),
.A2(n_1107),
.B(n_1003),
.C(n_1121),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1087),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_SL g1178 ( 
.A1(n_1095),
.A2(n_1020),
.B(n_1021),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1127),
.A2(n_1122),
.B(n_1054),
.Y(n_1179)
);

BUFx2_ASAP7_75t_SL g1180 ( 
.A(n_1098),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1135),
.B(n_1137),
.Y(n_1181)
);

BUFx8_ASAP7_75t_L g1182 ( 
.A(n_1042),
.Y(n_1182)
);

AO32x2_ASAP7_75t_L g1183 ( 
.A1(n_1095),
.A2(n_1080),
.A3(n_1021),
.B1(n_1058),
.B2(n_1111),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1122),
.A2(n_1028),
.B(n_1124),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_1098),
.Y(n_1185)
);

OAI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1073),
.A2(n_1018),
.B(n_1067),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1116),
.A2(n_1031),
.B1(n_1013),
.B2(n_1025),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1110),
.A2(n_1017),
.B(n_1056),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1042),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1055),
.A2(n_1071),
.B(n_1119),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1052),
.A2(n_1061),
.B(n_1030),
.C(n_1123),
.Y(n_1191)
);

CKINVDCx11_ASAP7_75t_R g1192 ( 
.A(n_1042),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1092),
.Y(n_1193)
);

AO32x2_ASAP7_75t_L g1194 ( 
.A1(n_1058),
.A2(n_1111),
.A3(n_1077),
.B1(n_1117),
.B2(n_1090),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1109),
.A2(n_1070),
.B(n_1099),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1113),
.B(n_1057),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1109),
.A2(n_1083),
.B(n_1032),
.C(n_1024),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_1100),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1051),
.B(n_1031),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1116),
.B(n_1062),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1043),
.B(n_1115),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1091),
.B(n_1108),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_SL g1203 ( 
.A1(n_1066),
.A2(n_1068),
.B(n_1043),
.C(n_1125),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1081),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1070),
.A2(n_1035),
.B(n_1038),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1051),
.B(n_1077),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1114),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1048),
.B(n_1069),
.Y(n_1208)
);

AO32x2_ASAP7_75t_L g1209 ( 
.A1(n_1115),
.A2(n_1104),
.A3(n_1101),
.B1(n_1065),
.B2(n_1089),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1069),
.B(n_1089),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1040),
.A2(n_1115),
.B(n_1089),
.Y(n_1211)
);

AO32x2_ASAP7_75t_L g1212 ( 
.A1(n_1069),
.A2(n_1045),
.A3(n_1059),
.B1(n_1095),
.B2(n_1036),
.Y(n_1212)
);

AO32x2_ASAP7_75t_L g1213 ( 
.A1(n_1097),
.A2(n_1045),
.A3(n_1059),
.B1(n_1095),
.B2(n_1036),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1097),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1100),
.B(n_1105),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1105),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1134),
.B(n_899),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1001),
.B(n_709),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1134),
.A2(n_750),
.B1(n_880),
.B2(n_564),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1220)
);

AO32x2_ASAP7_75t_L g1221 ( 
.A1(n_1045),
.A2(n_1059),
.A3(n_1095),
.B1(n_1036),
.B2(n_1079),
.Y(n_1221)
);

INVx5_ASAP7_75t_L g1222 ( 
.A(n_1013),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1072),
.A2(n_750),
.B(n_880),
.Y(n_1223)
);

CKINVDCx11_ASAP7_75t_R g1224 ( 
.A(n_1009),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1098),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1113),
.B(n_937),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1037),
.A2(n_1023),
.A3(n_893),
.B(n_1072),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1134),
.B(n_682),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1134),
.A2(n_827),
.B(n_996),
.C(n_1072),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1134),
.A2(n_827),
.B(n_996),
.C(n_1072),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_SL g1232 ( 
.A(n_1138),
.B(n_669),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_999),
.Y(n_1234)
);

AO21x1_ASAP7_75t_L g1235 ( 
.A1(n_1072),
.A2(n_1059),
.B(n_1064),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1009),
.B(n_842),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1134),
.B(n_899),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_R g1238 ( 
.A(n_1138),
.B(n_1015),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_SL g1239 ( 
.A1(n_1010),
.A2(n_1072),
.B(n_893),
.Y(n_1239)
);

INVx3_ASAP7_75t_SL g1240 ( 
.A(n_1138),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1088),
.A2(n_1085),
.B(n_1084),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1134),
.A2(n_827),
.B(n_996),
.C(n_1072),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1134),
.B(n_899),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_999),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_999),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1072),
.A2(n_750),
.B(n_880),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_999),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_L g1248 ( 
.A(n_1009),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1072),
.A2(n_750),
.B(n_880),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1134),
.B(n_682),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_1072),
.A2(n_1059),
.B(n_1064),
.Y(n_1251)
);

AOI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_1134),
.A2(n_682),
.B1(n_564),
.B2(n_666),
.C(n_786),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_999),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1134),
.B(n_682),
.Y(n_1254)
);

NOR3xp33_ASAP7_75t_L g1255 ( 
.A(n_1134),
.B(n_682),
.C(n_564),
.Y(n_1255)
);

AOI221xp5_ASAP7_75t_L g1256 ( 
.A1(n_1134),
.A2(n_682),
.B1(n_564),
.B2(n_666),
.C(n_786),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1009),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_SL g1260 ( 
.A(n_1138),
.B(n_669),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1098),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1086),
.A2(n_1076),
.B(n_1084),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_999),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1088),
.A2(n_1085),
.B(n_1084),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_999),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_L g1267 ( 
.A1(n_998),
.A2(n_1076),
.B(n_1088),
.Y(n_1267)
);

BUFx2_ASAP7_75t_R g1268 ( 
.A(n_1138),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1037),
.A2(n_1023),
.A3(n_893),
.B(n_1072),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1072),
.A2(n_750),
.B(n_880),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_999),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1138),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1134),
.A2(n_750),
.B1(n_880),
.B2(n_564),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1140),
.A2(n_750),
.B(n_564),
.C(n_1134),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1134),
.A2(n_827),
.B(n_996),
.C(n_1072),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1037),
.A2(n_1023),
.A3(n_893),
.B(n_1072),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1037),
.A2(n_1023),
.A3(n_893),
.B(n_1072),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1098),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1084),
.A2(n_594),
.B(n_533),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1072),
.A2(n_750),
.B(n_880),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1134),
.B(n_521),
.Y(n_1287)
);

NOR4xp25_ASAP7_75t_L g1288 ( 
.A(n_1059),
.B(n_944),
.C(n_831),
.D(n_1034),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1088),
.A2(n_1085),
.B(n_1084),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1134),
.B(n_682),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1072),
.A2(n_750),
.B(n_880),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1134),
.A2(n_827),
.B(n_996),
.C(n_1072),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1000),
.B(n_854),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1072),
.A2(n_514),
.B(n_594),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1182),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1224),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1252),
.B2(n_1256),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1229),
.A2(n_1250),
.B1(n_1290),
.B2(n_1254),
.Y(n_1298)
);

BUFx4f_ASAP7_75t_SL g1299 ( 
.A(n_1240),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1165),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1255),
.A2(n_1172),
.B1(n_1286),
.B2(n_1270),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1223),
.A2(n_1249),
.B1(n_1246),
.B2(n_1291),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1219),
.A2(n_1278),
.B1(n_1186),
.B2(n_1153),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1238),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_1192),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1217),
.A2(n_1237),
.B1(n_1243),
.B2(n_1157),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1145),
.A2(n_1239),
.B1(n_1144),
.B2(n_1221),
.Y(n_1307)
);

INVx3_ASAP7_75t_SL g1308 ( 
.A(n_1160),
.Y(n_1308)
);

INVx6_ASAP7_75t_L g1309 ( 
.A(n_1182),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1169),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1177),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1142),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1155),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1257),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1293),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1159),
.A2(n_1168),
.B1(n_1236),
.B2(n_1151),
.Y(n_1316)
);

BUFx2_ASAP7_75t_SL g1317 ( 
.A(n_1276),
.Y(n_1317)
);

BUFx2_ASAP7_75t_SL g1318 ( 
.A(n_1207),
.Y(n_1318)
);

CKINVDCx14_ASAP7_75t_R g1319 ( 
.A(n_1248),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1230),
.A2(n_1292),
.B1(n_1280),
.B2(n_1231),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1193),
.Y(n_1321)
);

INVx4_ASAP7_75t_SL g1322 ( 
.A(n_1225),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1164),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1166),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1287),
.B(n_1156),
.Y(n_1325)
);

BUFx2_ASAP7_75t_SL g1326 ( 
.A(n_1222),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1268),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1248),
.Y(n_1328)
);

CKINVDCx6p67_ASAP7_75t_R g1329 ( 
.A(n_1236),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1221),
.A2(n_1158),
.B1(n_1212),
.B2(n_1213),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1204),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1173),
.A2(n_1234),
.B1(n_1245),
.B2(n_1244),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1247),
.A2(n_1253),
.B1(n_1266),
.B2(n_1264),
.Y(n_1333)
);

INVx3_ASAP7_75t_SL g1334 ( 
.A(n_1218),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1215),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1162),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1275),
.A2(n_1150),
.B1(n_1147),
.B2(n_1200),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1199),
.A2(n_1221),
.B1(n_1181),
.B2(n_1202),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1232),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1208),
.A2(n_1174),
.B1(n_1187),
.B2(n_1242),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1222),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1225),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1216),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1175),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1214),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1288),
.A2(n_1260),
.B1(n_1206),
.B2(n_1201),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1212),
.A2(n_1213),
.B1(n_1195),
.B2(n_1178),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1209),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1212),
.A2(n_1213),
.B1(n_1148),
.B2(n_1167),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1171),
.A2(n_1179),
.B1(n_1163),
.B2(n_1184),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1189),
.Y(n_1351)
);

CKINVDCx6p67_ASAP7_75t_R g1352 ( 
.A(n_1180),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1163),
.A2(n_1152),
.B1(n_1226),
.B2(n_1166),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1152),
.A2(n_1211),
.B1(n_1294),
.B2(n_1188),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1210),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1143),
.A2(n_1183),
.B1(n_1176),
.B2(n_1196),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1161),
.Y(n_1357)
);

BUFx2_ASAP7_75t_SL g1358 ( 
.A(n_1185),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1198),
.Y(n_1359)
);

BUFx10_ASAP7_75t_L g1360 ( 
.A(n_1198),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1185),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1190),
.A2(n_1261),
.B1(n_1284),
.B2(n_1279),
.Y(n_1362)
);

INVx6_ASAP7_75t_L g1363 ( 
.A(n_1261),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1194),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1197),
.A2(n_1284),
.B1(n_1203),
.B2(n_1205),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1191),
.B(n_1283),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1267),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1220),
.A2(n_1263),
.B1(n_1285),
.B2(n_1274),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1183),
.A2(n_1262),
.B1(n_1282),
.B2(n_1233),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1194),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1227),
.A2(n_1258),
.B1(n_1272),
.B2(n_1277),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_SL g1372 ( 
.A(n_1228),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1271),
.B2(n_1170),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1146),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1269),
.A2(n_1281),
.B1(n_1283),
.B2(n_1265),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1269),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1241),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1289),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1283),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1149),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1192),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1256),
.B2(n_1252),
.Y(n_1382)
);

AO22x1_ASAP7_75t_L g1383 ( 
.A1(n_1229),
.A2(n_1254),
.B1(n_1250),
.B2(n_1290),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1252),
.A2(n_1256),
.B(n_1250),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1256),
.B2(n_1252),
.Y(n_1385)
);

CKINVDCx11_ASAP7_75t_R g1386 ( 
.A(n_1224),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1229),
.B(n_1250),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1256),
.B2(n_1252),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1224),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1224),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1229),
.A2(n_1250),
.B1(n_1290),
.B2(n_1254),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1252),
.A2(n_1256),
.B(n_1250),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1182),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1256),
.B2(n_1252),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1154),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1224),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_SL g1397 ( 
.A(n_1182),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1252),
.A2(n_1256),
.B(n_1250),
.Y(n_1398)
);

BUFx8_ASAP7_75t_L g1399 ( 
.A(n_1142),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1172),
.A2(n_1039),
.B1(n_729),
.B2(n_1044),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1256),
.B2(n_1252),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1256),
.B2(n_1252),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1169),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1229),
.A2(n_1250),
.B1(n_1290),
.B2(n_1254),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1229),
.A2(n_1250),
.B1(n_1290),
.B2(n_1254),
.Y(n_1405)
);

INVx4_ASAP7_75t_SL g1406 ( 
.A(n_1225),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1169),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1224),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1192),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1229),
.A2(n_809),
.B1(n_682),
.B2(n_990),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1192),
.Y(n_1411)
);

BUFx10_ASAP7_75t_L g1412 ( 
.A(n_1165),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1182),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1229),
.A2(n_1250),
.B1(n_1290),
.B2(n_1254),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1224),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1410),
.A2(n_1405),
.B1(n_1400),
.B2(n_1297),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1307),
.B(n_1302),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1367),
.A2(n_1366),
.B(n_1377),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1386),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1350),
.A2(n_1371),
.B(n_1368),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1384),
.B(n_1392),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1379),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1367),
.A2(n_1380),
.B(n_1320),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1323),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1376),
.A2(n_1372),
.B1(n_1414),
.B2(n_1298),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1350),
.A2(n_1379),
.B(n_1369),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1324),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1374),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1335),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1364),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1348),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1369),
.A2(n_1373),
.B(n_1354),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1330),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1330),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1378),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1372),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1349),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1307),
.B(n_1302),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1344),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1375),
.B(n_1347),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1347),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1363),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1410),
.A2(n_1400),
.B1(n_1401),
.B2(n_1297),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1353),
.A2(n_1354),
.B(n_1373),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1343),
.Y(n_1446)
);

CKINVDCx14_ASAP7_75t_R g1447 ( 
.A(n_1319),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1332),
.Y(n_1448)
);

AO21x1_ASAP7_75t_L g1449 ( 
.A1(n_1398),
.A2(n_1391),
.B(n_1365),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1353),
.B(n_1322),
.Y(n_1450)
);

OAI222xp33_ASAP7_75t_L g1451 ( 
.A1(n_1382),
.A2(n_1385),
.B1(n_1402),
.B2(n_1388),
.C1(n_1394),
.C2(n_1401),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1316),
.A2(n_1362),
.B(n_1340),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1389),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1332),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1316),
.A2(n_1362),
.B(n_1340),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1333),
.B(n_1306),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1333),
.B(n_1306),
.Y(n_1457)
);

AO31x2_ASAP7_75t_L g1458 ( 
.A1(n_1355),
.A2(n_1310),
.A3(n_1407),
.B(n_1403),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1363),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1303),
.A2(n_1337),
.B(n_1382),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1356),
.B(n_1385),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1361),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1390),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1309),
.Y(n_1464)
);

NOR2xp67_ASAP7_75t_L g1465 ( 
.A(n_1337),
.B(n_1351),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1336),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1356),
.B(n_1388),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1394),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1315),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1402),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1325),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1338),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1345),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1338),
.A2(n_1301),
.B(n_1346),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1301),
.A2(n_1322),
.B(n_1406),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_SL g1476 ( 
.A1(n_1387),
.A2(n_1404),
.B(n_1383),
.C(n_1317),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1341),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1358),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1334),
.B(n_1409),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1334),
.A2(n_1329),
.B(n_1326),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1381),
.B(n_1409),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1359),
.A2(n_1360),
.B(n_1357),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1318),
.B(n_1311),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1352),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1381),
.B(n_1411),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1309),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1321),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1381),
.B(n_1409),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1309),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1393),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1381),
.B(n_1411),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1393),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1397),
.A2(n_1342),
.B(n_1413),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1409),
.A2(n_1411),
.B1(n_1327),
.B2(n_1305),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1411),
.B(n_1305),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1421),
.A2(n_1408),
.B1(n_1396),
.B2(n_1331),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1421),
.A2(n_1339),
.B1(n_1395),
.B2(n_1308),
.C(n_1328),
.Y(n_1497)
);

AOI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1417),
.A2(n_1438),
.B1(n_1461),
.B2(n_1467),
.C(n_1416),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1471),
.B(n_1469),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1449),
.A2(n_1295),
.B(n_1313),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1440),
.B(n_1413),
.Y(n_1501)
);

NOR2x1_ASAP7_75t_L g1502 ( 
.A(n_1486),
.B(n_1296),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1416),
.A2(n_1397),
.B1(n_1299),
.B2(n_1304),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1440),
.B(n_1424),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1471),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1429),
.B(n_1299),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1443),
.A2(n_1312),
.B1(n_1399),
.B2(n_1415),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1436),
.B(n_1399),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1417),
.A2(n_1300),
.B1(n_1314),
.B2(n_1412),
.C(n_1438),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1440),
.B(n_1412),
.Y(n_1510)
);

AO21x1_ASAP7_75t_L g1511 ( 
.A1(n_1461),
.A2(n_1467),
.B(n_1474),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1429),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1423),
.A2(n_1418),
.B(n_1437),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1424),
.B(n_1437),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1436),
.B(n_1450),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1474),
.A2(n_1443),
.B(n_1476),
.C(n_1460),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1430),
.B(n_1429),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1473),
.B(n_1479),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1474),
.A2(n_1476),
.B(n_1460),
.C(n_1467),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1449),
.A2(n_1461),
.B1(n_1425),
.B2(n_1470),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1480),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1469),
.B(n_1466),
.Y(n_1523)
);

AO32x2_ASAP7_75t_L g1524 ( 
.A1(n_1428),
.A2(n_1435),
.A3(n_1442),
.B1(n_1489),
.B2(n_1464),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1473),
.B(n_1479),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1425),
.A2(n_1468),
.B1(n_1470),
.B2(n_1449),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1466),
.B(n_1462),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1430),
.B(n_1439),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1420),
.A2(n_1432),
.B(n_1426),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1439),
.B(n_1445),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1458),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1468),
.A2(n_1494),
.B1(n_1492),
.B2(n_1464),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1439),
.B(n_1445),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1450),
.B(n_1475),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1420),
.A2(n_1432),
.B(n_1455),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1460),
.A2(n_1451),
.B(n_1455),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1452),
.A2(n_1455),
.B(n_1465),
.C(n_1475),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1458),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1491),
.A2(n_1482),
.B(n_1465),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1446),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1447),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1451),
.A2(n_1452),
.B(n_1420),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1452),
.A2(n_1475),
.B(n_1422),
.Y(n_1543)
);

AO32x2_ASAP7_75t_L g1544 ( 
.A1(n_1428),
.A2(n_1435),
.A3(n_1442),
.B1(n_1492),
.B2(n_1464),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1483),
.B(n_1478),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1479),
.B(n_1481),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1433),
.A2(n_1434),
.B1(n_1441),
.B2(n_1456),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1524),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1528),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1504),
.B(n_1444),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1498),
.A2(n_1433),
.B1(n_1434),
.B2(n_1441),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1504),
.B(n_1444),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1515),
.Y(n_1553)
);

BUFx4f_ASAP7_75t_SL g1554 ( 
.A(n_1541),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1540),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1526),
.A2(n_1457),
.B1(n_1456),
.B2(n_1472),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1444),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1530),
.B(n_1444),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1533),
.B(n_1444),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1505),
.B(n_1431),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1521),
.B(n_1459),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1511),
.A2(n_1536),
.B1(n_1456),
.B2(n_1457),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1535),
.B(n_1435),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1542),
.A2(n_1457),
.B1(n_1472),
.B2(n_1448),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1499),
.B(n_1431),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1500),
.B(n_1483),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1517),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1547),
.A2(n_1454),
.B1(n_1448),
.B2(n_1453),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1514),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1516),
.A2(n_1494),
.B1(n_1454),
.B2(n_1491),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1543),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1519),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1543),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1516),
.A2(n_1487),
.B1(n_1486),
.B2(n_1490),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1545),
.B(n_1427),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1560),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1560),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1548),
.A2(n_1510),
.B1(n_1501),
.B2(n_1532),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1566),
.B(n_1508),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1555),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1570),
.A2(n_1520),
.B(n_1574),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1555),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1562),
.A2(n_1547),
.B1(n_1509),
.B2(n_1534),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1556),
.A2(n_1520),
.B1(n_1537),
.B2(n_1507),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1548),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1556),
.A2(n_1537),
.B1(n_1497),
.B2(n_1496),
.C(n_1503),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1548),
.Y(n_1587)
);

NOR3xp33_ASAP7_75t_L g1588 ( 
.A(n_1570),
.B(n_1487),
.C(n_1523),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1572),
.B(n_1525),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1554),
.A2(n_1541),
.B1(n_1496),
.B2(n_1453),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1553),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1571),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1569),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1566),
.B(n_1512),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1513),
.Y(n_1595)
);

AOI322xp5_ASAP7_75t_L g1596 ( 
.A1(n_1551),
.A2(n_1562),
.A3(n_1568),
.B1(n_1561),
.B2(n_1564),
.C1(n_1552),
.C2(n_1550),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1572),
.B(n_1546),
.Y(n_1597)
);

INVx5_ASAP7_75t_L g1598 ( 
.A(n_1563),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1554),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1553),
.B(n_1510),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1601)
);

OAI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1575),
.A2(n_1527),
.B(n_1529),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1567),
.B(n_1524),
.Y(n_1603)
);

OAI33xp33_ASAP7_75t_L g1604 ( 
.A1(n_1561),
.A2(n_1506),
.A3(n_1484),
.B1(n_1419),
.B2(n_1531),
.B3(n_1538),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1568),
.A2(n_1539),
.B1(n_1501),
.B2(n_1522),
.C(n_1518),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1563),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1567),
.B(n_1524),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1557),
.B(n_1544),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1598),
.B(n_1557),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1608),
.B(n_1601),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1580),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1580),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1582),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1585),
.B(n_1565),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1608),
.B(n_1557),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1598),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1598),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1606),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1585),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1608),
.B(n_1558),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1598),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1598),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1601),
.B(n_1558),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1603),
.B(n_1558),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1586),
.A2(n_1551),
.B1(n_1564),
.B2(n_1575),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1587),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1603),
.B(n_1559),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1582),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1587),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1607),
.B(n_1559),
.Y(n_1631)
);

AOI211xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1590),
.A2(n_1574),
.B(n_1508),
.C(n_1485),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1607),
.B(n_1549),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1606),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1593),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1593),
.Y(n_1637)
);

INVxp33_ASAP7_75t_L g1638 ( 
.A(n_1625),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1600),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1628),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1628),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1621),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1621),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1610),
.B(n_1615),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1628),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1611),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1611),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1610),
.B(n_1600),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1615),
.B(n_1591),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1621),
.B(n_1581),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1615),
.B(n_1591),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1612),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1636),
.B(n_1576),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1618),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1620),
.B(n_1591),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1620),
.B(n_1591),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1618),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1618),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1632),
.B(n_1597),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1619),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1634),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1636),
.B(n_1577),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1614),
.B(n_1577),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1614),
.B(n_1595),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1613),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1632),
.A2(n_1586),
.B1(n_1625),
.B2(n_1584),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1635),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1635),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1619),
.B(n_1596),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1626),
.B(n_1596),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1614),
.B(n_1594),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1621),
.B(n_1616),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1626),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1634),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1638),
.B(n_1623),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_SL g1680 ( 
.A(n_1661),
.B(n_1590),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1644),
.B(n_1616),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1668),
.B(n_1623),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1640),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1685)
);

INVxp33_ASAP7_75t_L g1686 ( 
.A(n_1650),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1617),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1668),
.B(n_1623),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1650),
.B(n_1621),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1650),
.B(n_1453),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1641),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1662),
.B(n_1602),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1676),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1639),
.B(n_1617),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1651),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1641),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1671),
.A2(n_1581),
.B1(n_1578),
.B2(n_1584),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1650),
.B(n_1617),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1639),
.B(n_1622),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1671),
.B(n_1622),
.C(n_1602),
.D(n_1609),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1651),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1645),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1648),
.B(n_1622),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1651),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1653),
.B(n_1630),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1662),
.B(n_1633),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1656),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1645),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1646),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1656),
.Y(n_1711)
);

INVxp33_ASAP7_75t_L g1712 ( 
.A(n_1661),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1672),
.A2(n_1578),
.B1(n_1583),
.B2(n_1579),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1672),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1646),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1698),
.A2(n_1677),
.B(n_1588),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1710),
.Y(n_1717)
);

AOI21xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1683),
.A2(n_1688),
.B(n_1690),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1712),
.A2(n_1648),
.B1(n_1658),
.B2(n_1609),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1714),
.A2(n_1588),
.B1(n_1604),
.B2(n_1605),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1679),
.A2(n_1658),
.B1(n_1609),
.B2(n_1677),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1701),
.A2(n_1666),
.B1(n_1605),
.B2(n_1653),
.C(n_1664),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1710),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1707),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1681),
.B(n_1685),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1715),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1713),
.A2(n_1604),
.B1(n_1552),
.B2(n_1550),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1680),
.A2(n_1573),
.B1(n_1522),
.B2(n_1518),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1686),
.B(n_1463),
.Y(n_1729)
);

OAI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1693),
.A2(n_1666),
.B1(n_1664),
.B2(n_1534),
.Y(n_1730)
);

NAND3x2_ASAP7_75t_L g1731 ( 
.A(n_1689),
.B(n_1674),
.C(n_1656),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1689),
.A2(n_1676),
.B(n_1495),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1699),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1694),
.A2(n_1643),
.B(n_1642),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1715),
.Y(n_1735)
);

OAI21xp33_ASAP7_75t_L g1736 ( 
.A1(n_1681),
.A2(n_1674),
.B(n_1657),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1685),
.B(n_1696),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1699),
.B(n_1652),
.C(n_1647),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1706),
.B(n_1665),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1696),
.B(n_1702),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1689),
.A2(n_1699),
.B1(n_1711),
.B2(n_1708),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1725),
.B(n_1706),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1727),
.A2(n_1711),
.B1(n_1708),
.B2(n_1705),
.C(n_1702),
.Y(n_1743)
);

OAI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1720),
.A2(n_1705),
.B1(n_1709),
.B2(n_1692),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1716),
.A2(n_1729),
.B1(n_1730),
.B2(n_1737),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1724),
.B(n_1733),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1722),
.A2(n_1738),
.B(n_1718),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1733),
.B(n_1699),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1717),
.Y(n_1749)
);

AOI322xp5_ASAP7_75t_L g1750 ( 
.A1(n_1728),
.A2(n_1631),
.A3(n_1624),
.B1(n_1627),
.B2(n_1552),
.C1(n_1592),
.C2(n_1629),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1739),
.B(n_1689),
.Y(n_1751)
);

OAI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1732),
.A2(n_1709),
.B1(n_1684),
.B2(n_1703),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1736),
.B(n_1682),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1732),
.A2(n_1592),
.B(n_1703),
.C(n_1691),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1723),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1726),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1741),
.A2(n_1463),
.B(n_1642),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1734),
.A2(n_1700),
.B(n_1695),
.Y(n_1758)
);

O2A1O1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1735),
.A2(n_1692),
.B(n_1691),
.C(n_1697),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1740),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1721),
.A2(n_1684),
.B1(n_1697),
.B2(n_1629),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1742),
.B(n_1731),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1747),
.A2(n_1676),
.B(n_1719),
.Y(n_1763)
);

INVx3_ASAP7_75t_SL g1764 ( 
.A(n_1748),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1751),
.B(n_1682),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1744),
.A2(n_1463),
.B1(n_1447),
.B2(n_1695),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1759),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1746),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1760),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1755),
.B(n_1687),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1749),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1756),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1744),
.B(n_1687),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1745),
.C(n_1758),
.Y(n_1774)
);

NOR3xp33_ASAP7_75t_L g1775 ( 
.A(n_1769),
.B(n_1761),
.C(n_1752),
.Y(n_1775)
);

NOR3xp33_ASAP7_75t_L g1776 ( 
.A(n_1768),
.B(n_1761),
.C(n_1752),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1764),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1765),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1770),
.Y(n_1779)
);

NAND4xp25_ASAP7_75t_L g1780 ( 
.A(n_1766),
.B(n_1757),
.C(n_1753),
.D(n_1743),
.Y(n_1780)
);

NAND4xp25_ASAP7_75t_L g1781 ( 
.A(n_1766),
.B(n_1754),
.C(n_1750),
.D(n_1704),
.Y(n_1781)
);

NAND3xp33_ASAP7_75t_SL g1782 ( 
.A(n_1773),
.B(n_1676),
.C(n_1700),
.Y(n_1782)
);

INVx6_ASAP7_75t_L g1783 ( 
.A(n_1762),
.Y(n_1783)
);

NOR3xp33_ASAP7_75t_L g1784 ( 
.A(n_1774),
.B(n_1763),
.C(n_1771),
.Y(n_1784)
);

AOI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1776),
.A2(n_1772),
.B(n_1704),
.C(n_1495),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1775),
.A2(n_1643),
.B(n_1642),
.Y(n_1786)
);

AOI211xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1777),
.A2(n_1495),
.B(n_1484),
.C(n_1508),
.Y(n_1787)
);

AOI21xp33_ASAP7_75t_SL g1788 ( 
.A1(n_1778),
.A2(n_1643),
.B(n_1665),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1781),
.A2(n_1678),
.B1(n_1654),
.B2(n_1655),
.C(n_1659),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1784),
.A2(n_1782),
.B(n_1780),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_SL g1791 ( 
.A(n_1785),
.B(n_1779),
.C(n_1783),
.Y(n_1791)
);

NOR3xp33_ASAP7_75t_L g1792 ( 
.A(n_1788),
.B(n_1786),
.C(n_1789),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1787),
.B(n_1649),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1784),
.A2(n_1678),
.B1(n_1654),
.B2(n_1655),
.C(n_1659),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1785),
.A2(n_1599),
.B1(n_1477),
.B2(n_1609),
.Y(n_1795)
);

AND4x1_ASAP7_75t_L g1796 ( 
.A(n_1790),
.B(n_1485),
.C(n_1481),
.D(n_1488),
.Y(n_1796)
);

XNOR2xp5_ASAP7_75t_L g1797 ( 
.A(n_1791),
.B(n_1493),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1792),
.A2(n_1655),
.B(n_1654),
.Y(n_1798)
);

NOR2x1_ASAP7_75t_L g1799 ( 
.A(n_1793),
.B(n_1477),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1795),
.A2(n_1481),
.B1(n_1485),
.B2(n_1488),
.Y(n_1800)
);

XNOR2xp5_ASAP7_75t_L g1801 ( 
.A(n_1797),
.B(n_1794),
.Y(n_1801)
);

NAND4xp75_ASAP7_75t_L g1802 ( 
.A(n_1799),
.B(n_1488),
.C(n_1502),
.D(n_1649),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1796),
.B(n_1477),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1803),
.B(n_1798),
.Y(n_1804)
);

CKINVDCx20_ASAP7_75t_R g1805 ( 
.A(n_1804),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1801),
.B(n_1800),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1805),
.A2(n_1802),
.B1(n_1678),
.B2(n_1659),
.Y(n_1807)
);

AO22x2_ASAP7_75t_L g1808 ( 
.A1(n_1806),
.A2(n_1660),
.B1(n_1663),
.B2(n_1669),
.Y(n_1808)
);

NAND2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1807),
.B(n_1493),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1808),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1809),
.A2(n_1663),
.B(n_1660),
.Y(n_1811)
);

AND3x1_ASAP7_75t_L g1812 ( 
.A(n_1810),
.B(n_1811),
.C(n_1663),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1812),
.A2(n_1660),
.B(n_1490),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1813),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1673),
.B1(n_1670),
.B2(n_1669),
.C(n_1667),
.Y(n_1815)
);

AOI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1493),
.B(n_1670),
.C(n_1667),
.Y(n_1816)
);


endmodule