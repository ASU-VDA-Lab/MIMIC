module fake_netlist_6_983_n_104 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_104);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_104;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_63;
wire n_39;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVxp33_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_25),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_29),
.C(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_30),
.B1(n_27),
.B2(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_47),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_46),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_45),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_48),
.B1(n_53),
.B2(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AO21x2_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_59),
.B(n_57),
.Y(n_69)
);

AND2x4_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_62),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_62),
.Y(n_74)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_68),
.B(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_68),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_66),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_80),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_85),
.B(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_92),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_89),
.Y(n_94)
);

OAI311xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_85),
.A3(n_39),
.B1(n_66),
.C1(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_93),
.Y(n_96)
);

OAI221xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_94),
.B1(n_39),
.B2(n_65),
.C(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

OAI211xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_40),
.B(n_7),
.C(n_11),
.Y(n_99)
);

NAND5xp2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_6),
.C(n_12),
.D(n_15),
.E(n_69),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_69),
.C(n_70),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_100),
.B1(n_40),
.B2(n_49),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_40),
.B1(n_56),
.B2(n_101),
.Y(n_104)
);


endmodule