module fake_jpeg_14444_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g155 ( 
.A(n_61),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_68),
.B(n_77),
.Y(n_154)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_29),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_90),
.Y(n_119)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_94),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_96),
.Y(n_143)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_29),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_104),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_31),
.B(n_16),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_25),
.B1(n_34),
.B2(n_36),
.Y(n_152)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_103),
.A2(n_49),
.B1(n_38),
.B2(n_21),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_29),
.Y(n_104)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_58),
.A2(n_52),
.B1(n_32),
.B2(n_43),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_110),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_45),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_142),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_42),
.B1(n_43),
.B2(n_32),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_43),
.B1(n_42),
.B2(n_32),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_60),
.A2(n_63),
.B1(n_42),
.B2(n_49),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_70),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_64),
.A2(n_51),
.B1(n_50),
.B2(n_48),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_69),
.A2(n_51),
.B1(n_50),
.B2(n_48),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_126),
.B1(n_141),
.B2(n_149),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_34),
.B1(n_46),
.B2(n_36),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_22),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_54),
.A2(n_48),
.B1(n_22),
.B2(n_46),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_96),
.A2(n_66),
.B1(n_92),
.B2(n_73),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_55),
.A2(n_22),
.B1(n_46),
.B2(n_25),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_152),
.B(n_1),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_74),
.B(n_25),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_34),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_87),
.A2(n_36),
.B1(n_38),
.B2(n_47),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_47),
.B1(n_38),
.B2(n_19),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_81),
.B1(n_65),
.B2(n_91),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_163),
.A2(n_164),
.B1(n_194),
.B2(n_207),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_19),
.B1(n_21),
.B2(n_47),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_167),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_116),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_208),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_62),
.B1(n_91),
.B2(n_85),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_109),
.B(n_103),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_173),
.B(n_174),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_85),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_62),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_176),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_15),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_177),
.B(n_180),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_88),
.B1(n_61),
.B2(n_102),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_179),
.A2(n_158),
.A3(n_150),
.B1(n_129),
.B2(n_137),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_14),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_111),
.B(n_16),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_185),
.B(n_196),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_28),
.B(n_27),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_106),
.B(n_28),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_195),
.Y(n_218)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_106),
.B(n_28),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_143),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_27),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_114),
.B(n_16),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_197),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_112),
.B(n_26),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_199),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_26),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_115),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_212),
.B1(n_145),
.B2(n_157),
.Y(n_226)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

BUFx12_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_146),
.A2(n_23),
.B1(n_29),
.B2(n_2),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_124),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_213),
.Y(n_225)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_121),
.B(n_0),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_217),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_0),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_3),
.Y(n_228)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_148),
.B(n_3),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_184),
.A2(n_140),
.B1(n_129),
.B2(n_158),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_226),
.A2(n_232),
.B1(n_241),
.B2(n_254),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_228),
.B(n_246),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_169),
.A3(n_166),
.B1(n_165),
.B2(n_195),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_231),
.A2(n_248),
.B(n_175),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_157),
.B1(n_144),
.B2(n_145),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_169),
.B(n_161),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_236),
.B(n_239),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_161),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_178),
.A2(n_138),
.B1(n_142),
.B2(n_131),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_162),
.Y(n_246)
);

AOI32xp33_ASAP7_75t_L g248 ( 
.A1(n_184),
.A2(n_188),
.A3(n_198),
.B1(n_199),
.B2(n_211),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_SL g252 ( 
.A(n_176),
.B(n_124),
.C(n_162),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_252),
.B(n_133),
.Y(n_294)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_202),
.A2(n_138),
.B1(n_131),
.B2(n_137),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_172),
.A2(n_151),
.B1(n_108),
.B2(n_150),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_262),
.A2(n_182),
.B1(n_179),
.B2(n_130),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_192),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_206),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_171),
.A2(n_151),
.B1(n_108),
.B2(n_124),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_174),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_270),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_218),
.B(n_191),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_272),
.B(n_279),
.Y(n_324)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_174),
.C(n_176),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_285),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_248),
.A2(n_187),
.B1(n_163),
.B2(n_170),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_276),
.A2(n_281),
.B1(n_305),
.B2(n_259),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_278),
.A2(n_306),
.B(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_197),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_235),
.A2(n_191),
.B(n_194),
.C(n_179),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_289),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_247),
.A2(n_201),
.B1(n_179),
.B2(n_210),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_205),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_311),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_284),
.A2(n_302),
.B1(n_250),
.B2(n_219),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_215),
.C(n_167),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_225),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_295),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_298),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_190),
.C(n_189),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_234),
.A2(n_212),
.B(n_216),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_297),
.A2(n_312),
.B(n_230),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_218),
.B(n_133),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_227),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_300),
.Y(n_339)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_250),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_223),
.B(n_186),
.C(n_139),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_266),
.Y(n_342)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_247),
.A2(n_133),
.B1(n_193),
.B2(n_204),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_193),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_233),
.B(n_193),
.Y(n_307)
);

OAI211xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_252),
.B(n_245),
.C(n_223),
.Y(n_322)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_308),
.Y(n_352)
);

AO21x2_ASAP7_75t_L g309 ( 
.A1(n_244),
.A2(n_204),
.B(n_139),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_3),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_235),
.A2(n_139),
.B(n_5),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_315),
.A2(n_328),
.B(n_353),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_282),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_330),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_274),
.A2(n_234),
.B1(n_219),
.B2(n_264),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_321),
.A2(n_325),
.B1(n_329),
.B2(n_336),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_322),
.B(n_294),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_256),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_334),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_288),
.A2(n_231),
.B1(n_229),
.B2(n_245),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_268),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_283),
.A2(n_229),
.B1(n_241),
.B2(n_233),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_332),
.A2(n_306),
.B1(n_305),
.B2(n_298),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_272),
.B(n_287),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_293),
.A2(n_243),
.B(n_253),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_335),
.B(n_278),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_283),
.A2(n_237),
.B1(n_240),
.B2(n_266),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_351),
.C(n_333),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_276),
.A2(n_237),
.B1(n_240),
.B2(n_263),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_343),
.A2(n_346),
.B1(n_309),
.B2(n_310),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_281),
.A2(n_263),
.B1(n_238),
.B2(n_224),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_270),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_301),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_257),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_317),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_312),
.A2(n_243),
.B(n_238),
.Y(n_353)
);

INVx5_ASAP7_75t_SL g355 ( 
.A(n_330),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_355),
.A2(n_375),
.B1(n_385),
.B2(n_387),
.Y(n_420)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

AO22x2_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_309),
.B1(n_290),
.B2(n_280),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_366),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_351),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_371),
.C(n_377),
.Y(n_393)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_364),
.Y(n_409)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_316),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_353),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_369),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_320),
.B(n_309),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_370),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_314),
.B(n_309),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_372),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_339),
.B(n_289),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_379),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_352),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_376),
.A2(n_309),
.B(n_340),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_275),
.C(n_285),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_380),
.B1(n_381),
.B2(n_388),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_350),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_306),
.B1(n_274),
.B2(n_288),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_331),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_349),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_382),
.B(n_386),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_286),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_389),
.C(n_347),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_384),
.Y(n_391)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_271),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_352),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_314),
.B(n_295),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_390),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_327),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_402),
.C(n_412),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_380),
.A2(n_367),
.B1(n_328),
.B2(n_378),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_396),
.A2(n_379),
.B1(n_358),
.B2(n_355),
.Y(n_424)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_325),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_406),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_319),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_374),
.A2(n_315),
.B(n_336),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_404),
.A2(n_280),
.B(n_387),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_383),
.C(n_361),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_388),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_319),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_414),
.B(n_415),
.C(n_416),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_318),
.C(n_317),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_318),
.C(n_323),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_323),
.C(n_303),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_418),
.C(n_419),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_347),
.C(n_343),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_369),
.C(n_356),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_304),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_354),
.C(n_308),
.Y(n_446)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_422),
.Y(n_423)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_423),
.Y(n_450)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_424),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_391),
.A2(n_358),
.B1(n_375),
.B2(n_385),
.Y(n_425)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_425),
.Y(n_470)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_405),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_427),
.Y(n_452)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_400),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_429),
.B(n_435),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_391),
.A2(n_297),
.B1(n_358),
.B2(n_346),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_431),
.A2(n_415),
.B1(n_404),
.B2(n_413),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_395),
.A2(n_358),
.B1(n_364),
.B2(n_365),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_433),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_407),
.A2(n_418),
.B1(n_419),
.B2(n_397),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_412),
.B(n_271),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_434),
.B(n_447),
.Y(n_468)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_403),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_438),
.B(n_410),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_362),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_437),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_396),
.A2(n_357),
.B1(n_337),
.B2(n_341),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_441),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_341),
.B1(n_338),
.B2(n_337),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_442),
.Y(n_466)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_338),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_326),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_449),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_402),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_354),
.B1(n_292),
.B2(n_299),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_296),
.C(n_291),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_393),
.C(n_399),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_313),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_460),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_448),
.B(n_392),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_453),
.B(n_454),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_406),
.C(n_394),
.Y(n_454)
);

OAI22x1_ASAP7_75t_L g475 ( 
.A1(n_459),
.A2(n_424),
.B1(n_432),
.B2(n_425),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_269),
.Y(n_462)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_430),
.B(n_401),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_4),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_465),
.A2(n_4),
.B(n_5),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_398),
.C(n_224),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_469),
.C(n_460),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_269),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_446),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_445),
.B(n_260),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_471),
.B(n_443),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_475),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_465),
.A2(n_436),
.B(n_438),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_452),
.B(n_8),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_485),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_443),
.C(n_428),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_440),
.C(n_449),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_455),
.C(n_454),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_457),
.A2(n_444),
.B1(n_437),
.B2(n_442),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_479),
.A2(n_455),
.B1(n_470),
.B2(n_464),
.Y(n_492)
);

INVx11_ASAP7_75t_L g482 ( 
.A(n_450),
.Y(n_482)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_482),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_431),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_483),
.B(n_461),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_470),
.A2(n_260),
.B1(n_5),
.B2(n_6),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_484),
.A2(n_466),
.B1(n_458),
.B2(n_457),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_456),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_459),
.A2(n_6),
.B(n_7),
.Y(n_488)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_488),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_498),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_493),
.Y(n_505)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_492),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_451),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_499),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_466),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_456),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_502),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_501),
.A2(n_488),
.B(n_484),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_12),
.C(n_9),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_481),
.A2(n_479),
.B1(n_482),
.B2(n_486),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_504),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_498),
.Y(n_509)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_509),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_487),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_513),
.Y(n_524)
);

AOI31xp33_ASAP7_75t_L g512 ( 
.A1(n_494),
.A2(n_480),
.A3(n_477),
.B(n_473),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_496),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_491),
.A2(n_475),
.B(n_485),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_514),
.B(n_516),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_500),
.B(n_12),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_515),
.B(n_517),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_489),
.B(n_10),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_506),
.Y(n_518)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_518),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_499),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_523),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_511),
.B(n_489),
.Y(n_523)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_525),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_511),
.B(n_502),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_506),
.C(n_508),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_530),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_509),
.C(n_514),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_529),
.A2(n_524),
.B(n_520),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_532),
.A2(n_528),
.B1(n_495),
.B2(n_513),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_521),
.C(n_519),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_534),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_533),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_535),
.B(n_495),
.Y(n_538)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_11),
.B(n_530),
.Y(n_539)
);


endmodule