module real_jpeg_5505_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_61),
.B1(n_73),
.B2(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_1),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_1),
.A2(n_76),
.B1(n_208),
.B2(n_312),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_1),
.A2(n_76),
.B1(n_163),
.B2(n_164),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_1),
.A2(n_76),
.B1(n_331),
.B2(n_396),
.Y(n_395)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_2),
.Y(n_195)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_2),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_2),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_2),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_3),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_3),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_3),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_3),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_57),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_57),
.B1(n_143),
.B2(n_147),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_4),
.A2(n_57),
.B1(n_205),
.B2(n_380),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_5),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_5),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_5),
.A2(n_282),
.B1(n_360),
.B2(n_363),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_5),
.A2(n_282),
.B1(n_391),
.B2(n_394),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_L g446 ( 
.A1(n_5),
.A2(n_53),
.B1(n_282),
.B2(n_447),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_52),
.B1(n_61),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_64),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_6),
.A2(n_64),
.B1(n_281),
.B2(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_6),
.A2(n_64),
.B1(n_363),
.B2(n_406),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_50),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_7),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_7),
.A2(n_79),
.B1(n_222),
.B2(n_230),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_7),
.A2(n_79),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_7),
.A2(n_79),
.B1(n_431),
.B2(n_432),
.Y(n_430)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_8),
.Y(n_329)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_10),
.A2(n_169),
.B1(n_204),
.B2(n_208),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_10),
.A2(n_169),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_10),
.A2(n_169),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_11),
.Y(n_125)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_11),
.Y(n_178)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_13),
.Y(n_137)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_13),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_13),
.Y(n_198)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_14),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_15),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_15),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_15),
.A2(n_188),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_15),
.A2(n_188),
.B1(n_271),
.B2(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_15),
.A2(n_188),
.B1(n_399),
.B2(n_401),
.Y(n_398)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_17),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_17),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_17),
.B(n_178),
.C(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_17),
.B(n_91),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_17),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_17),
.B(n_172),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_17),
.B(n_266),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_18),
.A2(n_96),
.B1(n_163),
.B2(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_18),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_18),
.A2(n_214),
.B1(n_229),
.B2(n_234),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_18),
.A2(n_36),
.B1(n_214),
.B2(n_273),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_18),
.A2(n_43),
.B1(n_44),
.B2(n_214),
.Y(n_419)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_66),
.B(n_523),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_58),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_27),
.B(n_58),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_40),
.B(n_48),
.Y(n_27)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_28),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_28),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_29),
.B(n_165),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_29),
.A2(n_59),
.B1(n_398),
.B2(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_29)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_31),
.Y(n_263)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_32),
.Y(n_431)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_34),
.Y(n_393)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_34),
.Y(n_434)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_40),
.A2(n_347),
.B(n_349),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_40),
.B(n_351),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_45),
.Y(n_326)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_58)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_53),
.B(n_165),
.Y(n_335)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_58),
.B(n_68),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_65),
.B1(n_72),
.B2(n_77),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_77),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_59),
.A2(n_350),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_59),
.A2(n_65),
.B1(n_72),
.B2(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_65),
.A2(n_419),
.B(n_449),
.Y(n_459)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_152),
.B(n_522),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_148),
.C(n_149),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_69),
.A2(n_70),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_80),
.C(n_115),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_71),
.B(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_75),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_80),
.A2(n_115),
.B1(n_116),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_80),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_103),
.B1(n_110),
.B2(n_111),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_81),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_81),
.A2(n_110),
.B1(n_305),
.B2(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_81),
.A2(n_110),
.B1(n_390),
.B2(n_395),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_81),
.A2(n_103),
.B1(n_110),
.B2(n_499),
.Y(n_498)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_82)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_83),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_90),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_90),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_90),
.Y(n_357)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_91),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

AOI22x1_ASAP7_75t_L g420 ( 
.A1(n_91),
.A2(n_150),
.B1(n_307),
.B2(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_91),
.A2(n_150),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_94),
.Y(n_292)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g293 ( 
.A(n_96),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_96),
.Y(n_385)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_97),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_99),
.Y(n_362)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_99),
.Y(n_365)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_105),
.Y(n_272)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_109),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_110),
.B(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_110),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_112),
.Y(n_396)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_115),
.A2(n_116),
.B1(n_497),
.B2(n_498),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_115),
.B(n_494),
.C(n_497),
.Y(n_505)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_133),
.B(n_142),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_162),
.B(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_117),
.A2(n_133),
.B1(n_213),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_117),
.A2(n_166),
.B(n_256),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_117),
.A2(n_133),
.B1(n_359),
.B2(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_118),
.B(n_167),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_118),
.A2(n_172),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_118),
.A2(n_172),
.B1(n_384),
.B2(n_405),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_118),
.A2(n_172),
.B1(n_405),
.B2(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_133),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_123),
.B1(n_126),
.B2(n_130),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx5_ASAP7_75t_SL g291 ( 
.A(n_130),
.Y(n_291)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_133),
.A2(n_213),
.B(n_215),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_133),
.A2(n_215),
.B(n_359),
.Y(n_358)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_136),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_137),
.Y(n_381)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_142),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_147),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_148),
.B(n_149),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_150),
.A2(n_262),
.B(n_269),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_150),
.B(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_150),
.A2(n_269),
.B(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_516),
.B(n_521),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_488),
.B(n_513),
.Y(n_153)
);

OAI311xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_368),
.A3(n_464),
.B1(n_482),
.C1(n_483),
.Y(n_154)
);

AOI21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_318),
.B(n_367),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_296),
.B(n_317),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_250),
.B(n_295),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_218),
.B(n_249),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_181),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_160),
.B(n_181),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_173),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_161),
.A2(n_173),
.B1(n_174),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_165),
.A2(n_192),
.B(n_199),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g262 ( 
.A1(n_165),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_165),
.A2(n_335),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_210),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_211),
.C(n_217),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_192),
.B(n_199),
.Y(n_182)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_185),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_192),
.A2(n_201),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_192),
.A2(n_374),
.B1(n_377),
.B2(n_379),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_192),
.A2(n_201),
.B(n_379),
.Y(n_407)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_203),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_193),
.A2(n_279),
.B1(n_311),
.B2(n_314),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_193),
.A2(n_340),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_195),
.Y(n_315)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_198),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_228),
.B(n_237),
.Y(n_227)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_240),
.B(n_248),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_226),
.B(n_239),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_238),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_238),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_237),
.A2(n_278),
.B(n_285),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_246),
.Y(n_248)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_252),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_276),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_260),
.B2(n_261),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_260),
.C(n_276),
.Y(n_297)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_259),
.Y(n_387)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_289),
.A3(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_275),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_288),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_287),
.Y(n_378)
);

INVx4_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_297),
.B(n_298),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_316),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_302),
.C(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_309),
.C(n_310),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_319),
.B(n_320),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_344),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_321)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_336),
.B2(n_337),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_324),
.B(n_336),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.A3(n_327),
.B1(n_330),
.B2(n_335),
.Y(n_324)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_341),
.B(n_343),
.C(n_344),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_354),
.B2(n_366),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_345),
.B(n_355),
.C(n_358),
.Y(n_473)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_356),
.Y(n_462)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_450),
.Y(n_368)
);

A2O1A1Ixp33_ASAP7_75t_SL g483 ( 
.A1(n_369),
.A2(n_450),
.B(n_484),
.C(n_487),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_422),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_370),
.B(n_422),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_402),
.C(n_409),
.Y(n_370)
);

FAx1_ASAP7_75t_SL g463 ( 
.A(n_371),
.B(n_402),
.CI(n_409),
.CON(n_463),
.SN(n_463)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_388),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_372),
.B(n_389),
.C(n_397),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_382),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_373),
.B(n_382),
.Y(n_456)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_374),
.Y(n_414)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_383),
.Y(n_412)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_397),
.Y(n_388)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_390),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx6_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_407),
.B2(n_408),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_407),
.A2(n_408),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_407),
.A2(n_441),
.B(n_444),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_417),
.C(n_420),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_411),
.B(n_413),
.Y(n_472)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_417),
.A2(n_418),
.B1(n_420),
.B2(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_420),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_423),
.B(n_426),
.C(n_439),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_439),
.B2(n_440),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_435),
.B(n_438),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_436),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_430),
.Y(n_499)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_438),
.B(n_491),
.CI(n_492),
.CON(n_490),
.SN(n_490)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_438),
.B(n_491),
.C(n_492),
.Y(n_512)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_449),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_446),
.Y(n_495)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_463),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_451),
.B(n_463),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_456),
.C(n_457),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_452),
.A2(n_453),
.B1(n_456),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_456),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_475),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.C(n_461),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_458),
.A2(n_459),
.B1(n_461),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_460),
.B(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_463),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_477),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_485),
.B(n_486),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_474),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_474),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_471),
.C(n_473),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_480),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_471),
.A2(n_472),
.B1(n_473),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_479),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_502),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_501),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_501),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_490),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B1(n_496),
.B2(n_500),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_494),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_504),
.C(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_496),
.Y(n_500)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_512),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_512),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_520),
.Y(n_521)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);


endmodule