module fake_jpeg_14876_n_122 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx5_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_35),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_10),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_16),
.B(n_12),
.C(n_11),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_51),
.B1(n_31),
.B2(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_26),
.B1(n_21),
.B2(n_25),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_64),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_43),
.B1(n_38),
.B2(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_63),
.B1(n_49),
.B2(n_52),
.Y(n_69)
);

AOI22x1_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_36),
.B1(n_40),
.B2(n_31),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_61),
.B1(n_21),
.B2(n_26),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_31),
.B1(n_43),
.B2(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_70),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_44),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_51),
.B(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_21),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_30),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_65),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_79),
.B(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_85),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_22),
.C(n_28),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_28),
.C(n_22),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_86),
.B(n_80),
.CI(n_76),
.CON(n_87),
.SN(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_9),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_71),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_90),
.C(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_3),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_22),
.C(n_28),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_4),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_92),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_82),
.B1(n_84),
.B2(n_29),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_23),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_87),
.B1(n_94),
.B2(n_23),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_87),
.B1(n_23),
.B2(n_12),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_11),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_96),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.C(n_113),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_4),
.B(n_7),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_8),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_9),
.B(n_7),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_115),
.C(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_119),
.B(n_4),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_121),
.Y(n_122)
);


endmodule