module fake_jpeg_31947_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_15),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_56),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_27),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_76),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_18),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_75),
.B(n_93),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_27),
.B(n_0),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_28),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_1),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_100),
.Y(n_139)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_28),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_104),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_40),
.B1(n_19),
.B2(n_42),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_106),
.A2(n_154),
.B1(n_88),
.B2(n_104),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_20),
.B(n_39),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_125),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_30),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_87),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_30),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_122),
.B(n_158),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_35),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_35),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_156),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_72),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_100),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_98),
.A2(n_103),
.B1(n_101),
.B2(n_97),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_138),
.A2(n_160),
.B1(n_43),
.B2(n_2),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_40),
.B1(n_19),
.B2(n_42),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_78),
.B(n_37),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_94),
.B(n_37),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_54),
.A2(n_36),
.B1(n_50),
.B2(n_25),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_117),
.A2(n_67),
.B1(n_89),
.B2(n_60),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_118),
.A2(n_63),
.B1(n_57),
.B2(n_65),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_175),
.A2(n_9),
.B(n_11),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_106),
.A2(n_61),
.B1(n_81),
.B2(n_79),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_186),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_133),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_197),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_39),
.B(n_20),
.C(n_44),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_181),
.A2(n_215),
.B(n_9),
.C(n_10),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_162),
.B1(n_147),
.B2(n_165),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_41),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_191),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_112),
.B(n_41),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_188),
.B(n_194),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_189),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_44),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_131),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_68),
.B1(n_74),
.B2(n_73),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_196),
.B(n_200),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_107),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_71),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_164),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_147),
.A2(n_50),
.B1(n_42),
.B2(n_25),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_201),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_51),
.B1(n_50),
.B2(n_53),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_202),
.A2(n_203),
.B1(n_217),
.B2(n_221),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_120),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_129),
.A2(n_51),
.B1(n_43),
.B2(n_34),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_204),
.A2(n_218),
.B1(n_144),
.B2(n_130),
.Y(n_259)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_205),
.B(n_208),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_108),
.A2(n_43),
.B1(n_2),
.B2(n_4),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_213),
.B1(n_216),
.B2(n_220),
.Y(n_232)
);

CKINVDCx6p67_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_210),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_145),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_123),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_108),
.A2(n_164),
.B1(n_126),
.B2(n_148),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_214),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_215)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_143),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_157),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g237 ( 
.A(n_219),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_126),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_120),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

CKINVDCx12_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_159),
.B(n_6),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_226),
.B(n_247),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_231),
.B(n_235),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_148),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_195),
.A2(n_177),
.B1(n_216),
.B2(n_204),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_242),
.A2(n_264),
.B1(n_263),
.B2(n_225),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_167),
.B(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_251),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_185),
.B(n_153),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_144),
.Y(n_251)
);

OR2x2_ASAP7_75t_SL g253 ( 
.A(n_171),
.B(n_150),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_207),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_258),
.B(n_220),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_259),
.A2(n_189),
.B1(n_176),
.B2(n_193),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_130),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_262),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_198),
.B(n_110),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_173),
.A2(n_115),
.B1(n_114),
.B2(n_113),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_196),
.B(n_115),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_261),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_196),
.B(n_9),
.CI(n_11),
.CON(n_269),
.SN(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_180),
.B(n_219),
.C(n_208),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_207),
.B(n_11),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_179),
.A2(n_181),
.B1(n_215),
.B2(n_178),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_218),
.B1(n_197),
.B2(n_170),
.Y(n_277)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_237),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_288),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_277),
.Y(n_349)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_166),
.B(n_194),
.C(n_186),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_279),
.A2(n_280),
.B(n_285),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_266),
.A2(n_253),
.B(n_243),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_183),
.B1(n_187),
.B2(n_207),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_282),
.B(n_287),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_222),
.B1(n_210),
.B2(n_183),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_283),
.A2(n_306),
.B1(n_239),
.B2(n_255),
.Y(n_339)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_286),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_246),
.B(n_205),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_232),
.A2(n_192),
.B1(n_184),
.B2(n_169),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_289),
.A2(n_305),
.B1(n_311),
.B2(n_225),
.Y(n_323)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_189),
.B(n_190),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_298),
.B(n_303),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_293),
.B(n_295),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_248),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_294),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_251),
.B(n_201),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_300),
.B1(n_308),
.B2(n_314),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_238),
.A2(n_211),
.B(n_217),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_248),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_128),
.B1(n_150),
.B2(n_200),
.Y(n_300)
);

BUFx24_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_301),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_235),
.B(n_209),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_302),
.B(n_307),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_233),
.A2(n_214),
.B1(n_176),
.B2(n_13),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_244),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_244),
.A2(n_17),
.B1(n_13),
.B2(n_14),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_233),
.A2(n_13),
.B(n_14),
.C(n_17),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_259),
.A2(n_14),
.B1(n_231),
.B2(n_264),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_265),
.A2(n_225),
.B1(n_263),
.B2(n_270),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_310),
.A2(n_245),
.B1(n_241),
.B2(n_256),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_14),
.B1(n_262),
.B2(n_230),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_229),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_258),
.B(n_226),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_313),
.B(n_250),
.Y(n_341)
);

O2A1O1Ixp33_ASAP7_75t_SL g314 ( 
.A1(n_255),
.A2(n_269),
.B(n_257),
.C(n_225),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_245),
.B1(n_260),
.B2(n_256),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_274),
.B(n_269),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_321),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_323),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_229),
.B1(n_228),
.B2(n_227),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_297),
.Y(n_381)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_274),
.B(n_273),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_334),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_267),
.C(n_254),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_343),
.C(n_356),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_254),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_338),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_340),
.Y(n_363)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_282),
.A2(n_228),
.A3(n_240),
.B1(n_245),
.B2(n_227),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_341),
.B(n_344),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_240),
.C(n_241),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_250),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_347),
.Y(n_358)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_350),
.A2(n_289),
.B1(n_302),
.B2(n_295),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_294),
.B(n_260),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_354),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_285),
.B(n_303),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_284),
.B(n_239),
.C(n_287),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_359),
.A2(n_371),
.B1(n_379),
.B2(n_324),
.Y(n_416)
);

AO22x1_ASAP7_75t_L g361 ( 
.A1(n_326),
.A2(n_279),
.B1(n_280),
.B2(n_312),
.Y(n_361)
);

AO21x2_ASAP7_75t_SL g411 ( 
.A1(n_361),
.A2(n_329),
.B(n_357),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_364),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_352),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_365),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_284),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_370),
.C(n_382),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_288),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_325),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_345),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_332),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_288),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_342),
.A2(n_309),
.B1(n_308),
.B2(n_313),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_298),
.B(n_292),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_372),
.A2(n_318),
.B(n_330),
.Y(n_398)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_374),
.Y(n_407)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_320),
.Y(n_378)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_378),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_342),
.A2(n_309),
.B1(n_299),
.B2(n_317),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_320),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_381),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_316),
.C(n_291),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_352),
.B(n_323),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_307),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_384),
.Y(n_394)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_388),
.Y(n_401)
);

O2A1O1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_318),
.A2(n_314),
.B(n_290),
.C(n_293),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_392),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_314),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_343),
.C(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

BUFx8_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_393),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_386),
.A2(n_349),
.B1(n_332),
.B2(n_334),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_395),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_384),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_396),
.B(n_397),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_SL g451 ( 
.A(n_398),
.B(n_417),
.C(n_301),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_356),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_404),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_384),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_405),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_357),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_408),
.B(n_419),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_361),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_373),
.Y(n_450)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_411),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_409),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_362),
.A2(n_363),
.B1(n_381),
.B2(n_365),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_413),
.A2(n_371),
.B1(n_359),
.B2(n_389),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_322),
.C(n_333),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_366),
.C(n_367),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_416),
.A2(n_423),
.B1(n_380),
.B2(n_378),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_372),
.A2(n_388),
.B(n_360),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_376),
.A2(n_330),
.B1(n_350),
.B2(n_355),
.Y(n_418)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_382),
.B(n_321),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_422),
.A2(n_424),
.B(n_390),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_379),
.A2(n_340),
.B1(n_346),
.B2(n_345),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_383),
.A2(n_337),
.B(n_348),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_426),
.A2(n_428),
.B1(n_450),
.B2(n_394),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_422),
.A2(n_391),
.B1(n_362),
.B2(n_367),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_429),
.A2(n_448),
.B(n_451),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_435),
.Y(n_465)
);

NOR3xp33_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_301),
.C(n_387),
.Y(n_431)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_431),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_351),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_433),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_351),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_434),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_392),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_441),
.C(n_415),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_438),
.A2(n_413),
.B1(n_402),
.B2(n_396),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_375),
.C(n_374),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_394),
.B(n_373),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_443),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_404),
.B(n_276),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_446),
.Y(n_461)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_401),
.A2(n_402),
.B(n_424),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_403),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_428),
.B(n_412),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_455),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_459),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_454),
.A2(n_439),
.B1(n_445),
.B2(n_447),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_430),
.B(n_417),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_440),
.B(n_393),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_468),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_406),
.C(n_423),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_462),
.C(n_463),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_425),
.B(n_429),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_435),
.C(n_436),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_406),
.C(n_416),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_398),
.C(n_397),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_471),
.C(n_472),
.Y(n_485)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_467),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_397),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_426),
.B(n_401),
.Y(n_472)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_427),
.C(n_450),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_459),
.Y(n_497)
);

BUFx24_ASAP7_75t_SL g476 ( 
.A(n_460),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_455),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_439),
.B1(n_438),
.B2(n_427),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_477),
.A2(n_483),
.B1(n_486),
.B2(n_369),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_471),
.B1(n_411),
.B2(n_461),
.Y(n_496)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_472),
.A2(n_445),
.B1(n_446),
.B2(n_443),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_473),
.A2(n_447),
.B1(n_400),
.B2(n_442),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_487),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_469),
.A2(n_449),
.B1(n_411),
.B2(n_393),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_400),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_465),
.C(n_453),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_489),
.B(n_465),
.C(n_452),
.Y(n_492)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_464),
.Y(n_490)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_490),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_492),
.B(n_500),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_479),
.A2(n_454),
.B1(n_458),
.B2(n_463),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_498),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_475),
.A2(n_469),
.B(n_466),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_495),
.A2(n_488),
.B(n_482),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_497),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_486),
.A2(n_432),
.B1(n_411),
.B2(n_421),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_503),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_474),
.A2(n_421),
.B1(n_420),
.B2(n_405),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_483),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_432),
.C(n_420),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_504),
.C(n_481),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_488),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_477),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_358),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_492),
.A2(n_481),
.B(n_485),
.Y(n_510)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_511),
.A2(n_495),
.B(n_497),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_515),
.C(n_517),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_482),
.C(n_369),
.Y(n_515)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_516),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_358),
.C(n_328),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_505),
.A2(n_496),
.B(n_501),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_513),
.B(n_505),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_521),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_508),
.A2(n_506),
.B1(n_493),
.B2(n_491),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_525),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_514),
.B(n_500),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_515),
.B(n_503),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_517),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_509),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_530),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_507),
.C(n_509),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_531),
.Y(n_532)
);

MAJx2_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_522),
.C(n_529),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_527),
.C(n_520),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_527),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_535),
.B(n_536),
.C(n_532),
.Y(n_537)
);

AOI322xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_524),
.A3(n_512),
.B1(n_346),
.B2(n_335),
.C1(n_337),
.C2(n_331),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_538),
.B(n_331),
.Y(n_539)
);

AOI21xp33_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_335),
.B(n_347),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_354),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_239),
.C(n_301),
.Y(n_542)
);


endmodule