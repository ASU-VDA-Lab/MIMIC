module real_jpeg_17620_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_522),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_0),
.B(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_1),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_1),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_1),
.A2(n_12),
.B1(n_259),
.B2(n_262),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_1),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_1),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_1),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_1),
.B(n_426),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_1),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_1),
.B(n_377),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_2),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_2),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_2),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_2),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_2),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_2),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_2),
.B(n_485),
.Y(n_484)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_3),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_3),
.Y(n_261)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_3),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_5),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_5),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_5),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_5),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_5),
.B(n_377),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_6),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_6),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_6),
.B(n_230),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_8),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_8),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_9),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_9),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_9),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_9),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_9),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_9),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_9),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_9),
.B(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_10),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_10),
.Y(n_236)
);

BUFx4f_ASAP7_75t_L g441 ( 
.A(n_10),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_11),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_12),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_12),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_12),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_12),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_12),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_12),
.B(n_87),
.Y(n_237)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_12),
.Y(n_375)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_14),
.Y(n_131)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_14),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_14),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_15),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_15),
.B(n_91),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_15),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_15),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_15),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_15),
.B(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_16),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_16),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_16),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_16),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_16),
.B(n_381),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_16),
.B(n_329),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_18),
.Y(n_139)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_198),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_197),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_161),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_24),
.B(n_161),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_108),
.C(n_122),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_25),
.A2(n_26),
.B1(n_108),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_66),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_48),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_28),
.B(n_48),
.C(n_163),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_42),
.C(n_44),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_29),
.A2(n_30),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.C(n_38),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_31),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_31),
.A2(n_36),
.B1(n_79),
.B2(n_157),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_35),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_36),
.B(n_146),
.C(n_149),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_36),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_36),
.A2(n_149),
.B1(n_157),
.B2(n_224),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g377 ( 
.A(n_37),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_38),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_38),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_38),
.A2(n_154),
.B1(n_269),
.B2(n_321),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_42),
.B(n_44),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_42),
.B(n_229),
.C(n_233),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_42),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_44),
.Y(n_140)
);

OAI22x1_ASAP7_75t_SL g243 ( 
.A1(n_44),
.A2(n_137),
.B1(n_140),
.B2(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_47),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_47),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g407 ( 
.A(n_47),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_49),
.B(n_53),
.C(n_65),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_51),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_60),
.B2(n_65),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_59),
.Y(n_335)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_64),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_80),
.C(n_95),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_67),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_76),
.C(n_79),
.Y(n_120)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_73),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_76),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_SL g170 ( 
.A(n_76),
.B(n_111),
.C(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_78),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_80),
.B(n_95),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.C(n_90),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_90),
.Y(n_144)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2x2_ASAP7_75t_SL g143 ( 
.A(n_86),
.B(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_88),
.Y(n_337)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_93),
.Y(n_424)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_100),
.C(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_108),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_120),
.C(n_121),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_111),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_111),
.A2(n_113),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_112),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_122),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_141),
.C(n_158),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_123),
.B(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_137),
.C(n_140),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_124),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_132),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_125),
.B(n_132),
.Y(n_226)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_127),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_128),
.B(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_136),
.Y(n_268)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_139),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_142),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_153),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_143),
.B(n_145),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_146),
.B(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_149),
.Y(n_224)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_152),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_153),
.B(n_305),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_154),
.B(n_265),
.C(n_269),
.Y(n_264)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_183),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_180),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_196),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_519),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_248),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_245),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_202),
.B(n_245),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.C(n_208),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_203),
.B(n_205),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_208),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_227),
.C(n_242),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_210),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_222),
.C(n_225),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_211),
.B(n_222),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.C(n_219),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_212),
.A2(n_219),
.B1(n_220),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_212),
.Y(n_346)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_215),
.B(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_219),
.B(n_402),
.C(n_406),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_219),
.A2(n_220),
.B1(n_406),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2x2_ASAP7_75t_SL g313 ( 
.A(n_225),
.B(n_314),
.Y(n_313)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_242),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_237),
.C(n_238),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_233),
.Y(n_256)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_236),
.Y(n_382)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_236),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_238),
.A2(n_239),
.B1(n_384),
.B2(n_385),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_239),
.B(n_379),
.C(n_384),
.Y(n_378)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AO21x2_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_353),
.B(n_516),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_347),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_308),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_251),
.B(n_308),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_301),
.Y(n_251)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_252),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_272),
.C(n_296),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_254),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.C(n_264),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_255),
.B(n_389),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_257),
.A2(n_258),
.B1(n_264),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_258),
.A2(n_369),
.B(n_374),
.Y(n_368)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_264),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_273),
.A2(n_297),
.B1(n_298),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_287),
.C(n_291),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_274),
.B(n_343),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_281),
.C(n_283),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_275),
.A2(n_283),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_275),
.Y(n_367)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_277),
.Y(n_457)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_280),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_281),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_283),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_283),
.B(n_422),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2x1_ASAP7_75t_L g343 ( 
.A(n_288),
.B(n_291),
.Y(n_343)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_351),
.C(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.C(n_315),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_309),
.A2(n_310),
.B1(n_313),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_342),
.C(n_344),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_317),
.B(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_322),
.C(n_332),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2x2_ASAP7_75t_L g410 ( 
.A(n_319),
.B(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_322),
.B(n_332),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_323),
.B(n_328),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_331),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.C(n_338),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_333),
.A2(n_336),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_336),
.A2(n_399),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_336),
.B(n_462),
.C(n_466),
.Y(n_493)
);

XOR2x2_ASAP7_75t_SL g396 ( 
.A(n_338),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_344),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_347),
.A2(n_517),
.B(n_518),
.Y(n_516)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_348),
.B(n_350),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_414),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.C(n_391),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_356),
.B(n_360),
.Y(n_515)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.C(n_387),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_388),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.C(n_378),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_368),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_366),
.B(n_423),
.C(n_425),
.Y(n_447)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_379),
.B(n_502),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_383),
.Y(n_454)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_380),
.A2(n_471),
.B1(n_472),
.B2(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_412),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_412),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_410),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_393),
.B(n_513),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_395),
.B(n_410),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_400),
.C(n_408),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_396),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_401),
.B(n_409),
.Y(n_507)
);

XOR2x2_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_406),
.Y(n_450)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_416),
.C(n_515),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_510),
.B(n_514),
.Y(n_416)
);

AOI21x1_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_496),
.B(n_509),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_458),
.B(n_495),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_445),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_420),
.B(n_445),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_428),
.C(n_437),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_421),
.B(n_491),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_425),
.Y(n_422)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_428),
.A2(n_429),
.B1(n_437),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_430),
.B(n_433),
.Y(n_463)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx6_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

AO22x1_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_442),
.B1(n_443),
.B2(n_444),
.Y(n_437)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_438),
.Y(n_443)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_442),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_443),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_484),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_451),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_447),
.B(n_448),
.C(n_451),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g504 ( 
.A(n_452),
.B(n_454),
.C(n_455),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_489),
.B(n_494),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_460),
.A2(n_473),
.B(n_488),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_470),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_470),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_472),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_483),
.B(n_487),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_481),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_481),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_493),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_SL g494 ( 
.A(n_490),
.B(n_493),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_508),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_497),
.B(n_508),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_499),
.B1(n_505),
.B2(n_506),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_503),
.B2(n_504),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_504),
.C(n_505),
.Y(n_511)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_512),
.Y(n_514)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);


endmodule