module fake_aes_8792_n_1395 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1395);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1395;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1390;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g318 ( .A(n_151), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_114), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_211), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_11), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_206), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_255), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_79), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_246), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_171), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_209), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_149), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_104), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_93), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_254), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_7), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_145), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_132), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_105), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_216), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_56), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_189), .Y(n_338) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_224), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_22), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_160), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_71), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_270), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_275), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_8), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_48), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_79), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_87), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_277), .Y(n_349) );
CKINVDCx14_ASAP7_75t_R g350 ( .A(n_207), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_219), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_205), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_118), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_247), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_74), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_187), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_282), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_38), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_308), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_248), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_41), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_287), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_36), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_43), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_200), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_62), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_143), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_6), .Y(n_368) );
INVxp33_ASAP7_75t_L g369 ( .A(n_122), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_84), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_123), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_299), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_115), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_176), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_263), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_5), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_227), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_288), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_226), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_44), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_190), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_34), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_193), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_61), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_24), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_95), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_113), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_310), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_42), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_126), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_97), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_197), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_273), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_291), .Y(n_394) );
INVxp33_ASAP7_75t_SL g395 ( .A(n_180), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_159), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_238), .Y(n_397) );
BUFx10_ASAP7_75t_L g398 ( .A(n_218), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_6), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_182), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_249), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_42), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_144), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_298), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_292), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_136), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_174), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_161), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_243), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_139), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_317), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_124), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_24), .Y(n_413) );
INVxp33_ASAP7_75t_L g414 ( .A(n_293), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_306), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_157), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_181), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_281), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_36), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_212), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_245), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_272), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_262), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_295), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_175), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_121), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_204), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_186), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_9), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_37), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_146), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_210), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_81), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_251), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_313), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_130), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_239), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_73), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_168), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_92), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_135), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_236), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_316), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_45), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_229), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_127), .Y(n_446) );
INVxp33_ASAP7_75t_L g447 ( .A(n_134), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_221), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_274), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_110), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_25), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_280), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_208), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_8), .Y(n_454) );
INVxp33_ASAP7_75t_SL g455 ( .A(n_279), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_244), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_39), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_55), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_88), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_233), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_294), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_39), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_158), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_286), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_109), .Y(n_465) );
INVxp33_ASAP7_75t_SL g466 ( .A(n_258), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_297), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_78), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_108), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_9), .Y(n_470) );
BUFx5_ASAP7_75t_L g471 ( .A(n_223), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_259), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_22), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_164), .B(n_152), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_194), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_203), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_68), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_260), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_267), .Y(n_479) );
INVxp33_ASAP7_75t_L g480 ( .A(n_234), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_369), .B(n_0), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_340), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_411), .B(n_0), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_382), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_471), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_369), .B(n_1), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_382), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_340), .B(n_1), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_389), .B(n_2), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_389), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_429), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_429), .B(n_2), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_471), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_318), .Y(n_494) );
NOR2xp33_ASAP7_75t_SL g495 ( .A(n_330), .B(n_86), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_471), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_319), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_322), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_411), .B(n_3), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_423), .B(n_3), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_471), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_471), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_323), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_328), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_329), .Y(n_506) );
BUFx12f_ASAP7_75t_L g507 ( .A(n_398), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_471), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_342), .B(n_4), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_331), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_423), .B(n_4), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_334), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_451), .B(n_327), .Y(n_513) );
BUFx12f_ASAP7_75t_L g514 ( .A(n_398), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_326), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_326), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_376), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_326), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_335), .Y(n_519) );
BUFx3_ASAP7_75t_L g520 ( .A(n_500), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_515), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_507), .B(n_391), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_482), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_507), .B(n_409), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_485), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_507), .B(n_418), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_485), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_514), .Y(n_529) );
INVx5_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
NAND2xp33_ASAP7_75t_L g531 ( .A(n_481), .B(n_320), .Y(n_531) );
NOR2x1p5_ASAP7_75t_L g532 ( .A(n_514), .B(n_364), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_493), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
NAND3x1_ASAP7_75t_L g535 ( .A(n_513), .B(n_332), .C(n_321), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_493), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_496), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_496), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_515), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_489), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_515), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_500), .B(n_469), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_496), .Y(n_543) );
AND3x2_ASAP7_75t_L g544 ( .A(n_495), .B(n_363), .C(n_358), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_499), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_482), .B(n_414), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_494), .B(n_414), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_481), .A2(n_354), .B1(n_403), .B2(n_401), .Y(n_549) );
INVx4_ASAP7_75t_L g550 ( .A(n_500), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_494), .B(n_497), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_500), .Y(n_552) );
BUFx3_ASAP7_75t_L g553 ( .A(n_501), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_515), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_497), .B(n_447), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_498), .B(n_447), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g558 ( .A(n_514), .B(n_436), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_489), .A2(n_337), .B1(n_346), .B2(n_345), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_501), .B(n_475), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_517), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_501), .B(n_347), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_498), .B(n_480), .Y(n_564) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_516), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_504), .B(n_480), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_499), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_502), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_548), .B(n_486), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_520), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_563), .A2(n_511), .B(n_501), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_559), .A2(n_354), .B1(n_403), .B2(n_401), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_556), .B(n_557), .Y(n_573) );
OR2x6_ASAP7_75t_L g574 ( .A(n_549), .B(n_486), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_532), .B(n_511), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_523), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_540), .A2(n_492), .B1(n_489), .B2(n_488), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_540), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_540), .Y(n_579) );
INVx5_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
INVxp33_ASAP7_75t_L g581 ( .A(n_546), .Y(n_581) );
INVx4_ASAP7_75t_L g582 ( .A(n_550), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g583 ( .A1(n_561), .A2(n_430), .B1(n_468), .B2(n_376), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_550), .B(n_511), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_542), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_555), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_555), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_520), .Y(n_588) );
NAND2xp33_ASAP7_75t_SL g589 ( .A(n_532), .B(n_511), .Y(n_589) );
INVx5_ASAP7_75t_L g590 ( .A(n_555), .Y(n_590) );
INVx6_ASAP7_75t_L g591 ( .A(n_563), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_564), .B(n_504), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_529), .B(n_509), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_566), .B(n_505), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_523), .B(n_488), .Y(n_595) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_558), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_563), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_542), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_542), .B(n_505), .Y(n_599) );
AND2x4_ASAP7_75t_SL g600 ( .A(n_542), .B(n_430), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_552), .A2(n_492), .B1(n_488), .B2(n_506), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_528), .A2(n_503), .B(n_502), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_563), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_551), .Y(n_604) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_552), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_560), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_553), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_560), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_560), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_560), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_565), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_535), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_528), .B(n_492), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_535), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_531), .B(n_506), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_533), .B(n_492), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_533), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_527), .B(n_510), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_SL g619 ( .A1(n_524), .A2(n_483), .B(n_350), .C(n_502), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_522), .B(n_355), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_534), .B(n_510), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_536), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_536), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_526), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_537), .B(n_512), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_544), .Y(n_626) );
OAI22xp5_ASAP7_75t_SL g627 ( .A1(n_525), .A2(n_477), .B1(n_468), .B2(n_364), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_537), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_538), .B(n_512), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_538), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_543), .B(n_419), .C(n_413), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_543), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_545), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_545), .Y(n_634) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_547), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_547), .B(n_519), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_526), .B(n_413), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_567), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_567), .A2(n_433), .B1(n_444), .B2(n_419), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_568), .Y(n_640) );
AO22x1_ASAP7_75t_L g641 ( .A1(n_530), .A2(n_455), .B1(n_466), .B2(n_395), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_530), .B(n_484), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_565), .B(n_503), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_565), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_565), .Y(n_645) );
NAND2xp33_ASAP7_75t_SL g646 ( .A(n_521), .B(n_333), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_521), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_530), .A2(n_508), .B(n_503), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_530), .B(n_508), .Y(n_649) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_521), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_530), .B(n_508), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_530), .A2(n_487), .B1(n_490), .B2(n_484), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_539), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_539), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_539), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_539), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_521), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_642), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_580), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_633), .Y(n_660) );
INVx3_ASAP7_75t_L g661 ( .A(n_580), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_SL g662 ( .A1(n_619), .A2(n_474), .B(n_336), .C(n_341), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_581), .B(n_395), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_580), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_635), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_604), .Y(n_666) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_580), .Y(n_667) );
INVx2_ASAP7_75t_SL g668 ( .A(n_600), .Y(n_668) );
OAI22xp5_ASAP7_75t_SL g669 ( .A1(n_583), .A2(n_477), .B1(n_444), .B2(n_366), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_582), .Y(n_670) );
NAND2xp33_ASAP7_75t_R g671 ( .A(n_574), .B(n_455), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_582), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_597), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_584), .A2(n_374), .B(n_339), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_590), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_603), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_596), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_572), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_609), .B(n_361), .Y(n_679) );
OR2x6_ASAP7_75t_L g680 ( .A(n_574), .B(n_368), .Y(n_680) );
BUFx2_ASAP7_75t_L g681 ( .A(n_574), .Y(n_681) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_570), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_573), .B(n_466), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_581), .B(n_385), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_585), .B(n_598), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_571), .A2(n_343), .B(n_338), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_593), .B(n_324), .Y(n_687) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_570), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_569), .B(n_384), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_621), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_590), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_610), .B(n_637), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_576), .Y(n_693) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_570), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_625), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_590), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_629), .Y(n_697) );
AO21x2_ASAP7_75t_L g698 ( .A1(n_619), .A2(n_348), .B(n_344), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_636), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_577), .A2(n_380), .B1(n_402), .B2(n_399), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_570), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_575), .Y(n_702) );
BUFx12f_ASAP7_75t_L g703 ( .A(n_626), .Y(n_703) );
BUFx12f_ASAP7_75t_L g704 ( .A(n_620), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_577), .A2(n_438), .B1(n_457), .B2(n_454), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_610), .B(n_370), .Y(n_706) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_642), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_615), .B(n_490), .C(n_487), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_606), .B(n_458), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_590), .Y(n_710) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_591), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_591), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_591), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_608), .A2(n_350), .B1(n_470), .B2(n_462), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_578), .Y(n_715) );
NAND2x1p5_ASAP7_75t_L g716 ( .A(n_640), .B(n_491), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_627), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_571), .A2(n_473), .B(n_491), .C(n_352), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_599), .B(n_333), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_639), .B(n_349), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_632), .B(n_349), .Y(n_721) );
BUFx3_ASAP7_75t_L g722 ( .A(n_653), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_607), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_632), .B(n_407), .Y(n_724) );
BUFx3_ASAP7_75t_L g725 ( .A(n_620), .Y(n_725) );
INVx5_ASAP7_75t_L g726 ( .A(n_607), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_595), .Y(n_727) );
INVx3_ASAP7_75t_L g728 ( .A(n_588), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_592), .A2(n_356), .B(n_351), .Y(n_729) );
BUFx4f_ASAP7_75t_L g730 ( .A(n_575), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_594), .B(n_407), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_615), .B(n_408), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_617), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_579), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g735 ( .A1(n_601), .A2(n_359), .B(n_360), .C(n_357), .Y(n_735) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_611), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_589), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_605), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_601), .B(n_408), .Y(n_739) );
BUFx4f_ASAP7_75t_SL g740 ( .A(n_612), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_614), .B(n_410), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_622), .B(n_412), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_623), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_595), .B(n_362), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_605), .B(n_425), .Y(n_745) );
BUFx8_ASAP7_75t_L g746 ( .A(n_655), .Y(n_746) );
O2A1O1Ixp33_ASAP7_75t_L g747 ( .A1(n_613), .A2(n_371), .B(n_373), .C(n_365), .Y(n_747) );
BUFx3_ASAP7_75t_L g748 ( .A(n_656), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_586), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_628), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_618), .B(n_425), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_630), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_631), .A2(n_398), .B1(n_378), .B2(n_386), .Y(n_753) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_587), .A2(n_434), .B1(n_441), .B2(n_428), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_634), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_641), .B(n_428), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_638), .B(n_434), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_613), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_616), .A2(n_387), .B1(n_390), .B2(n_377), .Y(n_759) );
O2A1O1Ixp5_ASAP7_75t_L g760 ( .A1(n_616), .A2(n_375), .B(n_388), .C(n_367), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_611), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_624), .A2(n_397), .B1(n_404), .B2(n_392), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_602), .B(n_441), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_652), .B(n_459), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_652), .A2(n_415), .B1(n_416), .B2(n_406), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_649), .A2(n_420), .B(n_421), .C(n_417), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_648), .A2(n_426), .B1(n_427), .B2(n_422), .Y(n_767) );
BUFx3_ASAP7_75t_L g768 ( .A(n_654), .Y(n_768) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_648), .A2(n_479), .B1(n_459), .B2(n_353), .Y(n_769) );
BUFx3_ASAP7_75t_L g770 ( .A(n_611), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_646), .B(n_479), .Y(n_771) );
OR2x6_ASAP7_75t_L g772 ( .A(n_649), .B(n_431), .Y(n_772) );
INVx2_ASAP7_75t_SL g773 ( .A(n_651), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_643), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_651), .A2(n_435), .B1(n_437), .B2(n_432), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_643), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_645), .A2(n_440), .B(n_439), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_611), .B(n_325), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_647), .A2(n_446), .B(n_442), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_644), .B(n_445), .Y(n_780) );
BUFx12f_ASAP7_75t_L g781 ( .A(n_644), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_644), .Y(n_782) );
INVxp67_ASAP7_75t_L g783 ( .A(n_644), .Y(n_783) );
OR2x6_ASAP7_75t_L g784 ( .A(n_650), .B(n_448), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_657), .A2(n_450), .B(n_449), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_650), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_650), .B(n_452), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_650), .B(n_372), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_577), .A2(n_460), .B1(n_461), .B2(n_456), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_580), .B(n_464), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_635), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_577), .A2(n_465), .B1(n_467), .B2(n_463), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_666), .Y(n_793) );
OAI21x1_ASAP7_75t_L g794 ( .A1(n_782), .A2(n_375), .B(n_367), .Y(n_794) );
OA21x2_ASAP7_75t_L g795 ( .A1(n_787), .A2(n_400), .B(n_388), .Y(n_795) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_716), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_662), .A2(n_405), .B(n_400), .Y(n_797) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_716), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_733), .Y(n_799) );
INVx6_ASAP7_75t_L g800 ( .A(n_746), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_743), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_750), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_680), .B(n_472), .Y(n_803) );
OAI21x1_ASAP7_75t_L g804 ( .A1(n_782), .A2(n_786), .B(n_787), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_690), .B(n_478), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_703), .Y(n_806) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_686), .A2(n_424), .B(n_405), .Y(n_807) );
OAI21x1_ASAP7_75t_L g808 ( .A1(n_790), .A2(n_443), .B(n_424), .Y(n_808) );
A2O1A1Ixp33_ASAP7_75t_L g809 ( .A1(n_718), .A2(n_443), .B(n_453), .C(n_464), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_695), .B(n_453), .Y(n_810) );
OAI21x1_ASAP7_75t_L g811 ( .A1(n_790), .A2(n_518), .B(n_516), .Y(n_811) );
NOR2xp33_ASAP7_75t_SL g812 ( .A(n_784), .B(n_379), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_697), .B(n_381), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_729), .A2(n_518), .B(n_521), .Y(n_814) );
OAI221xp5_ASAP7_75t_L g815 ( .A1(n_680), .A2(n_476), .B1(n_383), .B2(n_393), .C(n_394), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_747), .A2(n_476), .B(n_326), .C(n_396), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_738), .Y(n_817) );
BUFx3_ASAP7_75t_L g818 ( .A(n_704), .Y(n_818) );
AND2x4_ASAP7_75t_L g819 ( .A(n_693), .B(n_5), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_687), .B(n_539), .C(n_541), .Y(n_820) );
A2O1A1Ixp33_ASAP7_75t_L g821 ( .A1(n_699), .A2(n_539), .B(n_554), .C(n_541), .Y(n_821) );
BUFx8_ASAP7_75t_L g822 ( .A(n_668), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_680), .A2(n_554), .B1(n_562), .B2(n_541), .Y(n_823) );
AO21x1_ASAP7_75t_L g824 ( .A1(n_767), .A2(n_90), .B(n_89), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_752), .Y(n_825) );
AOI222xp33_ASAP7_75t_L g826 ( .A1(n_669), .A2(n_717), .B1(n_678), .B2(n_681), .C1(n_700), .C2(n_705), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_679), .Y(n_827) );
CKINVDCx6p67_ASAP7_75t_R g828 ( .A(n_725), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_700), .A2(n_554), .B1(n_562), .B2(n_541), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_664), .B(n_7), .Y(n_830) );
AO21x2_ASAP7_75t_L g831 ( .A1(n_698), .A2(n_554), .B(n_541), .Y(n_831) );
OR2x2_ASAP7_75t_L g832 ( .A(n_660), .B(n_10), .Y(n_832) );
OR3x4_ASAP7_75t_SL g833 ( .A(n_669), .B(n_10), .C(n_11), .Y(n_833) );
OA21x2_ASAP7_75t_L g834 ( .A1(n_760), .A2(n_562), .B(n_554), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_709), .Y(n_835) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_781), .Y(n_836) );
NAND2x1p5_ASAP7_75t_L g837 ( .A(n_738), .B(n_12), .Y(n_837) );
OAI21x1_ASAP7_75t_L g838 ( .A1(n_774), .A2(n_94), .B(n_91), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_677), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_752), .Y(n_840) );
INVx1_ASAP7_75t_SL g841 ( .A(n_660), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_755), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_684), .B(n_13), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_664), .B(n_13), .Y(n_844) );
OAI21x1_ASAP7_75t_L g845 ( .A1(n_755), .A2(n_98), .B(n_96), .Y(n_845) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_667), .Y(n_846) );
AO21x2_ASAP7_75t_L g847 ( .A1(n_698), .A2(n_562), .B(n_100), .Y(n_847) );
OA21x2_ASAP7_75t_L g848 ( .A1(n_779), .A2(n_562), .B(n_101), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_683), .B(n_663), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_709), .Y(n_850) );
OA21x2_ASAP7_75t_L g851 ( .A1(n_785), .A2(n_102), .B(n_99), .Y(n_851) );
OAI21x1_ASAP7_75t_L g852 ( .A1(n_777), .A2(n_106), .B(n_103), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_758), .Y(n_853) );
OAI21x1_ASAP7_75t_L g854 ( .A1(n_778), .A2(n_111), .B(n_107), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_665), .B(n_14), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_673), .Y(n_856) );
OA21x2_ASAP7_75t_L g857 ( .A1(n_783), .A2(n_116), .B(n_112), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g858 ( .A1(n_735), .A2(n_15), .B(n_16), .Y(n_858) );
OAI21xp5_ASAP7_75t_L g859 ( .A1(n_789), .A2(n_16), .B(n_17), .Y(n_859) );
NOR2x1_ASAP7_75t_R g860 ( .A(n_768), .B(n_17), .Y(n_860) );
BUFx5_ASAP7_75t_L g861 ( .A(n_770), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_676), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_705), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_766), .A2(n_18), .B(n_19), .C(n_20), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_791), .B(n_21), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_715), .Y(n_866) );
OAI21x1_ASAP7_75t_L g867 ( .A1(n_734), .A2(n_119), .B(n_117), .Y(n_867) );
OAI21x1_ASAP7_75t_L g868 ( .A1(n_749), .A2(n_125), .B(n_120), .Y(n_868) );
OAI21x1_ASAP7_75t_L g869 ( .A1(n_728), .A2(n_129), .B(n_128), .Y(n_869) );
OAI21x1_ASAP7_75t_L g870 ( .A1(n_728), .A2(n_133), .B(n_131), .Y(n_870) );
AND2x4_ASAP7_75t_L g871 ( .A(n_702), .B(n_21), .Y(n_871) );
OAI21x1_ASAP7_75t_L g872 ( .A1(n_723), .A2(n_138), .B(n_137), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_708), .A2(n_23), .B(n_25), .C(n_26), .Y(n_873) );
OAI21x1_ASAP7_75t_L g874 ( .A1(n_723), .A2(n_141), .B(n_140), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_744), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_720), .B(n_730), .Y(n_876) );
OAI21x1_ASAP7_75t_L g877 ( .A1(n_659), .A2(n_147), .B(n_142), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_730), .B(n_23), .Y(n_878) );
NOR2x1_ASAP7_75t_R g879 ( .A(n_667), .B(n_26), .Y(n_879) );
OAI21x1_ASAP7_75t_L g880 ( .A1(n_659), .A2(n_150), .B(n_148), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_784), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_881) );
NOR2xp67_ASAP7_75t_L g882 ( .A(n_756), .B(n_27), .Y(n_882) );
OAI21xp5_ASAP7_75t_L g883 ( .A1(n_789), .A2(n_28), .B(n_29), .Y(n_883) );
CKINVDCx11_ASAP7_75t_R g884 ( .A(n_737), .Y(n_884) );
OR2x2_ASAP7_75t_L g885 ( .A(n_689), .B(n_30), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_671), .Y(n_886) );
CKINVDCx11_ASAP7_75t_R g887 ( .A(n_667), .Y(n_887) );
OAI21x1_ASAP7_75t_L g888 ( .A1(n_661), .A2(n_154), .B(n_153), .Y(n_888) );
BUFx3_ASAP7_75t_L g889 ( .A(n_722), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_784), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_744), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_727), .Y(n_892) );
OAI21x1_ASAP7_75t_L g893 ( .A1(n_661), .A2(n_156), .B(n_155), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_692), .Y(n_894) );
INVx3_ASAP7_75t_L g895 ( .A(n_707), .Y(n_895) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_792), .A2(n_31), .B(n_32), .Y(n_896) );
BUFx6f_ASAP7_75t_L g897 ( .A(n_736), .Y(n_897) );
OAI22xp5_ASAP7_75t_SL g898 ( .A1(n_740), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_682), .Y(n_899) );
OAI21x1_ASAP7_75t_L g900 ( .A1(n_767), .A2(n_163), .B(n_162), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_792), .B(n_731), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g902 ( .A1(n_754), .A2(n_33), .B1(n_35), .B2(n_37), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_675), .A2(n_195), .B(n_314), .Y(n_903) );
AO21x2_ASAP7_75t_L g904 ( .A1(n_708), .A2(n_192), .B(n_312), .Y(n_904) );
OR2x6_ASAP7_75t_L g905 ( .A(n_772), .B(n_38), .Y(n_905) );
OAI21xp5_ASAP7_75t_L g906 ( .A1(n_674), .A2(n_40), .B(n_41), .Y(n_906) );
AO21x2_ASAP7_75t_L g907 ( .A1(n_775), .A2(n_196), .B(n_311), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_658), .B(n_40), .Y(n_908) );
OAI21x1_ASAP7_75t_L g909 ( .A1(n_691), .A2(n_198), .B(n_309), .Y(n_909) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_753), .B(n_43), .C(n_44), .Y(n_910) );
AOI21xp33_ASAP7_75t_L g911 ( .A1(n_772), .A2(n_45), .B(n_46), .Y(n_911) );
OAI21xp5_ASAP7_75t_L g912 ( .A1(n_739), .A2(n_46), .B(n_47), .Y(n_912) );
NOR2xp33_ASAP7_75t_SL g913 ( .A(n_736), .B(n_165), .Y(n_913) );
OAI21x1_ASAP7_75t_L g914 ( .A1(n_696), .A2(n_201), .B(n_307), .Y(n_914) );
NOR3xp33_ASAP7_75t_L g915 ( .A(n_751), .B(n_47), .C(n_48), .Y(n_915) );
BUFx4f_ASAP7_75t_L g916 ( .A(n_707), .Y(n_916) );
AOI22x1_ASAP7_75t_L g917 ( .A1(n_776), .A2(n_202), .B1(n_305), .B2(n_304), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_682), .Y(n_918) );
OAI21x1_ASAP7_75t_L g919 ( .A1(n_710), .A2(n_199), .B(n_303), .Y(n_919) );
INVx4_ASAP7_75t_L g920 ( .A(n_707), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_711), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_739), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_922) );
OAI22x1_ASAP7_75t_L g923 ( .A1(n_741), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_682), .Y(n_924) );
AND2x4_ASAP7_75t_L g925 ( .A(n_726), .B(n_52), .Y(n_925) );
INVx3_ASAP7_75t_L g926 ( .A(n_670), .Y(n_926) );
OAI21x1_ASAP7_75t_L g927 ( .A1(n_780), .A2(n_213), .B(n_302), .Y(n_927) );
AOI21xp33_ASAP7_75t_L g928 ( .A1(n_772), .A2(n_52), .B(n_53), .Y(n_928) );
OAI21x1_ASAP7_75t_L g929 ( .A1(n_670), .A2(n_214), .B(n_301), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_721), .B(n_53), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_742), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_742), .A2(n_191), .B(n_300), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_765), .Y(n_933) );
OAI21x1_ASAP7_75t_SL g934 ( .A1(n_721), .A2(n_54), .B(n_55), .Y(n_934) );
O2A1O1Ixp33_ASAP7_75t_SL g935 ( .A1(n_724), .A2(n_215), .B(n_296), .C(n_290), .Y(n_935) );
OAI21xp5_ASAP7_75t_L g936 ( .A1(n_765), .A2(n_54), .B(n_56), .Y(n_936) );
AO31x2_ASAP7_75t_L g937 ( .A1(n_775), .A2(n_57), .A3(n_58), .B(n_59), .Y(n_937) );
AOI21xp5_ASAP7_75t_L g938 ( .A1(n_724), .A2(n_763), .B(n_719), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_719), .B(n_741), .Y(n_939) );
BUFx3_ASAP7_75t_L g940 ( .A(n_711), .Y(n_940) );
AO21x2_ASAP7_75t_L g941 ( .A1(n_757), .A2(n_188), .B(n_289), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_826), .A2(n_706), .B1(n_714), .B2(n_732), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_835), .B(n_732), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_793), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_826), .A2(n_713), .B1(n_711), .B2(n_712), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_817), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_849), .A2(n_712), .B1(n_713), .B2(n_745), .Y(n_947) );
OAI21x1_ASAP7_75t_L g948 ( .A1(n_804), .A2(n_672), .B(n_685), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_796), .B(n_672), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_933), .A2(n_713), .B1(n_712), .B2(n_759), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_817), .Y(n_951) );
AOI222xp33_ASAP7_75t_L g952 ( .A1(n_860), .A2(n_762), .B1(n_764), .B2(n_726), .C1(n_771), .C2(n_773), .Y(n_952) );
AOI211xp5_ASAP7_75t_L g953 ( .A1(n_898), .A2(n_788), .B(n_748), .C(n_688), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_866), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_905), .A2(n_901), .B1(n_859), .B2(n_896), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_799), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_801), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g958 ( .A(n_806), .Y(n_958) );
AOI21xp5_ASAP7_75t_L g959 ( .A1(n_938), .A2(n_761), .B(n_736), .Y(n_959) );
OA21x2_ASAP7_75t_L g960 ( .A1(n_797), .A2(n_761), .B(n_688), .Y(n_960) );
INVx3_ASAP7_75t_L g961 ( .A(n_836), .Y(n_961) );
AOI22xp33_ASAP7_75t_SL g962 ( .A1(n_905), .A2(n_726), .B1(n_701), .B2(n_694), .Y(n_962) );
AOI222xp33_ASAP7_75t_L g963 ( .A1(n_894), .A2(n_688), .B1(n_694), .B2(n_701), .C1(n_60), .C2(n_61), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_796), .B(n_694), .Y(n_964) );
OAI21xp5_ASAP7_75t_L g965 ( .A1(n_901), .A2(n_931), .B(n_809), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_850), .B(n_769), .Y(n_966) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_798), .Y(n_967) );
OR2x6_ASAP7_75t_L g968 ( .A(n_905), .B(n_701), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_819), .A2(n_761), .B1(n_58), .B2(n_59), .Y(n_969) );
A2O1A1Ixp33_ASAP7_75t_L g970 ( .A1(n_859), .A2(n_57), .B(n_60), .C(n_62), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_802), .Y(n_971) );
CKINVDCx11_ASAP7_75t_R g972 ( .A(n_818), .Y(n_972) );
AO31x2_ASAP7_75t_L g973 ( .A1(n_824), .A2(n_63), .A3(n_64), .B(n_65), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_883), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_798), .B(n_66), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_876), .B(n_66), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_855), .Y(n_977) );
OAI211xp5_ASAP7_75t_L g978 ( .A1(n_902), .A2(n_863), .B(n_896), .C(n_883), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_812), .A2(n_225), .B(n_285), .Y(n_979) );
AO21x2_ASAP7_75t_L g980 ( .A1(n_831), .A2(n_222), .B(n_284), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g981 ( .A1(n_814), .A2(n_220), .B(n_283), .Y(n_981) );
CKINVDCx14_ASAP7_75t_R g982 ( .A(n_800), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_855), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_865), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_841), .B(n_67), .Y(n_985) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_803), .A2(n_68), .B1(n_69), .B2(n_70), .C(n_71), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_865), .Y(n_987) );
AND2x4_ASAP7_75t_L g988 ( .A(n_836), .B(n_69), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_819), .A2(n_70), .B1(n_72), .B2(n_73), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_871), .Y(n_990) );
A2O1A1Ixp33_ASAP7_75t_L g991 ( .A1(n_936), .A2(n_72), .B(n_74), .C(n_75), .Y(n_991) );
INVx4_ASAP7_75t_L g992 ( .A(n_836), .Y(n_992) );
OA21x2_ASAP7_75t_L g993 ( .A1(n_794), .A2(n_232), .B(n_278), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_841), .A2(n_75), .B1(n_76), .B2(n_77), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_856), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g996 ( .A1(n_837), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_996) );
OA21x2_ASAP7_75t_L g997 ( .A1(n_854), .A2(n_237), .B(n_276), .Y(n_997) );
INVxp67_ASAP7_75t_SL g998 ( .A(n_908), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_936), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_871), .Y(n_1000) );
OAI21xp5_ASAP7_75t_L g1001 ( .A1(n_930), .A2(n_80), .B(n_82), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_822), .Y(n_1002) );
AOI21xp5_ASAP7_75t_L g1003 ( .A1(n_814), .A2(n_821), .B(n_810), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_939), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_862), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_837), .A2(n_85), .B1(n_166), .B2(n_167), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_853), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_830), .Y(n_1008) );
AOI221xp5_ASAP7_75t_SL g1009 ( .A1(n_912), .A2(n_169), .B1(n_170), .B2(n_172), .C(n_173), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_830), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_805), .B(n_177), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_843), .B(n_178), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_844), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_881), .A2(n_179), .B1(n_183), .B2(n_184), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_889), .Y(n_1015) );
OAI21xp5_ASAP7_75t_L g1016 ( .A1(n_930), .A2(n_185), .B(n_217), .Y(n_1016) );
AOI211xp5_ASAP7_75t_L g1017 ( .A1(n_878), .A2(n_228), .B(n_230), .C(n_231), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_875), .B(n_235), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_891), .B(n_240), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_800), .A2(n_815), .B1(n_886), .B2(n_832), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_844), .Y(n_1021) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_915), .B(n_241), .C(n_242), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_908), .Y(n_1023) );
INVx2_ASAP7_75t_L g1024 ( .A(n_846), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_828), .B(n_250), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g1026 ( .A1(n_827), .A2(n_252), .B1(n_253), .B2(n_256), .C(n_257), .Y(n_1026) );
AO21x2_ASAP7_75t_L g1027 ( .A1(n_831), .A2(n_261), .B(n_264), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_805), .B(n_265), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_885), .A2(n_266), .B1(n_268), .B2(n_269), .Y(n_1029) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_800), .A2(n_271), .B1(n_315), .B2(n_815), .Y(n_1030) );
INVx2_ASAP7_75t_L g1031 ( .A(n_846), .Y(n_1031) );
AOI21xp5_ASAP7_75t_L g1032 ( .A1(n_932), .A2(n_834), .B(n_935), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_925), .A2(n_882), .B1(n_881), .B2(n_890), .Y(n_1033) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_892), .A2(n_912), .B1(n_858), .B2(n_890), .C(n_906), .Y(n_1034) );
OAI22xp33_ASAP7_75t_L g1035 ( .A1(n_813), .A2(n_923), .B1(n_858), .B2(n_911), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_825), .B(n_840), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_863), .A2(n_922), .B1(n_829), .B2(n_823), .Y(n_1037) );
OAI22x1_ASAP7_75t_L g1038 ( .A1(n_833), .A2(n_879), .B1(n_857), .B2(n_917), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_906), .A2(n_928), .B1(n_911), .B2(n_922), .C(n_807), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_910), .A2(n_887), .B1(n_928), .B2(n_884), .Y(n_1040) );
OAI222xp33_ASAP7_75t_L g1041 ( .A1(n_829), .A2(n_932), .B1(n_839), .B2(n_823), .C1(n_842), .C2(n_926), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_822), .A2(n_934), .B1(n_920), .B2(n_926), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_916), .A2(n_920), .B1(n_913), .B2(n_846), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_940), .A2(n_895), .B1(n_916), .B2(n_807), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_895), .A2(n_921), .B1(n_820), .B2(n_907), .Y(n_1045) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_897), .Y(n_1046) );
NAND2x1_ASAP7_75t_L g1047 ( .A(n_897), .B(n_899), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_816), .B(n_795), .Y(n_1048) );
AOI21xp5_ASAP7_75t_L g1049 ( .A1(n_834), .A2(n_847), .B(n_795), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1050 ( .A1(n_864), .A2(n_873), .B1(n_913), .B2(n_857), .C(n_851), .Y(n_1050) );
CKINVDCx6p67_ASAP7_75t_R g1051 ( .A(n_861), .Y(n_1051) );
INVx2_ASAP7_75t_L g1052 ( .A(n_808), .Y(n_1052) );
OAI21xp5_ASAP7_75t_L g1053 ( .A1(n_900), .A2(n_927), .B(n_811), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_907), .A2(n_861), .B1(n_941), .B2(n_924), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_861), .A2(n_941), .B1(n_918), .B2(n_904), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_937), .Y(n_1056) );
AOI21xp5_ASAP7_75t_L g1057 ( .A1(n_847), .A2(n_848), .B(n_851), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_861), .A2(n_904), .B1(n_848), .B2(n_897), .Y(n_1058) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_937), .A2(n_852), .B1(n_929), .B2(n_845), .C(n_868), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1060 ( .A1(n_937), .A2(n_867), .B1(n_914), .B2(n_919), .C(n_909), .Y(n_1060) );
AND2x4_ASAP7_75t_L g1061 ( .A(n_877), .B(n_893), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_880), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_888), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_861), .B(n_872), .Y(n_1064) );
OAI211xp5_ASAP7_75t_L g1065 ( .A1(n_874), .A2(n_869), .B(n_870), .C(n_903), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_861), .A2(n_680), .B1(n_826), .B2(n_574), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_838), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_793), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_793), .Y(n_1069) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_939), .A2(n_574), .B1(n_717), .B2(n_849), .C(n_826), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_894), .B(n_849), .Y(n_1071) );
INVx3_ASAP7_75t_L g1072 ( .A(n_1051), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1056), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_956), .B(n_957), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_971), .B(n_995), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_955), .B(n_1071), .Y(n_1076) );
INVx2_ASAP7_75t_SL g1077 ( .A(n_992), .Y(n_1077) );
AOI222xp33_ASAP7_75t_L g1078 ( .A1(n_1070), .A2(n_955), .B1(n_942), .B2(n_1066), .C1(n_1034), .C2(n_974), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1007), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_944), .B(n_954), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1005), .B(n_1068), .Y(n_1081) );
OAI21x1_ASAP7_75t_L g1082 ( .A1(n_1049), .A2(n_1057), .B(n_1032), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_967), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1084 ( .A(n_1023), .Y(n_1084) );
NAND2x1_ASAP7_75t_L g1085 ( .A(n_1061), .B(n_1064), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_998), .B(n_946), .Y(n_1086) );
INVx3_ASAP7_75t_L g1087 ( .A(n_964), .Y(n_1087) );
OR2x2_ASAP7_75t_L g1088 ( .A(n_951), .B(n_1021), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_960), .Y(n_1089) );
INVx4_ASAP7_75t_L g1090 ( .A(n_968), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1069), .Y(n_1091) );
AOI22xp33_ASAP7_75t_SL g1092 ( .A1(n_978), .A2(n_974), .B1(n_999), .B2(n_1006), .Y(n_1092) );
AND2x4_ASAP7_75t_L g1093 ( .A(n_968), .B(n_964), .Y(n_1093) );
BUFx2_ASAP7_75t_L g1094 ( .A(n_968), .Y(n_1094) );
INVx2_ASAP7_75t_L g1095 ( .A(n_960), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_977), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1063), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_985), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_975), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_1046), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1062), .Y(n_1101) );
INVx2_ASAP7_75t_L g1102 ( .A(n_1067), .Y(n_1102) );
INVxp67_ASAP7_75t_L g1103 ( .A(n_1002), .Y(n_1103) );
NOR2x1p5_ASAP7_75t_L g1104 ( .A(n_958), .B(n_992), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_983), .B(n_984), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_987), .B(n_965), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_965), .B(n_1001), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_945), .B(n_1033), .Y(n_1108) );
OAI21xp5_ASAP7_75t_L g1109 ( .A1(n_1037), .A2(n_1039), .B(n_1035), .Y(n_1109) );
NAND2xp5_ASAP7_75t_SL g1110 ( .A(n_1038), .B(n_1020), .Y(n_1110) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_1015), .Y(n_1111) );
INVxp67_ASAP7_75t_L g1112 ( .A(n_961), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1001), .B(n_963), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_943), .B(n_1008), .Y(n_1114) );
OA21x2_ASAP7_75t_L g1115 ( .A1(n_1054), .A2(n_1055), .B(n_1058), .Y(n_1115) );
INVx1_ASAP7_75t_SL g1116 ( .A(n_972), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_990), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_963), .B(n_999), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1000), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_943), .B(n_949), .Y(n_1120) );
INVx2_ASAP7_75t_SL g1121 ( .A(n_949), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_966), .B(n_1018), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1036), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1036), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_976), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_966), .B(n_1018), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_988), .B(n_1010), .Y(n_1127) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_1013), .B(n_1024), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_988), .Y(n_1129) );
AOI22xp33_ASAP7_75t_SL g1130 ( .A1(n_1006), .A2(n_1014), .B1(n_1037), .B2(n_982), .Y(n_1130) );
OR2x6_ASAP7_75t_L g1131 ( .A(n_1014), .B(n_1061), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_1031), .Y(n_1132) );
AND2x4_ASAP7_75t_SL g1133 ( .A(n_1025), .B(n_950), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_970), .B(n_991), .Y(n_1134) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_1047), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1012), .B(n_973), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_973), .B(n_996), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_1042), .B(n_1040), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_994), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_973), .B(n_962), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_989), .Y(n_1141) );
INVx2_ASAP7_75t_L g1142 ( .A(n_993), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_953), .B(n_1028), .Y(n_1143) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_1016), .B(n_948), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_986), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1011), .B(n_1004), .Y(n_1146) );
INVx3_ASAP7_75t_L g1147 ( .A(n_1052), .Y(n_1147) );
INVx2_ASAP7_75t_L g1148 ( .A(n_997), .Y(n_1148) );
NOR2x1_ASAP7_75t_L g1149 ( .A(n_1030), .B(n_1022), .Y(n_1149) );
INVx5_ASAP7_75t_L g1150 ( .A(n_1043), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_980), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_980), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_952), .B(n_947), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_969), .B(n_1044), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1048), .B(n_1045), .Y(n_1155) );
NOR2xp33_ASAP7_75t_L g1156 ( .A(n_1041), .B(n_1019), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1027), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1027), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1048), .Y(n_1159) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_1017), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1029), .B(n_1009), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1003), .B(n_1059), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1060), .B(n_1053), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1050), .Y(n_1164) );
INVx2_ASAP7_75t_SL g1165 ( .A(n_979), .Y(n_1165) );
AND2x4_ASAP7_75t_L g1166 ( .A(n_1053), .B(n_959), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1065), .Y(n_1167) );
INVx2_ASAP7_75t_SL g1168 ( .A(n_1026), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_981), .Y(n_1169) );
INVx2_ASAP7_75t_SL g1170 ( .A(n_1072), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1106), .B(n_1120), .Y(n_1171) );
INVx3_ASAP7_75t_L g1172 ( .A(n_1085), .Y(n_1172) );
INVx3_ASAP7_75t_L g1173 ( .A(n_1085), .Y(n_1173) );
INVx3_ASAP7_75t_L g1174 ( .A(n_1131), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1073), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1073), .Y(n_1176) );
NOR2x1_ASAP7_75t_L g1177 ( .A(n_1110), .B(n_1090), .Y(n_1177) );
INVx1_ASAP7_75t_SL g1178 ( .A(n_1100), .Y(n_1178) );
BUFx2_ASAP7_75t_L g1179 ( .A(n_1131), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1076), .B(n_1108), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1097), .Y(n_1181) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_1083), .Y(n_1182) );
INVx2_ASAP7_75t_L g1183 ( .A(n_1097), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1102), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1106), .B(n_1120), .Y(n_1185) );
NOR2x1_ASAP7_75t_L g1186 ( .A(n_1104), .B(n_1072), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1102), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1107), .B(n_1080), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1131), .B(n_1140), .Y(n_1189) );
HB1xp67_ASAP7_75t_L g1190 ( .A(n_1111), .Y(n_1190) );
INVx4_ASAP7_75t_L g1191 ( .A(n_1072), .Y(n_1191) );
AOI221xp5_ASAP7_75t_L g1192 ( .A1(n_1109), .A2(n_1099), .B1(n_1145), .B2(n_1113), .C(n_1125), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1096), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1107), .B(n_1080), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1096), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1136), .B(n_1075), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1136), .B(n_1075), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1079), .Y(n_1198) );
INVx4_ASAP7_75t_L g1199 ( .A(n_1090), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1074), .B(n_1163), .Y(n_1200) );
OAI211xp5_ASAP7_75t_SL g1201 ( .A1(n_1103), .A2(n_1138), .B(n_1081), .C(n_1098), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1105), .B(n_1074), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1163), .B(n_1122), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1114), .B(n_1091), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1159), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1076), .B(n_1108), .Y(n_1206) );
NOR2xp67_ASAP7_75t_L g1207 ( .A(n_1077), .B(n_1138), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1122), .B(n_1126), .Y(n_1208) );
AO21x2_ASAP7_75t_L g1209 ( .A1(n_1157), .A2(n_1158), .B(n_1148), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1101), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1101), .Y(n_1211) );
AOI22xp5_ASAP7_75t_L g1212 ( .A1(n_1113), .A2(n_1118), .B1(n_1130), .B2(n_1078), .Y(n_1212) );
AOI21xp5_ASAP7_75t_SL g1213 ( .A1(n_1131), .A2(n_1118), .B(n_1090), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_1092), .A2(n_1153), .B1(n_1126), .B2(n_1168), .Y(n_1214) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1089), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1086), .B(n_1088), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1217 ( .A1(n_1168), .A2(n_1133), .B1(n_1160), .B2(n_1141), .Y(n_1217) );
AND2x2_ASAP7_75t_SL g1218 ( .A(n_1094), .B(n_1133), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1162), .B(n_1140), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1162), .B(n_1137), .Y(n_1220) );
HB1xp67_ASAP7_75t_L g1221 ( .A(n_1086), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1147), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1095), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1147), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1123), .Y(n_1225) );
BUFx3_ASAP7_75t_L g1226 ( .A(n_1077), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1137), .B(n_1164), .Y(n_1227) );
AOI22xp5_ASAP7_75t_L g1228 ( .A1(n_1143), .A2(n_1146), .B1(n_1127), .B2(n_1156), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_1139), .A2(n_1143), .B1(n_1146), .B2(n_1134), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1114), .B(n_1124), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1155), .B(n_1084), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1164), .B(n_1119), .Y(n_1232) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_1117), .A2(n_1134), .B1(n_1129), .B2(n_1127), .C(n_1154), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1167), .Y(n_1234) );
NOR2xp33_ASAP7_75t_R g1235 ( .A(n_1116), .B(n_1121), .Y(n_1235) );
BUFx3_ASAP7_75t_L g1236 ( .A(n_1121), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1167), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1155), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1198), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_1216), .B(n_1132), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1188), .B(n_1128), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1219), .B(n_1166), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1188), .B(n_1128), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1244 ( .A(n_1212), .B(n_1112), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1219), .B(n_1166), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1220), .B(n_1166), .Y(n_1246) );
INVxp67_ASAP7_75t_SL g1247 ( .A(n_1207), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1194), .B(n_1200), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1221), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1200), .B(n_1087), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1201), .B(n_1087), .Y(n_1251) );
OAI21xp5_ASAP7_75t_L g1252 ( .A1(n_1214), .A2(n_1161), .B(n_1149), .Y(n_1252) );
NOR2xp33_ASAP7_75t_R g1253 ( .A(n_1218), .B(n_1150), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1215), .Y(n_1254) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1215), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1196), .B(n_1197), .Y(n_1256) );
NAND5xp2_ASAP7_75t_L g1257 ( .A(n_1192), .B(n_1169), .C(n_1150), .D(n_1093), .E(n_1165), .Y(n_1257) );
BUFx2_ASAP7_75t_L g1258 ( .A(n_1226), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1196), .B(n_1115), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1197), .B(n_1115), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1193), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1231), .B(n_1152), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1171), .B(n_1144), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1185), .B(n_1144), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1195), .Y(n_1265) );
INVx1_ASAP7_75t_SL g1266 ( .A(n_1235), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1185), .B(n_1135), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1195), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1227), .B(n_1144), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1202), .B(n_1151), .Y(n_1270) );
NOR2x1_ASAP7_75t_L g1271 ( .A(n_1186), .B(n_1152), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1272 ( .A(n_1228), .B(n_1180), .Y(n_1272) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_1190), .Y(n_1273) );
NAND2x1p5_ASAP7_75t_L g1274 ( .A(n_1191), .B(n_1150), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1203), .B(n_1082), .Y(n_1275) );
INVx1_ASAP7_75t_SL g1276 ( .A(n_1178), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1203), .B(n_1208), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1204), .B(n_1142), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1230), .B(n_1225), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1182), .B(n_1231), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1175), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1180), .B(n_1206), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1206), .B(n_1205), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1189), .B(n_1238), .Y(n_1284) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_1189), .B(n_1174), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1175), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1287 ( .A(n_1191), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1239), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1256), .B(n_1229), .Y(n_1289) );
AOI22x1_ASAP7_75t_L g1290 ( .A1(n_1266), .A2(n_1191), .B1(n_1199), .B2(n_1170), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1282), .B(n_1179), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1261), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1256), .B(n_1179), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1277), .B(n_1225), .Y(n_1294) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1254), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1259), .B(n_1174), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1280), .B(n_1234), .Y(n_1297) );
HB1xp67_ASAP7_75t_L g1298 ( .A(n_1273), .Y(n_1298) );
INVx2_ASAP7_75t_SL g1299 ( .A(n_1258), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1260), .B(n_1176), .Y(n_1300) );
INVx2_ASAP7_75t_L g1301 ( .A(n_1254), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1275), .B(n_1234), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1277), .B(n_1232), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1265), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1275), .B(n_1237), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1249), .B(n_1237), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1242), .B(n_1183), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1242), .B(n_1183), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1268), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1281), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1245), .B(n_1187), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1245), .B(n_1187), .Y(n_1312) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_1247), .A2(n_1213), .B1(n_1218), .B2(n_1217), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1272), .B(n_1233), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1286), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1283), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1255), .Y(n_1317) );
NOR2x1p5_ASAP7_75t_L g1318 ( .A(n_1267), .B(n_1172), .Y(n_1318) );
OR2x6_ASAP7_75t_L g1319 ( .A(n_1287), .B(n_1213), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1246), .B(n_1223), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1246), .B(n_1223), .Y(n_1321) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1255), .Y(n_1322) );
AOI221x1_ASAP7_75t_L g1323 ( .A1(n_1252), .A2(n_1222), .B1(n_1224), .B2(n_1172), .C(n_1173), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1270), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1248), .B(n_1184), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1303), .B(n_1240), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1327 ( .A(n_1314), .B(n_1276), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1298), .Y(n_1328) );
AOI21xp5_ASAP7_75t_L g1329 ( .A1(n_1319), .A2(n_1313), .B(n_1290), .Y(n_1329) );
NAND2xp5_ASAP7_75t_SL g1330 ( .A(n_1290), .B(n_1287), .Y(n_1330) );
AOI21xp5_ASAP7_75t_L g1331 ( .A1(n_1319), .A2(n_1257), .B(n_1177), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1324), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1300), .B(n_1284), .Y(n_1333) );
NOR2xp67_ASAP7_75t_SL g1334 ( .A(n_1299), .B(n_1199), .Y(n_1334) );
OAI21xp33_ASAP7_75t_L g1335 ( .A1(n_1293), .A2(n_1244), .B(n_1251), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1306), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1297), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1325), .Y(n_1338) );
NOR2xp33_ASAP7_75t_L g1339 ( .A(n_1289), .B(n_1279), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1302), .B(n_1250), .Y(n_1340) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1295), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1325), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1288), .Y(n_1343) );
AOI21xp5_ASAP7_75t_L g1344 ( .A1(n_1319), .A2(n_1274), .B(n_1172), .Y(n_1344) );
OAI21xp5_ASAP7_75t_L g1345 ( .A1(n_1330), .A2(n_1323), .B(n_1299), .Y(n_1345) );
NAND2xp33_ASAP7_75t_SL g1346 ( .A(n_1334), .B(n_1253), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1343), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_1330), .A2(n_1319), .B1(n_1318), .B2(n_1291), .Y(n_1348) );
A2O1A1Ixp33_ASAP7_75t_L g1349 ( .A1(n_1329), .A2(n_1291), .B(n_1294), .C(n_1173), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1338), .B(n_1296), .Y(n_1350) );
INVx2_ASAP7_75t_SL g1351 ( .A(n_1328), .Y(n_1351) );
AO22x2_ASAP7_75t_L g1352 ( .A1(n_1332), .A2(n_1316), .B1(n_1323), .B2(n_1310), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1342), .Y(n_1353) );
AOI21xp5_ASAP7_75t_L g1354 ( .A1(n_1331), .A2(n_1274), .B(n_1271), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1336), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1339), .B(n_1305), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1339), .B(n_1305), .Y(n_1357) );
INVx2_ASAP7_75t_SL g1358 ( .A(n_1326), .Y(n_1358) );
NAND2xp33_ASAP7_75t_SL g1359 ( .A(n_1337), .B(n_1253), .Y(n_1359) );
AOI322xp5_ASAP7_75t_L g1360 ( .A1(n_1327), .A2(n_1307), .A3(n_1311), .B1(n_1312), .B2(n_1308), .C1(n_1320), .C2(n_1321), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1360), .B(n_1335), .Y(n_1361) );
OAI21xp5_ASAP7_75t_L g1362 ( .A1(n_1349), .A2(n_1327), .B(n_1344), .Y(n_1362) );
OAI21xp33_ASAP7_75t_SL g1363 ( .A1(n_1345), .A2(n_1333), .B(n_1340), .Y(n_1363) );
AOI32xp33_ASAP7_75t_L g1364 ( .A1(n_1346), .A2(n_1321), .A3(n_1320), .B1(n_1311), .B2(n_1312), .Y(n_1364) );
AOI22xp5_ASAP7_75t_L g1365 ( .A1(n_1348), .A2(n_1285), .B1(n_1263), .B2(n_1264), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1347), .Y(n_1366) );
INVx2_ASAP7_75t_SL g1367 ( .A(n_1358), .Y(n_1367) );
AOI221x1_ASAP7_75t_L g1368 ( .A1(n_1352), .A2(n_1315), .B1(n_1288), .B2(n_1292), .C(n_1309), .Y(n_1368) );
NOR2xp33_ASAP7_75t_L g1369 ( .A(n_1356), .B(n_1285), .Y(n_1369) );
XOR2x2_ASAP7_75t_L g1370 ( .A(n_1357), .B(n_1241), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1366), .Y(n_1371) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_1363), .A2(n_1359), .B1(n_1354), .B2(n_1351), .C(n_1353), .Y(n_1372) );
AND2x4_ASAP7_75t_L g1373 ( .A(n_1367), .B(n_1355), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1361), .B(n_1350), .Y(n_1374) );
AOI211x1_ASAP7_75t_SL g1375 ( .A1(n_1362), .A2(n_1352), .B(n_1341), .C(n_1243), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1373), .B(n_1365), .Y(n_1376) );
NAND3xp33_ASAP7_75t_SL g1377 ( .A(n_1375), .B(n_1364), .C(n_1369), .Y(n_1377) );
HB1xp67_ASAP7_75t_L g1378 ( .A(n_1371), .Y(n_1378) );
NAND2x1p5_ASAP7_75t_L g1379 ( .A(n_1373), .B(n_1236), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1374), .Y(n_1380) );
AOI21xp5_ASAP7_75t_L g1381 ( .A1(n_1372), .A2(n_1368), .B(n_1370), .Y(n_1381) );
XNOR2xp5_ASAP7_75t_L g1382 ( .A(n_1380), .B(n_1236), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1383 ( .A(n_1377), .B(n_1262), .Y(n_1383) );
NOR3xp33_ASAP7_75t_L g1384 ( .A(n_1381), .B(n_1378), .C(n_1376), .Y(n_1384) );
NOR3x1_ASAP7_75t_L g1385 ( .A(n_1381), .B(n_1304), .C(n_1262), .Y(n_1385) );
INVx2_ASAP7_75t_SL g1386 ( .A(n_1382), .Y(n_1386) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1383), .Y(n_1387) );
OAI221xp5_ASAP7_75t_SL g1388 ( .A1(n_1384), .A2(n_1379), .B1(n_1269), .B2(n_1278), .C(n_1317), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1385), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1386), .B(n_1269), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1387), .Y(n_1391) );
OAI22xp5_ASAP7_75t_SL g1392 ( .A1(n_1391), .A2(n_1389), .B1(n_1388), .B2(n_1322), .Y(n_1392) );
AOI222xp33_ASAP7_75t_L g1393 ( .A1(n_1392), .A2(n_1390), .B1(n_1184), .B2(n_1181), .C1(n_1301), .C2(n_1211), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1393), .Y(n_1394) );
AOI21xp5_ASAP7_75t_L g1395 ( .A1(n_1394), .A2(n_1209), .B(n_1210), .Y(n_1395) );
endmodule