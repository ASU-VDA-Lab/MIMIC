module real_aes_8572_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g164 ( .A1(n_0), .A2(n_165), .B(n_166), .C(n_170), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_1), .B(n_159), .Y(n_172) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_2), .B(n_431), .C(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_3), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_4), .A2(n_153), .B(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_5), .A2(n_133), .B(n_150), .C(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_6), .A2(n_153), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_7), .B(n_159), .Y(n_456) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_8), .A2(n_125), .B(n_247), .Y(n_246) );
AND2x6_ASAP7_75t_L g150 ( .A(n_9), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_10), .A2(n_133), .B(n_150), .C(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g547 ( .A(n_11), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_12), .B(n_39), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_13), .B(n_169), .Y(n_496) );
INVx1_ASAP7_75t_L g130 ( .A(n_14), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_15), .B(n_144), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_16), .A2(n_145), .B(n_505), .C(n_507), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_17), .B(n_159), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_18), .B(n_187), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_19), .A2(n_133), .B(n_179), .C(n_186), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_20), .A2(n_168), .B(n_221), .C(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_21), .B(n_169), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_22), .B(n_169), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g474 ( .A(n_23), .Y(n_474) );
INVx1_ASAP7_75t_L g444 ( .A(n_24), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_25), .A2(n_133), .B(n_186), .C(n_250), .Y(n_249) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_26), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_27), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_28), .A2(n_100), .B1(n_709), .B2(n_716), .Y(n_99) );
INVx1_ASAP7_75t_L g468 ( .A(n_29), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_30), .A2(n_153), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g135 ( .A(n_31), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_32), .A2(n_148), .B(n_202), .C(n_203), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_33), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_34), .A2(n_168), .B(n_453), .C(n_455), .Y(n_452) );
INVxp67_ASAP7_75t_L g469 ( .A(n_35), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_36), .B(n_252), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_37), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_38), .A2(n_133), .B(n_186), .C(n_443), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_40), .A2(n_170), .B(n_545), .C(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_41), .B(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_42), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_43), .B(n_144), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_44), .B(n_153), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_45), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_46), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_47), .A2(n_148), .B(n_202), .C(n_230), .Y(n_229) );
AOI222xp33_ASAP7_75t_L g113 ( .A1(n_48), .A2(n_67), .B1(n_114), .B2(n_694), .C1(n_698), .C2(n_699), .Y(n_113) );
INVx1_ASAP7_75t_L g167 ( .A(n_49), .Y(n_167) );
INVx1_ASAP7_75t_L g231 ( .A(n_50), .Y(n_231) );
INVx1_ASAP7_75t_L g512 ( .A(n_51), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_52), .B(n_153), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_53), .Y(n_191) );
CKINVDCx14_ASAP7_75t_R g543 ( .A(n_54), .Y(n_543) );
INVx1_ASAP7_75t_L g151 ( .A(n_55), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_56), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_57), .B(n_159), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_58), .A2(n_140), .B(n_185), .C(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g129 ( .A(n_59), .Y(n_129) );
INVx1_ASAP7_75t_SL g454 ( .A(n_60), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_61), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_62), .B(n_144), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_63), .B(n_159), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_64), .B(n_145), .Y(n_218) );
INVx1_ASAP7_75t_L g477 ( .A(n_65), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_66), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_67), .Y(n_698) );
OAI22xp5_ASAP7_75t_SL g703 ( .A1(n_68), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_68), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_69), .B(n_181), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g132 ( .A1(n_70), .A2(n_133), .B(n_138), .C(n_148), .Y(n_132) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_71), .Y(n_240) );
INVx1_ASAP7_75t_L g714 ( .A(n_72), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_73), .A2(n_153), .B(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_74), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_75), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_76), .A2(n_153), .B(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_77), .A2(n_177), .B(n_464), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_78), .Y(n_441) );
INVx1_ASAP7_75t_L g503 ( .A(n_79), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_80), .B(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_81), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_82), .A2(n_153), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g506 ( .A(n_83), .Y(n_506) );
INVx2_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVx1_ASAP7_75t_L g495 ( .A(n_85), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_86), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_87), .B(n_169), .Y(n_219) );
OR2x2_ASAP7_75t_L g108 ( .A(n_88), .B(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g117 ( .A(n_88), .B(n_110), .Y(n_117) );
INVx2_ASAP7_75t_L g431 ( .A(n_88), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_89), .A2(n_133), .B(n_148), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_90), .B(n_153), .Y(n_200) );
INVx1_ASAP7_75t_L g204 ( .A(n_91), .Y(n_204) );
INVxp67_ASAP7_75t_L g243 ( .A(n_92), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_93), .B(n_125), .Y(n_548) );
INVx1_ASAP7_75t_L g139 ( .A(n_94), .Y(n_139) );
INVx1_ASAP7_75t_L g214 ( .A(n_95), .Y(n_214) );
INVx2_ASAP7_75t_L g515 ( .A(n_96), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_97), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g233 ( .A(n_98), .B(n_189), .Y(n_233) );
AOI22x1_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_113), .B1(n_700), .B2(n_702), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g701 ( .A(n_103), .Y(n_701) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_105), .A2(n_703), .B(n_707), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g708 ( .A(n_107), .Y(n_708) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2x2_ASAP7_75t_L g699 ( .A(n_109), .B(n_431), .Y(n_699) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g430 ( .A(n_110), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVxp67_ASAP7_75t_L g715 ( .A(n_112), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B1(n_428), .B2(n_432), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g696 ( .A(n_116), .Y(n_696) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g695 ( .A(n_118), .Y(n_695) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_118), .Y(n_704) );
OR3x1_ASAP7_75t_L g118 ( .A(n_119), .B(n_336), .C(n_385), .Y(n_118) );
NAND5xp2_ASAP7_75t_L g119 ( .A(n_120), .B(n_270), .C(n_299), .D(n_307), .E(n_322), .Y(n_119) );
O2A1O1Ixp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_193), .B(n_209), .C(n_254), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_173), .Y(n_121) );
AND2x2_ASAP7_75t_L g265 ( .A(n_122), .B(n_262), .Y(n_265) );
AND2x2_ASAP7_75t_L g298 ( .A(n_122), .B(n_174), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_122), .B(n_197), .Y(n_391) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_158), .Y(n_122) );
INVx2_ASAP7_75t_L g196 ( .A(n_123), .Y(n_196) );
BUFx2_ASAP7_75t_L g365 ( .A(n_123), .Y(n_365) );
AO21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_131), .B(n_156), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_124), .B(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_124), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_124), .B(n_208), .Y(n_207) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_124), .A2(n_213), .B(n_223), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_124), .B(n_447), .Y(n_446) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_124), .A2(n_473), .B(n_480), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_124), .B(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_125), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_125), .A2(n_248), .B(n_249), .Y(n_247) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g225 ( .A(n_126), .Y(n_225) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_127), .B(n_128), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_152), .Y(n_131) );
INVx5_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
BUFx3_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
INVx1_ASAP7_75t_L g222 ( .A(n_135), .Y(n_222) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_137), .Y(n_142) );
INVx3_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
AND2x2_ASAP7_75t_L g154 ( .A(n_137), .B(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
INVx1_ASAP7_75t_L g252 ( .A(n_137), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_143), .C(n_146), .Y(n_138) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_141), .A2(n_144), .B1(n_468), .B2(n_469), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_141), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_141), .B(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
INVx2_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_144), .B(n_243), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_144), .A2(n_184), .B(n_444), .C(n_445), .Y(n_443) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_145), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g455 ( .A(n_147), .Y(n_455) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_SL g161 ( .A1(n_149), .A2(n_162), .B(n_163), .C(n_164), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_149), .A2(n_163), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_149), .A2(n_163), .B(n_451), .C(n_452), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_149), .A2(n_163), .B(n_465), .C(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_149), .A2(n_163), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_149), .A2(n_163), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_SL g542 ( .A1(n_149), .A2(n_163), .B(n_543), .C(n_544), .Y(n_542) );
INVx4_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g153 ( .A(n_150), .B(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_150), .B(n_154), .Y(n_215) );
BUFx2_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
INVx1_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
AND2x2_ASAP7_75t_L g173 ( .A(n_158), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g263 ( .A(n_158), .Y(n_263) );
AND2x2_ASAP7_75t_L g349 ( .A(n_158), .B(n_262), .Y(n_349) );
AND2x2_ASAP7_75t_L g404 ( .A(n_158), .B(n_196), .Y(n_404) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_172), .Y(n_158) );
INVx2_ASAP7_75t_L g202 ( .A(n_163), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_168), .B(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g545 ( .A(n_169), .Y(n_545) );
INVx2_ASAP7_75t_L g479 ( .A(n_170), .Y(n_479) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
INVx1_ASAP7_75t_L g507 ( .A(n_171), .Y(n_507) );
INVx1_ASAP7_75t_L g321 ( .A(n_173), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_173), .B(n_197), .Y(n_368) );
INVx5_ASAP7_75t_L g262 ( .A(n_174), .Y(n_262) );
AND2x4_ASAP7_75t_L g283 ( .A(n_174), .B(n_263), .Y(n_283) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
AND2x2_ASAP7_75t_L g380 ( .A(n_174), .B(n_365), .Y(n_380) );
AND2x2_ASAP7_75t_L g383 ( .A(n_174), .B(n_198), .Y(n_383) );
OR2x6_ASAP7_75t_L g174 ( .A(n_175), .B(n_190), .Y(n_174) );
AOI21xp5_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_178), .B(n_187), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_182), .B(n_184), .Y(n_179) );
INVx2_ASAP7_75t_L g183 ( .A(n_181), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_183), .A2(n_204), .B(n_205), .C(n_206), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_183), .A2(n_206), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_183), .A2(n_477), .B(n_478), .C(n_479), .Y(n_476) );
O2A1O1Ixp5_ASAP7_75t_L g494 ( .A1(n_183), .A2(n_479), .B(n_495), .C(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_185), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_188), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g192 ( .A(n_189), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_189), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_189), .A2(n_228), .B(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_189), .A2(n_215), .B(n_441), .C(n_442), .Y(n_440) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_189), .A2(n_541), .B(n_548), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_192), .A2(n_491), .B(n_497), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_193), .B(n_263), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_193), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_197), .Y(n_194) );
AND2x2_ASAP7_75t_L g288 ( .A(n_195), .B(n_263), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_195), .B(n_198), .Y(n_306) );
INVx1_ASAP7_75t_L g326 ( .A(n_195), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_195), .B(n_262), .Y(n_371) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_195), .Y(n_413) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_196), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_197), .B(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_197), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_197), .A2(n_258), .B(n_319), .C(n_321), .Y(n_318) );
AND2x2_ASAP7_75t_L g325 ( .A(n_197), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g334 ( .A(n_197), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g338 ( .A(n_197), .B(n_262), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_197), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g353 ( .A(n_197), .B(n_263), .Y(n_353) );
AND2x2_ASAP7_75t_L g403 ( .A(n_197), .B(n_404), .Y(n_403) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g267 ( .A(n_198), .Y(n_267) );
AND2x2_ASAP7_75t_L g308 ( .A(n_198), .B(n_261), .Y(n_308) );
AND2x2_ASAP7_75t_L g320 ( .A(n_198), .B(n_295), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_198), .B(n_349), .Y(n_367) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_207), .Y(n_198) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_234), .Y(n_209) );
INVx1_ASAP7_75t_L g256 ( .A(n_210), .Y(n_256) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_226), .Y(n_210) );
OR2x2_ASAP7_75t_L g258 ( .A(n_211), .B(n_226), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g264 ( .A(n_211), .B(n_265), .C(n_266), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_211), .B(n_236), .Y(n_275) );
OR2x2_ASAP7_75t_L g290 ( .A(n_211), .B(n_278), .Y(n_290) );
AND2x2_ASAP7_75t_L g296 ( .A(n_211), .B(n_245), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_211), .B(n_427), .Y(n_426) );
INVx5_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_212), .B(n_236), .Y(n_293) );
AND2x2_ASAP7_75t_L g332 ( .A(n_212), .B(n_246), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_212), .B(n_245), .Y(n_360) );
OR2x2_ASAP7_75t_L g363 ( .A(n_212), .B(n_245), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_215), .A2(n_474), .B(n_475), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_215), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_220), .A2(n_251), .B(n_253), .Y(n_250) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g462 ( .A(n_225), .Y(n_462) );
INVx5_ASAP7_75t_SL g278 ( .A(n_226), .Y(n_278) );
OR2x2_ASAP7_75t_L g284 ( .A(n_226), .B(n_235), .Y(n_284) );
AND2x2_ASAP7_75t_L g300 ( .A(n_226), .B(n_301), .Y(n_300) );
AOI321xp33_ASAP7_75t_L g307 ( .A1(n_226), .A2(n_308), .A3(n_309), .B1(n_310), .B2(n_316), .C(n_318), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_226), .B(n_234), .Y(n_317) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_226), .Y(n_330) );
OR2x2_ASAP7_75t_L g377 ( .A(n_226), .B(n_275), .Y(n_377) );
AND2x2_ASAP7_75t_L g399 ( .A(n_226), .B(n_296), .Y(n_399) );
AND2x2_ASAP7_75t_L g418 ( .A(n_226), .B(n_236), .Y(n_418) );
OR2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
INVx1_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_245), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_236), .B(n_245), .Y(n_259) );
AND2x2_ASAP7_75t_L g268 ( .A(n_236), .B(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g295 ( .A(n_236), .Y(n_295) );
AND2x2_ASAP7_75t_L g301 ( .A(n_236), .B(n_296), .Y(n_301) );
INVxp67_ASAP7_75t_L g331 ( .A(n_236), .Y(n_331) );
OR2x2_ASAP7_75t_L g373 ( .A(n_236), .B(n_278), .Y(n_373) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_244), .Y(n_236) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_237), .A2(n_449), .B(n_456), .Y(n_448) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_237), .A2(n_501), .B(n_508), .Y(n_500) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_237), .A2(n_510), .B(n_516), .Y(n_509) );
OR2x2_ASAP7_75t_L g255 ( .A(n_245), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_SL g269 ( .A(n_245), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_245), .B(n_258), .Y(n_302) );
AND2x2_ASAP7_75t_L g351 ( .A(n_245), .B(n_295), .Y(n_351) );
AND2x2_ASAP7_75t_L g389 ( .A(n_245), .B(n_278), .Y(n_389) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_246), .B(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_257), .B(n_260), .C(n_264), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_255), .A2(n_257), .B1(n_382), .B2(n_384), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_257), .A2(n_280), .B1(n_335), .B2(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_SL g409 ( .A(n_258), .Y(n_409) );
INVx1_ASAP7_75t_SL g309 ( .A(n_259), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_261), .B(n_281), .Y(n_311) );
AOI222xp33_ASAP7_75t_L g322 ( .A1(n_261), .A2(n_302), .B1(n_309), .B2(n_323), .C1(n_327), .C2(n_333), .Y(n_322) );
AND2x2_ASAP7_75t_L g412 ( .A(n_261), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_262), .B(n_282), .Y(n_357) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_262), .Y(n_394) );
AND2x2_ASAP7_75t_L g397 ( .A(n_262), .B(n_306), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_262), .B(n_413), .Y(n_423) );
INVx1_ASAP7_75t_L g314 ( .A(n_263), .Y(n_314) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_263), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g405 ( .A1(n_265), .A2(n_406), .B(n_407), .C(n_410), .Y(n_405) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g328 ( .A(n_267), .B(n_329), .C(n_332), .Y(n_328) );
OR2x2_ASAP7_75t_L g356 ( .A(n_267), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_267), .B(n_283), .Y(n_384) );
OR2x2_ASAP7_75t_L g289 ( .A(n_269), .B(n_290), .Y(n_289) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_273), .B(n_279), .C(n_291), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_272), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g378 ( .A(n_273), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_274), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g292 ( .A(n_277), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_278), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g346 ( .A(n_278), .B(n_296), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_278), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_278), .B(n_295), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B1(n_285), .B2(n_289), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_281), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_283), .B(n_325), .Y(n_324) );
OAI221xp5_ASAP7_75t_SL g347 ( .A1(n_284), .A2(n_348), .B1(n_350), .B2(n_352), .C(n_354), .Y(n_347) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g402 ( .A(n_287), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g415 ( .A(n_287), .B(n_404), .Y(n_415) );
INVx1_ASAP7_75t_L g335 ( .A(n_288), .Y(n_335) );
INVx1_ASAP7_75t_L g406 ( .A(n_289), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_290), .A2(n_373), .B(n_396), .Y(n_395) );
AOI21xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B(n_297), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI21xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_303), .Y(n_299) );
INVx1_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_301), .A2(n_387), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_386) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_309), .A2(n_399), .B1(n_400), .B2(n_402), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g375 ( .A(n_311), .Y(n_375) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp67_ASAP7_75t_SL g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g379 ( .A(n_315), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g344 ( .A(n_320), .Y(n_344) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_325), .B(n_349), .Y(n_401) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_331), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g417 ( .A(n_332), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g424 ( .A(n_332), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI211xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_339), .B(n_340), .C(n_374), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B(n_347), .C(n_366), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g427 ( .A(n_351), .Y(n_427) );
AND2x2_ASAP7_75t_L g364 ( .A(n_353), .B(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_362), .B2(n_364), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
OR2x2_ASAP7_75t_L g372 ( .A(n_360), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g425 ( .A(n_361), .Y(n_425) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI31xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .A3(n_369), .B(n_372), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI211xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B(n_378), .C(n_381), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
CKINVDCx16_ASAP7_75t_R g382 ( .A(n_383), .Y(n_382) );
NAND5xp2_ASAP7_75t_L g385 ( .A(n_386), .B(n_398), .C(n_405), .D(n_419), .E(n_422), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_397), .A2(n_423), .B1(n_424), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_SL g421 ( .A(n_399), .Y(n_421) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .B(n_416), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g694 ( .A1(n_430), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_432), .Y(n_697) );
OR3x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_605), .C(n_652), .Y(n_432) );
NAND3xp33_ASAP7_75t_SL g433 ( .A(n_434), .B(n_551), .C(n_576), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_489), .B1(n_517), .B2(n_520), .C(n_528), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_457), .B(n_482), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_437), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_437), .B(n_533), .Y(n_649) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_448), .Y(n_437) );
AND2x2_ASAP7_75t_L g519 ( .A(n_438), .B(n_488), .Y(n_519) );
AND2x2_ASAP7_75t_L g569 ( .A(n_438), .B(n_487), .Y(n_569) );
AND2x2_ASAP7_75t_L g590 ( .A(n_438), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g595 ( .A(n_438), .B(n_562), .Y(n_595) );
OR2x2_ASAP7_75t_L g603 ( .A(n_438), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g675 ( .A(n_438), .B(n_471), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_438), .B(n_624), .Y(n_689) );
INVx3_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g534 ( .A(n_439), .B(n_448), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_439), .B(n_471), .Y(n_535) );
AND2x4_ASAP7_75t_L g557 ( .A(n_439), .B(n_488), .Y(n_557) );
AND2x2_ASAP7_75t_L g587 ( .A(n_439), .B(n_459), .Y(n_587) );
AND2x2_ASAP7_75t_L g596 ( .A(n_439), .B(n_586), .Y(n_596) );
AND2x2_ASAP7_75t_L g612 ( .A(n_439), .B(n_472), .Y(n_612) );
OR2x2_ASAP7_75t_L g621 ( .A(n_439), .B(n_604), .Y(n_621) );
AND2x2_ASAP7_75t_L g627 ( .A(n_439), .B(n_562), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_439), .B(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g641 ( .A(n_439), .B(n_484), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_439), .B(n_530), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_439), .B(n_591), .Y(n_680) );
OR2x6_ASAP7_75t_L g439 ( .A(n_440), .B(n_446), .Y(n_439) );
INVx2_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
AND2x2_ASAP7_75t_L g586 ( .A(n_448), .B(n_471), .Y(n_586) );
AND2x2_ASAP7_75t_L g591 ( .A(n_448), .B(n_472), .Y(n_591) );
INVx1_ASAP7_75t_L g647 ( .A(n_448), .Y(n_647) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g556 ( .A(n_458), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_471), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_459), .B(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g533 ( .A(n_459), .Y(n_533) );
OR2x2_ASAP7_75t_L g604 ( .A(n_459), .B(n_471), .Y(n_604) );
OR2x2_ASAP7_75t_L g665 ( .A(n_459), .B(n_572), .Y(n_665) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B(n_470), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_461), .A2(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g485 ( .A(n_463), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_470), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_471), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g624 ( .A(n_471), .B(n_484), .Y(n_624) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g563 ( .A(n_472), .Y(n_563) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_483), .A2(n_669), .B1(n_673), .B2(n_676), .C(n_677), .Y(n_668) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_SL g531 ( .A(n_484), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_484), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_484), .B(n_519), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_487), .B(n_533), .Y(n_655) );
AND2x2_ASAP7_75t_L g562 ( .A(n_488), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_SL g566 ( .A(n_489), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_489), .B(n_572), .Y(n_602) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
AND2x2_ASAP7_75t_L g527 ( .A(n_490), .B(n_500), .Y(n_527) );
INVx4_ASAP7_75t_L g539 ( .A(n_490), .Y(n_539) );
BUFx3_ASAP7_75t_L g582 ( .A(n_490), .Y(n_582) );
AND3x2_ASAP7_75t_L g597 ( .A(n_490), .B(n_598), .C(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g679 ( .A(n_499), .B(n_593), .Y(n_679) );
AND2x2_ASAP7_75t_L g687 ( .A(n_499), .B(n_572), .Y(n_687) );
INVx1_ASAP7_75t_SL g692 ( .A(n_499), .Y(n_692) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .Y(n_499) );
INVx1_ASAP7_75t_SL g550 ( .A(n_500), .Y(n_550) );
AND2x2_ASAP7_75t_L g573 ( .A(n_500), .B(n_539), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_500), .B(n_523), .Y(n_575) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_500), .Y(n_615) );
OR2x2_ASAP7_75t_L g620 ( .A(n_500), .B(n_539), .Y(n_620) );
INVx2_ASAP7_75t_L g525 ( .A(n_509), .Y(n_525) );
AND2x2_ASAP7_75t_L g560 ( .A(n_509), .B(n_540), .Y(n_560) );
OR2x2_ASAP7_75t_L g580 ( .A(n_509), .B(n_540), .Y(n_580) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_509), .Y(n_600) );
INVx1_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_518), .A2(n_559), .B(n_651), .Y(n_650) );
AOI322xp5_ASAP7_75t_L g686 ( .A1(n_520), .A2(n_530), .A3(n_557), .B1(n_687), .B2(n_688), .C1(n_690), .C2(n_693), .Y(n_686) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_522), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_523), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g549 ( .A(n_524), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g617 ( .A(n_525), .B(n_539), .Y(n_617) );
AND2x2_ASAP7_75t_L g684 ( .A(n_525), .B(n_540), .Y(n_684) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g625 ( .A(n_527), .B(n_579), .Y(n_625) );
AOI31xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .A3(n_535), .B(n_536), .Y(n_528) );
AND2x2_ASAP7_75t_L g584 ( .A(n_530), .B(n_562), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_530), .B(n_554), .Y(n_666) );
AND2x2_ASAP7_75t_L g685 ( .A(n_530), .B(n_590), .Y(n_685) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_533), .B(n_562), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g608 ( .A(n_533), .B(n_591), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_533), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_533), .B(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_534), .B(n_591), .Y(n_623) );
INVx1_ASAP7_75t_L g667 ( .A(n_534), .Y(n_667) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_549), .Y(n_537) );
INVxp67_ASAP7_75t_L g619 ( .A(n_538), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_539), .B(n_550), .Y(n_555) );
INVx1_ASAP7_75t_L g661 ( .A(n_539), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_539), .B(n_638), .Y(n_672) );
BUFx3_ASAP7_75t_L g572 ( .A(n_540), .Y(n_572) );
AND2x2_ASAP7_75t_L g598 ( .A(n_540), .B(n_550), .Y(n_598) );
INVx2_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_549), .B(n_671), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_556), .B(n_558), .C(n_567), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI21xp33_ASAP7_75t_L g601 ( .A1(n_553), .A2(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_554), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_554), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g634 ( .A(n_555), .B(n_580), .Y(n_634) );
INVx3_ASAP7_75t_L g565 ( .A(n_557), .Y(n_565) );
OAI22xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_561), .B1(n_564), .B2(n_566), .Y(n_558) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_560), .A2(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g609 ( .A(n_560), .B(n_573), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_560), .B(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g564 ( .A(n_563), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g633 ( .A(n_563), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g577 ( .A1(n_564), .A2(n_578), .B(n_583), .Y(n_577) );
OAI22xp33_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_570), .B1(n_574), .B2(n_575), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_569), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g593 ( .A(n_572), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_572), .B(n_615), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_588), .C(n_601), .Y(n_576) );
OAI22xp5_ASAP7_75t_SL g643 ( .A1(n_578), .A2(n_644), .B1(n_648), .B2(n_649), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g648 ( .A(n_580), .B(n_581), .Y(n_648) );
AND2x2_ASAP7_75t_L g656 ( .A(n_581), .B(n_637), .Y(n_656) );
CKINVDCx16_ASAP7_75t_R g581 ( .A(n_582), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_SL g664 ( .A1(n_582), .A2(n_665), .B(n_666), .C(n_667), .Y(n_664) );
OR2x2_ASAP7_75t_L g691 ( .A(n_582), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B(n_594), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_590), .A2(n_627), .B(n_628), .C(n_631), .Y(n_626) );
OAI21xp33_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_596), .B(n_597), .Y(n_594) );
AND2x2_ASAP7_75t_L g659 ( .A(n_598), .B(n_617), .Y(n_659) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g637 ( .A(n_600), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g642 ( .A(n_602), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g605 ( .A(n_606), .B(n_626), .C(n_639), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B(n_610), .C(n_618), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g676 ( .A(n_613), .Y(n_676) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g636 ( .A(n_615), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_615), .B(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_621), .C(n_622), .Y(n_618) );
INVx2_ASAP7_75t_SL g630 ( .A(n_620), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_621), .A2(n_632), .B1(n_634), .B2(n_635), .Y(n_631) );
OAI21xp33_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_624), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B(n_643), .C(n_650), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVxp33_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g693 ( .A(n_647), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_668), .C(n_681), .D(n_686), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_656), .B(n_657), .C(n_664), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B(n_662), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_658), .A2(n_678), .B(n_680), .Y(n_677) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_665), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g706 ( .A(n_704), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_710), .Y(n_716) );
OR2x2_ASAP7_75t_SL g710 ( .A(n_711), .B(n_715), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
endmodule