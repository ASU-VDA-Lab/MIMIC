module fake_jpeg_22862_n_193 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_2),
.B(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_36),
.B(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_44),
.B1(n_41),
.B2(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_44),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_21),
.B1(n_30),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_56),
.B1(n_62),
.B2(n_69),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_31),
.C(n_11),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_31),
.C(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_39),
.B1(n_21),
.B2(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_16),
.B1(n_6),
.B2(n_7),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_20),
.B1(n_23),
.B2(n_30),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_23),
.B(n_27),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_16),
.B(n_33),
.C(n_24),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_70),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_22),
.B1(n_27),
.B2(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_4),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_16),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_3),
.Y(n_74)
);

OAI22x1_ASAP7_75t_SL g75 ( 
.A1(n_34),
.A2(n_33),
.B1(n_17),
.B2(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_94),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_25),
.A3(n_24),
.B1(n_18),
.B2(n_47),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_58),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_22),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_66),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_47),
.B1(n_33),
.B2(n_17),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_49),
.B1(n_70),
.B2(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_89),
.B1(n_96),
.B2(n_99),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_3),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_8),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_93),
.B(n_95),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_16),
.B(n_8),
.C(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_49),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_72),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_8),
.B1(n_10),
.B2(n_58),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_67),
.C(n_71),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_113),
.C(n_115),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_59),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_67),
.C(n_68),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_63),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_68),
.B(n_58),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_92),
.B(n_83),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_85),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_79),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_61),
.C(n_10),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_87),
.C(n_103),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

NOR4xp25_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.D(n_110),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_87),
.C(n_82),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_120),
.B1(n_123),
.B2(n_89),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_87),
.C(n_82),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_144),
.A2(n_110),
.B(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_156),
.C(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_143),
.B1(n_127),
.B2(n_90),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_138),
.B1(n_140),
.B2(n_139),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_115),
.B(n_106),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_157),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_121),
.C(n_88),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_141),
.B(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_158),
.B1(n_146),
.B2(n_145),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_161),
.C(n_169),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_137),
.C(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_166),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_134),
.A3(n_107),
.B1(n_81),
.B2(n_137),
.C1(n_108),
.C2(n_78),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_165),
.A2(n_90),
.B1(n_153),
.B2(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_137),
.C(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_145),
.B(n_153),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_156),
.B1(n_129),
.B2(n_91),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_177),
.C(n_61),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_154),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_159),
.A3(n_161),
.B1(n_163),
.B2(n_164),
.C1(n_160),
.C2(n_129),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_181),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_182),
.B(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_80),
.B1(n_88),
.B2(n_121),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_61),
.B1(n_12),
.B2(n_14),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_187),
.Y(n_188)
);

AOI221xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_182),
.B1(n_179),
.B2(n_177),
.C(n_171),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_190),
.C(n_14),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_171),
.B(n_12),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_192),
.Y(n_193)
);


endmodule