module fake_jpeg_2791_n_223 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_223);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_16),
.B(n_40),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_21),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_83),
.Y(n_90)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_68),
.Y(n_94)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_66),
.B1(n_56),
.B2(n_67),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_67),
.B1(n_56),
.B2(n_70),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_101),
.B1(n_88),
.B2(n_65),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_103),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_92),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_55),
.B1(n_74),
.B2(n_72),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_117),
.B1(n_63),
.B2(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_60),
.Y(n_109)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_57),
.B1(n_59),
.B2(n_54),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_116),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_115),
.C(n_121),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_74),
.B1(n_72),
.B2(n_65),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_62),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_77),
.A3(n_57),
.B1(n_59),
.B2(n_54),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_101),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_1),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_126),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_58),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_88),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_6),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_63),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_136),
.B(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_138),
.A2(n_144),
.B1(n_140),
.B2(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_2),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_141),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_120),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_2),
.B(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_5),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_160),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_110),
.B1(n_23),
.B2(n_25),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_153),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_135),
.B1(n_132),
.B2(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_162),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_52),
.B1(n_46),
.B2(n_45),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_159),
.B(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_42),
.B1(n_39),
.B2(n_35),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_6),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_137),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_12),
.B(n_13),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_7),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_123),
.B(n_8),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_11),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_20),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_179),
.C(n_182),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_9),
.B(n_10),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_188),
.B(n_147),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_154),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_181),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_9),
.C(n_10),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_169),
.B(n_19),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_11),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_187),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_12),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_13),
.C(n_15),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_194),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_156),
.B1(n_168),
.B2(n_163),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_197),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_186),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_198),
.A2(n_185),
.B(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_180),
.B(n_183),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_203),
.B(n_194),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_174),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_146),
.C(n_182),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_196),
.C(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_207),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_189),
.B1(n_164),
.B2(n_185),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_201),
.B1(n_166),
.B2(n_205),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_213),
.C(n_211),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_209),
.C(n_211),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_218),
.A2(n_217),
.B(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_219),
.B(n_193),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_179),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_15),
.Y(n_223)
);


endmodule