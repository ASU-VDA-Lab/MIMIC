module fake_jpeg_21910_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_8),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_30),
.B(n_26),
.C(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_15),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_57),
.C(n_24),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_31),
.B1(n_17),
.B2(n_22),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_29),
.B(n_23),
.C(n_16),
.Y(n_85)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_56),
.B1(n_40),
.B2(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_56)
);

NOR3xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_25),
.C(n_27),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_85),
.B1(n_48),
.B2(n_63),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_35),
.C(n_33),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_86),
.B1(n_25),
.B2(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_98),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_68),
.C(n_52),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_60),
.B(n_15),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_71),
.B1(n_51),
.B2(n_55),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_48),
.B1(n_59),
.B2(n_53),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_72),
.B1(n_70),
.B2(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_99),
.Y(n_126)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_37),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_45),
.B1(n_51),
.B2(n_18),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_15),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_106),
.B(n_87),
.Y(n_113)
);

NAND2x1_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_62),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_47),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_124),
.B1(n_102),
.B2(n_110),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_118),
.B(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_32),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_129),
.C(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_119),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_0),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_128),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_53),
.B1(n_39),
.B2(n_35),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_106),
.B(n_93),
.C(n_89),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_130),
.B1(n_132),
.B2(n_96),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_27),
.C(n_28),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_35),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_91),
.A2(n_39),
.B1(n_77),
.B2(n_28),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_105),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_136),
.B(n_140),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_99),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_146),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_95),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_150),
.C(n_60),
.Y(n_177)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_147),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_149),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_108),
.C(n_100),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_118),
.B(n_112),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_15),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_112),
.B1(n_104),
.B2(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_37),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_172),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_133),
.B(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_147),
.B1(n_144),
.B2(n_141),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_0),
.Y(n_167)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_116),
.B(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_145),
.C(n_150),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_184),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_190),
.C(n_195),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

BUFx12f_ASAP7_75t_SL g186 ( 
.A(n_175),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_186),
.A2(n_161),
.B(n_164),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_197),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_139),
.C(n_137),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_152),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_159),
.B(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_166),
.B1(n_167),
.B2(n_176),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_138),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_168),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_165),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_189),
.C(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_173),
.B1(n_162),
.B2(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_210),
.B1(n_179),
.B2(n_192),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_202),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_135),
.B(n_140),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_185),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_183),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_171),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_211),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_136),
.C(n_167),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_184),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_182),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_218),
.C(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_220),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_183),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_202),
.B(n_181),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_189),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_207),
.B(n_203),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_228),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_200),
.B1(n_181),
.B2(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_229),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_201),
.B(n_199),
.Y(n_229)
);

NAND2x1p5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_205),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_230),
.A2(n_234),
.B(n_219),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_29),
.B1(n_23),
.B2(n_15),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_29),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_9),
.B(n_1),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_237),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_213),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_239),
.C(n_225),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_10),
.B(n_2),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_23),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_14),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_7),
.C(n_3),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_246),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_5),
.C(n_6),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_250),
.B(n_13),
.Y(n_251)
);

FAx1_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_11),
.CI(n_12),
.CON(n_248),
.SN(n_248)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_249),
.B(n_13),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_252),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_13),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_14),
.B(n_0),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_255),
.Y(n_256)
);


endmodule