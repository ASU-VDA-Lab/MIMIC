module real_jpeg_14218_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_0),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_26),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_5),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_18),
.B1(n_19),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_29),
.B1(n_52),
.B2(n_53),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_9),
.B(n_24),
.C(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_9),
.B(n_88),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_9),
.A2(n_20),
.B(n_23),
.C(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_9),
.B(n_37),
.C(n_40),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_9),
.B(n_91),
.Y(n_135)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_107),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_105),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_93),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_14),
.B(n_93),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_14),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_60),
.CI(n_77),
.CON(n_14),
.SN(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_32),
.C(n_46),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_16),
.A2(n_32),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_16),
.A2(n_71),
.B1(n_76),
.B2(n_98),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B(n_27),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_18),
.A2(n_19),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_18),
.A2(n_21),
.B(n_29),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_19),
.B(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_28),
.A2(n_30),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_29),
.B(n_64),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_29),
.B(n_43),
.Y(n_147)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_43),
.B(n_44),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_45),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g124 ( 
.A1(n_34),
.A2(n_38),
.B1(n_45),
.B2(n_73),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_39),
.B(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_72),
.B(n_74),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_47),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OA21x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_56),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_81),
.Y(n_80)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_58),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_64),
.B(n_66),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_68),
.B1(n_70),
.B2(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_66),
.B(n_83),
.Y(n_102)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_98),
.C(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_71),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_71),
.A2(n_76),
.B1(n_131),
.B2(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_82),
.A2(n_100),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_82),
.B(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_124),
.C(n_136),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_92),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_102),
.C(n_103),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.C(n_101),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_101),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_158),
.B(n_162),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_127),
.B(n_157),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_117),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_110),
.B(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_112),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_124),
.C(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_123),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_126),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_151),
.B(n_156),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_138),
.B(n_150),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_142),
.B(n_149),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B(n_148),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);


endmodule