module fake_jpeg_29064_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx11_ASAP7_75t_SL g77 ( 
.A(n_75),
.Y(n_77)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_21),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_85),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

OR2x2_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_0),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_68),
.B1(n_60),
.B2(n_76),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_99),
.B1(n_55),
.B2(n_71),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_57),
.B1(n_70),
.B2(n_66),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_68),
.B1(n_57),
.B2(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_74),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_84),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_112),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_72),
.B(n_64),
.C(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_3),
.Y(n_122)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_55),
.B1(n_73),
.B2(n_75),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_114),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_2),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_89),
.B1(n_88),
.B2(n_67),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_61),
.B(n_56),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_4),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_1),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_118),
.Y(n_131)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_1),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_86),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_130),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_136),
.B1(n_120),
.B2(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_36),
.B1(n_50),
.B2(n_48),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_7),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_9),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_140),
.B(n_10),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_37),
.C(n_47),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_143),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_106),
.B(n_31),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_43),
.B(n_24),
.Y(n_167)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_52),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_150),
.C(n_131),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_152),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_154),
.B(n_13),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_38),
.C(n_45),
.Y(n_150)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_151),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_124),
.B(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_42),
.C(n_20),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_29),
.C(n_40),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_170),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_154),
.C(n_157),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_153),
.C(n_150),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_152),
.B1(n_145),
.B2(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_161),
.B1(n_165),
.B2(n_149),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_161),
.B1(n_165),
.B2(n_158),
.Y(n_179)
);

AOI321xp33_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_162),
.A3(n_146),
.B1(n_178),
.B2(n_175),
.C(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_172),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_174),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_182),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_156),
.B1(n_125),
.B2(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_159),
.C(n_44),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_46),
.Y(n_186)
);


endmodule