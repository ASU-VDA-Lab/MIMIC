module real_jpeg_33206_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g171 ( 
.A(n_0),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_0),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g374 ( 
.A(n_0),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_0),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_0),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_1),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_2),
.B(n_159),
.Y(n_158)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_2),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_2),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_2),
.B(n_283),
.Y(n_282)
);

NAND2x1_ASAP7_75t_L g371 ( 
.A(n_2),
.B(n_372),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_15),
.B1(n_21),
.B2(n_24),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_4),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_4),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_4),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_4),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_4),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_4),
.B(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_4),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_4),
.B(n_421),
.Y(n_420)
);

AND2x4_ASAP7_75t_SL g191 ( 
.A(n_5),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_129),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_5),
.B(n_195),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g428 ( 
.A(n_5),
.B(n_429),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_5),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_5),
.B(n_261),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_5),
.B(n_357),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_5),
.B(n_564),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_6),
.B(n_222),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_6),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_6),
.B(n_403),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_6),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_6),
.B(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_6),
.B(n_530),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_6),
.B(n_537),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_7),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_7),
.B(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_7),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_7),
.B(n_170),
.Y(n_169)
);

NAND2x1p5_ASAP7_75t_L g182 ( 
.A(n_7),
.B(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_9),
.Y(n_409)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_10),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_10),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_10),
.Y(n_262)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_10),
.Y(n_438)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_11),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_12),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_12),
.B(n_39),
.Y(n_209)
);

AND2x4_ASAP7_75t_SL g227 ( 
.A(n_12),
.B(n_228),
.Y(n_227)
);

AND2x4_ASAP7_75t_SL g256 ( 
.A(n_12),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_12),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_12),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_12),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_12),
.B(n_357),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_13),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_13),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_13),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_13),
.B(n_222),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_13),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_13),
.B(n_510),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_13),
.B(n_353),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_14),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_14),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_14),
.B(n_368),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_14),
.B(n_44),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_14),
.B(n_411),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_14),
.B(n_478),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_14),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_14),
.B(n_522),
.Y(n_521)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_16),
.B(n_67),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g194 ( 
.A(n_16),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_16),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_16),
.B(n_416),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_16),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_16),
.B(n_560),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_17),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_17),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_18),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_18),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_19),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_19),
.B(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_19),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_19),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_19),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_19),
.B(n_287),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_138),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_137),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_120),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_27),
.B(n_120),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_91),
.C(n_93),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_29),
.B(n_328),
.Y(n_327)
);

MAJx2_ASAP7_75t_R g29 ( 
.A(n_30),
.B(n_60),
.C(n_77),
.Y(n_29)
);

XNOR2x1_ASAP7_75t_L g334 ( 
.A(n_30),
.B(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_48),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_49),
.C(n_55),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.C(n_43),
.Y(n_31)
);

XNOR2x1_ASAP7_75t_L g320 ( 
.A(n_32),
.B(n_43),
.Y(n_320)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_37),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_37),
.Y(n_404)
);

XOR2x1_ASAP7_75t_L g319 ( 
.A(n_38),
.B(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_47),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_47),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_54),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_60),
.B(n_336),
.Y(n_335)
);

XOR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_62),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_62),
.A2(n_70),
.B1(n_87),
.B2(n_297),
.Y(n_311)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_69),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_86),
.C(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_76),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_78),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.C(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_80),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_87),
.A2(n_182),
.B1(n_186),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_87),
.Y(n_297)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_90),
.Y(n_533)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_92),
.B(n_94),
.Y(n_328)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_103),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_106),
.C(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_101),
.Y(n_379)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_108),
.C(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_109),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_114),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_119),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_135),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21x1_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_342),
.B(n_627),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_326),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_298),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_142),
.B(n_298),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_213),
.C(n_269),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_144),
.A2(n_145),
.B1(n_270),
.B2(n_607),
.Y(n_606)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_187),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_146),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_162),
.C(n_176),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_148),
.B(n_611),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_150),
.B(n_157),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_150),
.B(n_157),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_153),
.Y(n_400)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_153),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_153),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_156),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_160),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_161),
.Y(n_413)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_162),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.C(n_172),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_164),
.B(n_169),
.Y(n_236)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_166),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_167),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_169),
.B1(n_182),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_178),
.C(n_182),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_169),
.B(n_178),
.C(n_182),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_170),
.Y(n_538)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_172),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_242)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_176),
.B(n_610),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_185),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_186),
.B(n_291),
.C(n_297),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_207),
.B1(n_211),
.B2(n_212),
.Y(n_187)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_201),
.C(n_203),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.C(n_197),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_194),
.C(n_197),
.Y(n_246)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_198),
.Y(n_218)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_194),
.B(n_218),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g322 ( 
.A(n_203),
.B(n_323),
.C(n_324),
.Y(n_322)
);

INVx3_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_205),
.Y(n_564)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_206),
.Y(n_370)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_207),
.Y(n_302)
);

XOR2x1_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_209),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_211),
.Y(n_301)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_214),
.B(n_606),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_243),
.C(n_247),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_216),
.B(n_616),
.Y(n_615)
);

AO22x1_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_219),
.B1(n_239),
.B2(n_242),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_234),
.C(n_237),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_226),
.C(n_230),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_221),
.A2(n_226),
.B1(n_227),
.B2(n_241),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_231),
.C(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_230),
.B(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_236),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g585 ( 
.A(n_240),
.B(n_242),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_243),
.B(n_248),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.C(n_258),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22x1_ASAP7_75t_L g592 ( 
.A1(n_250),
.A2(n_256),
.B1(n_593),
.B2(n_594),
.Y(n_592)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_250),
.Y(n_594)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_255),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_256),
.Y(n_593)
);

XNOR2x1_ASAP7_75t_L g591 ( 
.A(n_258),
.B(n_592),
.Y(n_591)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.C(n_267),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_574)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_266),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_267),
.B(n_574),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_270),
.Y(n_607)
);

XOR2x1_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_289),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_272)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_308),
.C(n_309),
.Y(n_307)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_286),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_314),
.C(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_314),
.C(n_315),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_303),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_304),
.C(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.C(n_302),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_312),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_316),
.B1(n_317),
.B2(n_325),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_322),
.C(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_318),
.Y(n_331)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_329),
.B(n_337),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_327),
.B(n_329),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_327),
.B(n_329),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.C(n_333),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_341),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_334),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_337),
.A2(n_629),
.B(n_630),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_338),
.B(n_340),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_603),
.B(n_624),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_550),
.B(n_601),
.Y(n_343)
);

OAI21x1_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_465),
.B(n_548),
.Y(n_344)
);

NOR3xp33_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_446),
.C(n_449),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_347),
.B(n_447),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_391),
.Y(n_347)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_348),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_348),
.B(n_599),
.C(n_600),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_365),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_349),
.B(n_366),
.C(n_376),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_358),
.C(n_363),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_350),
.B(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_351),
.A2(n_352),
.B1(n_355),
.B2(n_356),
.Y(n_453)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_358),
.A2(n_359),
.B1(n_363),
.B2(n_364),
.Y(n_464)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_376),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_371),
.B(n_375),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_371),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx8_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_375),
.A2(n_576),
.B1(n_577),
.B2(n_578),
.Y(n_575)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_375),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_SL g587 ( 
.A(n_375),
.B(n_573),
.C(n_577),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_380),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_378),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_385),
.B1(n_389),
.B2(n_390),
.Y(n_380)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_381),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_381),
.B(n_389),
.C(n_557),
.Y(n_556)
);

INVx3_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_383),
.Y(n_513)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_384),
.Y(n_475)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_385),
.Y(n_389)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_388),
.Y(n_562)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_425),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_393),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.C(n_414),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_394),
.B(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_397),
.C(n_398),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_401),
.B(n_414),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_405),
.C(n_410),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_402),
.B(n_405),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_409),
.Y(n_485)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_419),
.B1(n_420),
.B2(n_424),
.Y(n_414)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_415),
.Y(n_424)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_424),
.Y(n_442)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_425),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_441),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g553 ( 
.A(n_426),
.B(n_442),
.C(n_445),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_428),
.B(n_434),
.C(n_439),
.Y(n_576)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_434),
.B1(n_439),
.B2(n_440),
.Y(n_432)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_433),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_434),
.Y(n_440)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_444),
.B2(n_445),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_442),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_443),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_449),
.B(n_549),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.C(n_462),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_450),
.B(n_546),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_452),
.B(n_463),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.C(n_457),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_454),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_494),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

AO22x1_ASAP7_75t_SL g491 ( 
.A1(n_458),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_491)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_543),
.B(n_547),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_504),
.B(n_542),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_492),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_468),
.B(n_492),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_486),
.C(n_491),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_469),
.A2(n_470),
.B1(n_515),
.B2(n_517),
.Y(n_514)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_476),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_498),
.C(n_499),
.Y(n_497)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_481),
.Y(n_476)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_477),
.Y(n_499)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_481),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_483),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_486),
.A2(n_487),
.B1(n_491),
.B2(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_490),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_491),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_495),
.B1(n_496),
.B2(n_503),
.Y(n_492)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_493),
.Y(n_503)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_500),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_497),
.B(n_500),
.C(n_503),
.Y(n_544)
);

XOR2x1_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

AOI21x1_ASAP7_75t_SL g504 ( 
.A1(n_505),
.A2(n_518),
.B(n_541),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_514),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_SL g541 ( 
.A(n_506),
.B(n_514),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.C(n_511),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_526),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_508),
.A2(n_509),
.B1(n_511),
.B2(n_512),
.Y(n_526)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_515),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_519),
.A2(n_527),
.B(n_540),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_525),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_520),
.B(n_525),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_521),
.B(n_524),
.Y(n_534)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_524),
.B(n_536),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_535),
.B(n_539),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_534),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_534),
.Y(n_539)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_SL g543 ( 
.A(n_544),
.B(n_545),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_545),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_551),
.A2(n_579),
.B(n_595),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_551),
.B(n_579),
.C(n_602),
.Y(n_601)
);

MAJx2_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_569),
.C(n_571),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_552),
.B(n_597),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_553),
.B(n_554),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_553),
.B(n_555),
.C(n_581),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_567),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_558),
.Y(n_555)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_556),
.A2(n_563),
.B(n_566),
.C(n_590),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_559),
.A2(n_563),
.B1(n_565),
.B2(n_566),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_559),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_565),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_561),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_563),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_567),
.Y(n_581)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_570),
.B(n_572),
.Y(n_597)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_575),
.Y(n_572)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_576),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_582),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_580),
.B(n_619),
.C(n_620),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_586),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_583),
.Y(n_620)
);

XNOR2x1_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_585),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_586),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_587),
.B(n_588),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_R g612 ( 
.A(n_587),
.B(n_613),
.C(n_614),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_587),
.B(n_613),
.C(n_614),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_591),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_589),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_591),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_598),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_598),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_604),
.B(n_617),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_604),
.A2(n_625),
.B(n_626),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_608),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_608),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_609),
.B(n_612),
.C(n_615),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_609),
.B(n_623),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_622),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_621),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_618),
.B(n_621),
.Y(n_625)
);

OAI21x1_ASAP7_75t_SL g627 ( 
.A1(n_628),
.A2(n_631),
.B(n_632),
.Y(n_627)
);


endmodule