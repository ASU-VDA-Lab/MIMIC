module real_aes_7894_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g499 ( .A(n_1), .Y(n_499) );
INVx1_ASAP7_75t_L g180 ( .A(n_2), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_3), .A2(n_38), .B1(n_142), .B2(n_441), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g121 ( .A1(n_4), .A2(n_122), .B(n_129), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_5), .B(n_115), .Y(n_490) );
AND2x6_ASAP7_75t_L g127 ( .A(n_6), .B(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_7), .A2(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_8), .B(n_39), .Y(n_105) );
INVx1_ASAP7_75t_L g139 ( .A(n_9), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_10), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_12), .B(n_152), .Y(n_436) );
INVx1_ASAP7_75t_L g227 ( .A(n_13), .Y(n_227) );
INVx1_ASAP7_75t_L g494 ( .A(n_14), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_15), .B(n_116), .Y(n_475) );
AO32x2_ASAP7_75t_L g456 ( .A1(n_16), .A2(n_115), .A3(n_149), .B1(n_457), .B2(n_461), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_17), .B(n_142), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_18), .B(n_168), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_19), .B(n_116), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_20), .A2(n_49), .B1(n_142), .B2(n_441), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_21), .B(n_122), .Y(n_192) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_22), .A2(n_74), .B1(n_142), .B2(n_152), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_23), .B(n_142), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_24), .B(n_113), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_25), .A2(n_225), .B(n_226), .C(n_228), .Y(n_224) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_26), .A2(n_100), .B1(n_708), .B2(n_715), .C1(n_716), .C2(n_719), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_26), .Y(n_715) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_27), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_28), .B(n_145), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_29), .B(n_137), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_30), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_31), .Y(n_719) );
INVx1_ASAP7_75t_L g158 ( .A(n_32), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_33), .B(n_145), .Y(n_454) );
INVx2_ASAP7_75t_L g125 ( .A(n_34), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_35), .B(n_142), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_36), .B(n_145), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_37), .A2(n_127), .B(n_132), .C(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g156 ( .A(n_40), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_41), .B(n_137), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_42), .B(n_142), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_43), .A2(n_84), .B1(n_199), .B2(n_441), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_44), .B(n_142), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_45), .B(n_142), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g159 ( .A(n_46), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_47), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_48), .B(n_122), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_50), .A2(n_59), .B1(n_142), .B2(n_152), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_51), .A2(n_132), .B1(n_152), .B2(n_154), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_52), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_53), .B(n_142), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_54), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_55), .B(n_142), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_56), .A2(n_136), .B(n_138), .C(n_141), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_57), .Y(n_245) );
INVx1_ASAP7_75t_L g130 ( .A(n_58), .Y(n_130) );
INVx1_ASAP7_75t_L g128 ( .A(n_60), .Y(n_128) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_61), .A2(n_99), .B1(n_720), .B2(n_729), .C1(n_742), .C2(n_748), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_61), .A2(n_732), .B1(n_733), .B2(n_735), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_61), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_62), .B(n_142), .Y(n_500) );
INVx1_ASAP7_75t_L g119 ( .A(n_63), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_64), .Y(n_725) );
AO32x2_ASAP7_75t_L g466 ( .A1(n_65), .A2(n_115), .A3(n_207), .B1(n_461), .B2(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g511 ( .A(n_66), .Y(n_511) );
INVx1_ASAP7_75t_L g449 ( .A(n_67), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_68), .A2(n_141), .B(n_168), .C(n_169), .Y(n_167) );
INVxp67_ASAP7_75t_L g170 ( .A(n_69), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_70), .B(n_152), .Y(n_450) );
INVx1_ASAP7_75t_L g724 ( .A(n_71), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_72), .Y(n_162) );
INVx1_ASAP7_75t_L g238 ( .A(n_73), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_75), .A2(n_127), .B(n_132), .C(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_76), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_77), .B(n_152), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_78), .B(n_181), .Y(n_195) );
INVx2_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_80), .B(n_168), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_81), .B(n_152), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_82), .A2(n_127), .B(n_132), .C(n_179), .Y(n_178) );
OR2x2_ASAP7_75t_L g102 ( .A(n_83), .B(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g425 ( .A(n_83), .Y(n_425) );
OR2x2_ASAP7_75t_L g728 ( .A(n_83), .B(n_718), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_85), .A2(n_97), .B1(n_152), .B2(n_153), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_86), .B(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_87), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_88), .A2(n_127), .B(n_132), .C(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_89), .Y(n_217) );
INVx1_ASAP7_75t_L g166 ( .A(n_90), .Y(n_166) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_91), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_92), .B(n_181), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_93), .B(n_152), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_94), .B(n_115), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_95), .A2(n_122), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_96), .B(n_724), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_106), .B1(n_423), .B2(n_426), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g711 ( .A(n_102), .Y(n_711) );
OR2x2_ASAP7_75t_L g424 ( .A(n_103), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g718 ( .A(n_103), .Y(n_718) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx1_ASAP7_75t_L g734 ( .A(n_106), .Y(n_734) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g712 ( .A(n_107), .Y(n_712) );
AND3x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_345), .C(n_390), .Y(n_107) );
NOR4xp25_ASAP7_75t_L g108 ( .A(n_109), .B(n_268), .C(n_309), .D(n_326), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_172), .B(n_188), .C(n_230), .Y(n_109) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_146), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_111), .B(n_173), .Y(n_172) );
NOR4xp25_ASAP7_75t_L g292 ( .A(n_111), .B(n_286), .C(n_293), .D(n_299), .Y(n_292) );
AND2x2_ASAP7_75t_L g365 ( .A(n_111), .B(n_254), .Y(n_365) );
AND2x2_ASAP7_75t_L g384 ( .A(n_111), .B(n_330), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_111), .B(n_379), .Y(n_393) );
AND2x2_ASAP7_75t_L g406 ( .A(n_111), .B(n_187), .Y(n_406) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_SL g251 ( .A(n_112), .Y(n_251) );
AND2x2_ASAP7_75t_L g258 ( .A(n_112), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g308 ( .A(n_112), .B(n_147), .Y(n_308) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_112), .B(n_254), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_112), .B(n_147), .Y(n_323) );
AND2x2_ASAP7_75t_L g332 ( .A(n_112), .B(n_257), .Y(n_332) );
BUFx2_ASAP7_75t_L g355 ( .A(n_112), .Y(n_355) );
AND2x2_ASAP7_75t_L g359 ( .A(n_112), .B(n_163), .Y(n_359) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_121), .B(n_144), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_SL g201 ( .A(n_114), .B(n_202), .Y(n_201) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_114), .B(n_461), .C(n_477), .Y(n_476) );
AO21x1_ASAP7_75t_L g514 ( .A1(n_114), .A2(n_477), .B(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_115), .A2(n_164), .B(n_171), .Y(n_163) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_115), .A2(n_482), .B(n_490), .Y(n_481) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_117), .B(n_118), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
BUFx2_ASAP7_75t_L g221 ( .A(n_122), .Y(n_221) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_127), .Y(n_122) );
NAND2x1p5_ASAP7_75t_L g160 ( .A(n_123), .B(n_127), .Y(n_160) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g489 ( .A(n_124), .Y(n_489) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
INVx1_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx1_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_126), .Y(n_137) );
INVx3_ASAP7_75t_L g140 ( .A(n_126), .Y(n_140) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
INVx1_ASAP7_75t_L g168 ( .A(n_126), .Y(n_168) );
INVx4_ASAP7_75t_SL g143 ( .A(n_127), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_127), .A2(n_434), .B(n_438), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_127), .A2(n_448), .B(n_451), .Y(n_447) );
BUFx3_ASAP7_75t_L g461 ( .A(n_127), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_127), .A2(n_483), .B(n_486), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_127), .A2(n_493), .B(n_497), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_135), .C(n_143), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_131), .A2(n_143), .B(n_166), .C(n_167), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_131), .A2(n_143), .B(n_223), .C(n_224), .Y(n_222) );
INVx5_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_133), .Y(n_142) );
BUFx3_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
INVx1_ASAP7_75t_L g441 ( .A(n_133), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_136), .A2(n_439), .B(n_440), .Y(n_438) );
O2A1O1Ixp5_ASAP7_75t_L g510 ( .A1(n_136), .A2(n_498), .B(n_511), .C(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx4_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_137), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g467 ( .A1(n_137), .A2(n_140), .B1(n_468), .B2(n_469), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_137), .A2(n_459), .B1(n_478), .B2(n_479), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_140), .B(n_170), .Y(n_169) );
INVx5_ASAP7_75t_L g181 ( .A(n_140), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_SL g448 ( .A1(n_141), .A2(n_181), .B(n_449), .C(n_450), .Y(n_448) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g150 ( .A1(n_143), .A2(n_151), .B1(n_159), .B2(n_160), .Y(n_150) );
INVx1_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
INVx2_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_145), .A2(n_220), .B(n_229), .Y(n_219) );
OA21x2_ASAP7_75t_L g432 ( .A1(n_145), .A2(n_433), .B(n_442), .Y(n_432) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_145), .A2(n_447), .B(n_454), .Y(n_446) );
OR2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_163), .Y(n_146) );
AND2x2_ASAP7_75t_L g187 ( .A(n_147), .B(n_163), .Y(n_187) );
BUFx2_ASAP7_75t_L g261 ( .A(n_147), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_147), .A2(n_294), .B1(n_296), .B2(n_297), .Y(n_293) );
OR2x2_ASAP7_75t_L g315 ( .A(n_147), .B(n_175), .Y(n_315) );
AND2x2_ASAP7_75t_L g379 ( .A(n_147), .B(n_257), .Y(n_379) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g247 ( .A(n_148), .B(n_175), .Y(n_247) );
AND2x2_ASAP7_75t_L g254 ( .A(n_148), .B(n_163), .Y(n_254) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_148), .Y(n_296) );
OR2x2_ASAP7_75t_L g331 ( .A(n_148), .B(n_174), .Y(n_331) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_161), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_149), .B(n_162), .Y(n_161) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_149), .A2(n_176), .B(n_184), .Y(n_175) );
INVx2_ASAP7_75t_L g200 ( .A(n_149), .Y(n_200) );
INVx2_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_156), .B1(n_157), .B2(n_158), .Y(n_154) );
INVx2_ASAP7_75t_L g157 ( .A(n_155), .Y(n_157) );
INVx4_ASAP7_75t_L g225 ( .A(n_155), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_160), .A2(n_177), .B(n_178), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_160), .A2(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g250 ( .A(n_163), .Y(n_250) );
INVx3_ASAP7_75t_L g259 ( .A(n_163), .Y(n_259) );
BUFx2_ASAP7_75t_L g283 ( .A(n_163), .Y(n_283) );
AND2x2_ASAP7_75t_L g316 ( .A(n_163), .B(n_251), .Y(n_316) );
INVx1_ASAP7_75t_L g437 ( .A(n_168), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_172), .A2(n_402), .B1(n_403), .B2(n_404), .Y(n_401) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_187), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_174), .B(n_259), .Y(n_263) );
INVx1_ASAP7_75t_L g291 ( .A(n_174), .Y(n_291) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_183), .Y(n_179) );
INVx2_ASAP7_75t_L g459 ( .A(n_181), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_181), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_181), .A2(n_508), .B(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_183), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_186), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_186), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g269 ( .A(n_187), .Y(n_269) );
NAND2x1_ASAP7_75t_SL g188 ( .A(n_189), .B(n_203), .Y(n_188) );
AND2x2_ASAP7_75t_L g267 ( .A(n_189), .B(n_218), .Y(n_267) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_189), .Y(n_341) );
AND2x2_ASAP7_75t_L g368 ( .A(n_189), .B(n_288), .Y(n_368) );
AND2x2_ASAP7_75t_L g376 ( .A(n_189), .B(n_338), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_189), .B(n_233), .Y(n_403) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g234 ( .A(n_190), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g252 ( .A(n_190), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g273 ( .A(n_190), .Y(n_273) );
INVx1_ASAP7_75t_L g279 ( .A(n_190), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_190), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g312 ( .A(n_190), .B(n_236), .Y(n_312) );
OR2x2_ASAP7_75t_L g350 ( .A(n_190), .B(n_305), .Y(n_350) );
AOI32xp33_ASAP7_75t_L g362 ( .A1(n_190), .A2(n_363), .A3(n_366), .B1(n_367), .B2(n_368), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_190), .B(n_338), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_190), .B(n_298), .Y(n_413) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_201), .Y(n_190) );
AOI21xp5_ASAP7_75t_SL g191 ( .A1(n_192), .A2(n_193), .B(n_200), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_197), .A2(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g228 ( .A(n_199), .Y(n_228) );
INVx1_ASAP7_75t_L g243 ( .A(n_200), .Y(n_243) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_200), .A2(n_492), .B(n_501), .Y(n_491) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_200), .A2(n_506), .B(n_513), .Y(n_505) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g324 ( .A(n_204), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_218), .Y(n_204) );
INVx1_ASAP7_75t_L g286 ( .A(n_205), .Y(n_286) );
AND2x2_ASAP7_75t_L g288 ( .A(n_205), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_205), .B(n_235), .Y(n_305) );
AND2x2_ASAP7_75t_L g338 ( .A(n_205), .B(n_314), .Y(n_338) );
AND2x2_ASAP7_75t_L g375 ( .A(n_205), .B(n_236), .Y(n_375) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g233 ( .A(n_206), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_206), .B(n_235), .Y(n_265) );
AND2x2_ASAP7_75t_L g272 ( .A(n_206), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g313 ( .A(n_206), .B(n_314), .Y(n_313) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_216), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_215), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_214), .Y(n_210) );
INVx2_ASAP7_75t_L g289 ( .A(n_218), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_218), .B(n_235), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_218), .B(n_280), .Y(n_361) );
INVx1_ASAP7_75t_L g383 ( .A(n_218), .Y(n_383) );
INVx1_ASAP7_75t_L g400 ( .A(n_218), .Y(n_400) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g253 ( .A(n_219), .B(n_235), .Y(n_253) );
AND2x2_ASAP7_75t_L g275 ( .A(n_219), .B(n_236), .Y(n_275) );
INVx1_ASAP7_75t_L g314 ( .A(n_219), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_225), .B(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_225), .A2(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g496 ( .A(n_225), .Y(n_496) );
AOI221x1_ASAP7_75t_SL g230 ( .A1(n_231), .A2(n_246), .B1(n_252), .B2(n_254), .C(n_255), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_231), .A2(n_319), .B1(n_386), .B2(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
AND2x2_ASAP7_75t_L g277 ( .A(n_232), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g372 ( .A(n_232), .B(n_252), .Y(n_372) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g328 ( .A(n_233), .B(n_253), .Y(n_328) );
INVx1_ASAP7_75t_L g340 ( .A(n_234), .Y(n_340) );
AND2x2_ASAP7_75t_L g351 ( .A(n_234), .B(n_338), .Y(n_351) );
AND2x2_ASAP7_75t_L g418 ( .A(n_234), .B(n_313), .Y(n_418) );
INVx2_ASAP7_75t_L g280 ( .A(n_235), .Y(n_280) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_243), .B(n_244), .Y(n_236) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_247), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g370 ( .A(n_247), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_248), .B(n_331), .Y(n_334) );
INVx3_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_249), .A2(n_370), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NOR2xp33_ASAP7_75t_SL g392 ( .A(n_252), .B(n_278), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_253), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g344 ( .A(n_253), .B(n_272), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_253), .B(n_279), .Y(n_421) );
AND2x2_ASAP7_75t_L g290 ( .A(n_254), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g357 ( .A(n_254), .Y(n_357) );
AOI21xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_260), .B(n_264), .Y(n_255) );
NAND2x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_257), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g306 ( .A(n_257), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g318 ( .A(n_257), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_257), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g342 ( .A(n_258), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_258), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_258), .B(n_261), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_261), .A2(n_300), .B(n_330), .C(n_332), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_261), .A2(n_348), .B1(n_351), .B2(n_352), .C(n_356), .Y(n_347) );
AND2x2_ASAP7_75t_L g343 ( .A(n_262), .B(n_296), .Y(n_343) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g303 ( .A(n_267), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g374 ( .A(n_267), .B(n_375), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_276), .C(n_301), .Y(n_268) );
NAND3xp33_ASAP7_75t_SL g387 ( .A(n_269), .B(n_388), .C(n_389), .Y(n_387) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
OR2x2_ASAP7_75t_L g360 ( .A(n_271), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B1(n_284), .B2(n_290), .C(n_292), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_278), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_278), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g300 ( .A(n_283), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_283), .A2(n_340), .B1(n_341), .B2(n_342), .Y(n_339) );
OR2x2_ASAP7_75t_L g420 ( .A(n_283), .B(n_331), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVxp67_ASAP7_75t_L g394 ( .A(n_286), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_288), .B(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g295 ( .A(n_289), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_291), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_291), .B(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_291), .B(n_358), .Y(n_397) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g411 ( .A(n_300), .B(n_331), .Y(n_411) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g389 ( .A(n_306), .Y(n_389) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI322xp33_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_315), .A3(n_316), .B1(n_317), .B2(n_320), .C1(n_322), .C2(n_324), .Y(n_309) );
OAI322xp33_ASAP7_75t_L g391 ( .A1(n_310), .A2(n_392), .A3(n_393), .B1(n_394), .B2(n_395), .C1(n_396), .C2(n_398), .Y(n_391) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx4_ASAP7_75t_L g325 ( .A(n_312), .Y(n_325) );
AND2x2_ASAP7_75t_L g386 ( .A(n_312), .B(n_338), .Y(n_386) );
AND2x2_ASAP7_75t_L g399 ( .A(n_312), .B(n_400), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_315), .Y(n_410) );
INVx1_ASAP7_75t_L g388 ( .A(n_316), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OR2x2_ASAP7_75t_L g322 ( .A(n_318), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g405 ( .A(n_318), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_318), .B(n_359), .Y(n_416) );
OR2x2_ASAP7_75t_L g349 ( .A(n_321), .B(n_350), .Y(n_349) );
INVxp33_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g326 ( .A1(n_325), .A2(n_327), .B1(n_329), .B2(n_333), .C(n_335), .Y(n_326) );
NOR2xp67_ASAP7_75t_L g382 ( .A(n_325), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g409 ( .A(n_325), .Y(n_409) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
AOI322xp5_ASAP7_75t_L g373 ( .A1(n_332), .A2(n_357), .A3(n_374), .B1(n_376), .B2(n_377), .C1(n_380), .C2(n_384), .Y(n_373) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_339), .B1(n_343), .B2(n_344), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_369), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_362), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_350), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_353), .B(n_364), .Y(n_367) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OAI322xp33_ASAP7_75t_L g407 ( .A1(n_355), .A2(n_408), .A3(n_410), .B1(n_411), .B2(n_412), .C1(n_414), .C2(n_417), .Y(n_407) );
AOI21xp33_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_358), .B(n_360), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_365), .B(n_413), .Y(n_422) );
OAI211xp5_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B(n_373), .C(n_385), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR4xp25_ASAP7_75t_L g390 ( .A(n_391), .B(n_401), .C(n_407), .D(n_419), .Y(n_390) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
CKINVDCx14_ASAP7_75t_R g417 ( .A(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B(n_422), .Y(n_419) );
INVx6_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g713 ( .A(n_424), .Y(n_713) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_425), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g714 ( .A(n_426), .Y(n_714) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_630), .Y(n_426) );
NAND5xp2_ASAP7_75t_L g427 ( .A(n_428), .B(n_549), .C(n_564), .D(n_590), .E(n_612), .Y(n_427) );
NOR2xp33_ASAP7_75t_SL g428 ( .A(n_429), .B(n_529), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_470), .B1(n_502), .B2(n_518), .C(n_519), .Y(n_429) );
NOR2xp33_ASAP7_75t_SL g430 ( .A(n_431), .B(n_462), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_431), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g706 ( .A(n_431), .Y(n_706) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_443), .Y(n_431) );
INVx1_ASAP7_75t_L g546 ( .A(n_432), .Y(n_546) );
AND2x2_ASAP7_75t_L g548 ( .A(n_432), .B(n_456), .Y(n_548) );
AND2x2_ASAP7_75t_L g558 ( .A(n_432), .B(n_455), .Y(n_558) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_432), .Y(n_576) );
INVx1_ASAP7_75t_L g586 ( .A(n_432), .Y(n_586) );
OR2x2_ASAP7_75t_L g624 ( .A(n_432), .B(n_523), .Y(n_624) );
INVx2_ASAP7_75t_L g674 ( .A(n_432), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_432), .B(n_522), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B(n_437), .Y(n_434) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_444), .B(n_455), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_445), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_445), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_SL g606 ( .A(n_445), .B(n_546), .Y(n_606) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_446), .Y(n_464) );
INVx2_ASAP7_75t_L g523 ( .A(n_446), .Y(n_523) );
OR2x2_ASAP7_75t_L g585 ( .A(n_446), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g524 ( .A(n_455), .B(n_466), .Y(n_524) );
AND2x2_ASAP7_75t_L g541 ( .A(n_455), .B(n_521), .Y(n_541) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g465 ( .A(n_456), .B(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g544 ( .A(n_456), .Y(n_544) );
AND2x2_ASAP7_75t_L g673 ( .A(n_456), .B(n_674), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_459), .A2(n_487), .B(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_459), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_461), .A2(n_507), .B(n_510), .Y(n_506) );
INVx1_ASAP7_75t_L g518 ( .A(n_462), .Y(n_518) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
AND2x2_ASAP7_75t_L g636 ( .A(n_463), .B(n_524), .Y(n_636) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g637 ( .A(n_464), .B(n_548), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_465), .A2(n_605), .B(n_607), .C(n_609), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_465), .B(n_605), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_465), .A2(n_535), .B1(n_678), .B2(n_679), .C(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g521 ( .A(n_466), .Y(n_521) );
INVx1_ASAP7_75t_L g557 ( .A(n_466), .Y(n_557) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_466), .Y(n_566) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_480), .Y(n_471) );
AND2x2_ASAP7_75t_L g583 ( .A(n_472), .B(n_528), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_472), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_473), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g675 ( .A(n_473), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g707 ( .A(n_473), .Y(n_707) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g537 ( .A(n_474), .Y(n_537) );
AND2x2_ASAP7_75t_L g563 ( .A(n_474), .B(n_517), .Y(n_563) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_474), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_474), .B(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_480), .B(n_619), .Y(n_654) );
INVx1_ASAP7_75t_SL g658 ( .A(n_480), .Y(n_658) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
INVx3_ASAP7_75t_L g517 ( .A(n_481), .Y(n_517) );
AND2x2_ASAP7_75t_L g528 ( .A(n_481), .B(n_505), .Y(n_528) );
AND2x2_ASAP7_75t_L g550 ( .A(n_481), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g595 ( .A(n_481), .B(n_589), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_481), .B(n_527), .Y(n_676) );
INVx2_ASAP7_75t_L g498 ( .A(n_489), .Y(n_498) );
AND2x2_ASAP7_75t_L g516 ( .A(n_491), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g527 ( .A(n_491), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_491), .B(n_505), .Y(n_552) );
AND2x2_ASAP7_75t_L g588 ( .A(n_491), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_516), .Y(n_503) );
INVx1_ASAP7_75t_L g568 ( .A(n_504), .Y(n_568) );
AND2x2_ASAP7_75t_L g610 ( .A(n_504), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_504), .B(n_531), .Y(n_616) );
AOI21xp5_ASAP7_75t_SL g690 ( .A1(n_504), .A2(n_522), .B(n_545), .Y(n_690) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
OR2x2_ASAP7_75t_L g533 ( .A(n_505), .B(n_514), .Y(n_533) );
AND2x2_ASAP7_75t_L g580 ( .A(n_505), .B(n_517), .Y(n_580) );
INVx2_ASAP7_75t_L g589 ( .A(n_505), .Y(n_589) );
INVx1_ASAP7_75t_L g695 ( .A(n_505), .Y(n_695) );
AND2x2_ASAP7_75t_L g619 ( .A(n_514), .B(n_589), .Y(n_619) );
INVx1_ASAP7_75t_L g644 ( .A(n_514), .Y(n_644) );
AND2x2_ASAP7_75t_L g553 ( .A(n_516), .B(n_537), .Y(n_553) );
AND2x2_ASAP7_75t_L g565 ( .A(n_516), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g683 ( .A(n_516), .Y(n_683) );
INVx2_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g611 ( .A(n_517), .B(n_527), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_517), .B(n_695), .Y(n_694) );
OAI21xp33_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_524), .B(n_525), .Y(n_519) );
AND2x2_ASAP7_75t_L g626 ( .A(n_520), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g680 ( .A(n_520), .Y(n_680) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
BUFx2_ASAP7_75t_L g699 ( .A(n_521), .Y(n_699) );
BUFx2_ASAP7_75t_L g570 ( .A(n_522), .Y(n_570) );
AND2x2_ASAP7_75t_L g672 ( .A(n_522), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g655 ( .A(n_523), .Y(n_655) );
AND2x4_ASAP7_75t_L g582 ( .A(n_524), .B(n_545), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_524), .B(n_606), .Y(n_618) );
AOI32xp33_ASAP7_75t_L g542 ( .A1(n_525), .A2(n_543), .A3(n_545), .B1(n_547), .B2(n_548), .Y(n_542) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
INVx3_ASAP7_75t_L g531 ( .A(n_526), .Y(n_531) );
OR2x2_ASAP7_75t_L g667 ( .A(n_526), .B(n_623), .Y(n_667) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g536 ( .A(n_527), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g643 ( .A(n_527), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g535 ( .A(n_528), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g547 ( .A(n_528), .B(n_537), .Y(n_547) );
INVx1_ASAP7_75t_L g668 ( .A(n_528), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_528), .B(n_643), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_534), .B(n_538), .C(n_542), .Y(n_529) );
OAI322xp33_ASAP7_75t_L g638 ( .A1(n_530), .A2(n_575), .A3(n_639), .B1(n_641), .B2(n_645), .C1(n_646), .C2(n_650), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVxp67_ASAP7_75t_L g603 ( .A(n_531), .Y(n_603) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g657 ( .A(n_533), .B(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_533), .B(n_573), .Y(n_704) );
INVxp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g596 ( .A(n_536), .Y(n_596) );
OR2x2_ASAP7_75t_L g682 ( .A(n_537), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_540), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g591 ( .A(n_541), .B(n_570), .Y(n_591) );
AND2x2_ASAP7_75t_L g662 ( .A(n_541), .B(n_575), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_541), .B(n_649), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_543), .A2(n_550), .B1(n_553), .B2(n_554), .C(n_559), .Y(n_549) );
OR2x2_ASAP7_75t_L g560 ( .A(n_543), .B(n_556), .Y(n_560) );
AND2x2_ASAP7_75t_L g648 ( .A(n_543), .B(n_649), .Y(n_648) );
AOI32xp33_ASAP7_75t_L g687 ( .A1(n_543), .A2(n_573), .A3(n_688), .B1(n_689), .B2(n_692), .Y(n_687) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_544), .B(n_580), .C(n_603), .Y(n_621) );
AND2x2_ASAP7_75t_L g647 ( .A(n_544), .B(n_640), .Y(n_647) );
INVxp67_ASAP7_75t_L g627 ( .A(n_545), .Y(n_627) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_548), .B(n_600), .Y(n_656) );
INVx2_ASAP7_75t_L g666 ( .A(n_548), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_548), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g635 ( .A(n_551), .Y(n_635) );
OR2x2_ASAP7_75t_L g561 ( .A(n_552), .B(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_554), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_557), .Y(n_640) );
AND2x2_ASAP7_75t_L g599 ( .A(n_558), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g645 ( .A(n_558), .Y(n_645) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_558), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_560), .A2(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g678 ( .A(n_563), .B(n_588), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B(n_577), .C(n_584), .Y(n_564) );
AND2x2_ASAP7_75t_L g608 ( .A(n_566), .B(n_576), .Y(n_608) );
INVx2_ASAP7_75t_L g623 ( .A(n_566), .Y(n_623) );
OR2x2_ASAP7_75t_L g661 ( .A(n_566), .B(n_624), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_566), .B(n_704), .Y(n_703) );
AOI211xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_569), .B(n_571), .C(n_574), .Y(n_567) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_570), .B(n_608), .Y(n_607) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_571), .A2(n_666), .B(n_690), .C(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g587 ( .A(n_572), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g629 ( .A(n_573), .B(n_619), .Y(n_629) );
INVx1_ASAP7_75t_L g634 ( .A(n_573), .Y(n_634) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_578), .B(n_581), .Y(n_577) );
INVxp33_ASAP7_75t_L g685 ( .A(n_579), .Y(n_685) );
AND2x2_ASAP7_75t_L g664 ( .A(n_580), .B(n_643), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_585), .A2(n_647), .B(n_648), .Y(n_646) );
OAI322xp33_ASAP7_75t_L g665 ( .A1(n_587), .A2(n_666), .A3(n_667), .B1(n_668), .B2(n_669), .C1(n_671), .C2(n_675), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_597), .B2(n_601), .C(n_604), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g642 ( .A(n_595), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g686 ( .A(n_599), .Y(n_686) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_602), .B(n_622), .Y(n_688) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g651 ( .A(n_611), .B(n_619), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B1(n_617), .B2(n_619), .C(n_620), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_615), .A2(n_632), .B1(n_636), .B2(n_637), .C(n_638), .Y(n_631) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVxp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_619), .B(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_625), .B2(n_628), .Y(n_620) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx2_ASAP7_75t_SL g649 ( .A(n_624), .Y(n_649) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND5xp2_ASAP7_75t_L g630 ( .A(n_631), .B(n_652), .C(n_677), .D(n_687), .E(n_697), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_633), .B(n_635), .Y(n_632) );
NOR4xp25_ASAP7_75t_L g705 ( .A(n_634), .B(n_640), .C(n_706), .D(n_707), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_637), .A2(n_698), .B1(n_700), .B2(n_702), .C(n_705), .Y(n_697) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g696 ( .A(n_643), .Y(n_696) );
OAI322xp33_ASAP7_75t_L g653 ( .A1(n_647), .A2(n_654), .A3(n_655), .B1(n_656), .B2(n_657), .C1(n_659), .C2(n_663), .Y(n_653) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_665), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g698 ( .A(n_673), .B(n_699), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_681) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx2_ASAP7_75t_L g735 ( .A(n_712), .Y(n_735) );
INVx3_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_726), .Y(n_721) );
NOR2xp33_ASAP7_75t_SL g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_SL g747 ( .A(n_723), .Y(n_747) );
INVx1_ASAP7_75t_L g746 ( .A(n_725), .Y(n_746) );
OA21x2_ASAP7_75t_L g749 ( .A1(n_725), .A2(n_740), .B(n_747), .Y(n_749) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_728), .Y(n_738) );
BUFx2_ASAP7_75t_L g740 ( .A(n_728), .Y(n_740) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_736), .B(n_739), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g739 ( .A(n_740), .B(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
endmodule