module fake_jpeg_24036_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_24),
.B1(n_19),
.B2(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_58),
.B1(n_64),
.B2(n_66),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_29),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_34),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_26),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_35),
.B1(n_30),
.B2(n_33),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_21),
.B1(n_27),
.B2(n_33),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_34),
.B1(n_23),
.B2(n_31),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_0),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_72),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_81),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_35),
.B1(n_44),
.B2(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_87),
.B1(n_95),
.B2(n_0),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_80),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_37),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_94),
.B(n_100),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_61),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_91),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_45),
.B1(n_22),
.B2(n_17),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_96),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_101),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_45),
.B(n_22),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_17),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_50),
.B(n_65),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_84),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_50),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_109),
.C(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_111),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_50),
.B(n_65),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_116),
.Y(n_152)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_46),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_123),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_88),
.B1(n_69),
.B2(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_46),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_104),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_134),
.B(n_141),
.C(n_154),
.D(n_118),
.Y(n_169)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_137),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_127),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_142),
.B(n_112),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_144),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_70),
.Y(n_141)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_86),
.C(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_147),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_86),
.B1(n_87),
.B2(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_77),
.B1(n_78),
.B2(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_76),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_147),
.Y(n_191)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_160),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_134),
.C(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_177),
.Y(n_194)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_154),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_107),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_103),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_187),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_71),
.B(n_122),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_141),
.C(n_146),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_195),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_139),
.B1(n_148),
.B2(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

AOI22x1_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_137),
.B1(n_133),
.B2(n_113),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_188),
.B1(n_197),
.B2(n_78),
.Y(n_210)
);

OAI322xp33_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_167),
.A3(n_169),
.B1(n_168),
.B2(n_156),
.C1(n_165),
.C2(n_173),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_113),
.B1(n_153),
.B2(n_90),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_103),
.C(n_111),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_163),
.C(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_125),
.B1(n_108),
.B2(n_81),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_108),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_216)
);

AOI221xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_174),
.B1(n_162),
.B2(n_160),
.C(n_155),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_209),
.C(n_188),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_171),
.C(n_166),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_125),
.C(n_172),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_188),
.B1(n_194),
.B2(n_193),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_85),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_189),
.B(n_116),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_201),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_223),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_217),
.B1(n_197),
.B2(n_212),
.Y(n_230)
);

XOR2x2_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_188),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_221),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_205),
.B(n_198),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_184),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_208),
.A2(n_179),
.B(n_180),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_225),
.B(n_219),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_203),
.C(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_211),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.Y(n_241)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_15),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_232),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_16),
.A3(n_15),
.B1(n_14),
.B2(n_12),
.C1(n_10),
.C2(n_90),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_242),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_227),
.B1(n_232),
.B2(n_226),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_246),
.B(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_228),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_240),
.C(n_3),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_251),
.B(n_243),
.Y(n_253)
);

AOI31xp33_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_3),
.A3(n_6),
.B(n_7),
.Y(n_251)
);

AOI321xp33_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_8),
.A3(n_9),
.B1(n_243),
.B2(n_246),
.C(n_183),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);


endmodule