module fake_jpeg_24080_n_301 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_20),
.B1(n_25),
.B2(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_53),
.B1(n_61),
.B2(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_30),
.B1(n_35),
.B2(n_20),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_58),
.C(n_15),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_56),
.Y(n_65)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_20),
.B1(n_25),
.B2(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_14),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_14),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_18),
.B1(n_17),
.B2(n_29),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_75),
.B1(n_28),
.B2(n_24),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_67),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_33),
.B1(n_38),
.B2(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_17),
.B1(n_29),
.B2(n_21),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_34),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_44),
.C(n_34),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_29),
.B1(n_28),
.B2(n_21),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_29),
.B1(n_28),
.B2(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_81),
.B(n_82),
.Y(n_88)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_51),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_105),
.C(n_44),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_95),
.B1(n_97),
.B2(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_101),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_58),
.B(n_56),
.C(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_84),
.Y(n_112)
);

XNOR2x1_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_48),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_108),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_54),
.B1(n_41),
.B2(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_54),
.B1(n_46),
.B2(n_60),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_15),
.B1(n_16),
.B2(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_47),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_60),
.B1(n_55),
.B2(n_32),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_15),
.B(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_25),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_11),
.B(n_9),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_7),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_16),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_116),
.B1(n_89),
.B2(n_87),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_89),
.B(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_101),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_79),
.B1(n_80),
.B2(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_124),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_99),
.C(n_86),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_81),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_152)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_131),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_93),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_135),
.C(n_138),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_88),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_38),
.B(n_33),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_109),
.B1(n_116),
.B2(n_117),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_147),
.C(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_86),
.B1(n_87),
.B2(n_69),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_112),
.B1(n_115),
.B2(n_119),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_69),
.C(n_100),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_131),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_69),
.B1(n_68),
.B2(n_100),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_155),
.B1(n_113),
.B2(n_114),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_32),
.B1(n_92),
.B2(n_70),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_70),
.B1(n_24),
.B2(n_15),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_158),
.B1(n_67),
.B2(n_125),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_24),
.B1(n_16),
.B2(n_27),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_169),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_164),
.B1(n_156),
.B2(n_136),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_147),
.B1(n_141),
.B2(n_140),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_174),
.B1(n_135),
.B2(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_120),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_118),
.B1(n_121),
.B2(n_27),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_175),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_27),
.B(n_19),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_177),
.B(n_179),
.Y(n_198)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_19),
.B(n_1),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_148),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_19),
.B(n_2),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_191),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_138),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_168),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_205),
.B1(n_174),
.B2(n_169),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_38),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_164),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_83),
.B1(n_33),
.B2(n_3),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_83),
.C(n_2),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_201),
.C(n_182),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_83),
.C(n_3),
.Y(n_201)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_171),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_167),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_183),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_206),
.B(n_197),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_175),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_189),
.B(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_219),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_190),
.CI(n_206),
.CON(n_228),
.SN(n_228)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_162),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_172),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_179),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_177),
.C(n_161),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_200),
.C(n_205),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_198),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_176),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_198),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_8),
.B(n_11),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_224),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_202),
.B1(n_188),
.B2(n_195),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_207),
.B1(n_225),
.B2(n_219),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_235),
.C(n_244),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_192),
.C(n_200),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_0),
.Y(n_254)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_193),
.C(n_4),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_229),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_246),
.B1(n_228),
.B2(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_209),
.C(n_222),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_258),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_4),
.C(n_5),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_256),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_5),
.C(n_6),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_7),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_6),
.CI(n_7),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_6),
.C(n_9),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_231),
.B(n_239),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_270),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_262),
.A2(n_248),
.B1(n_254),
.B2(n_241),
.Y(n_280)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_264),
.B(n_268),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_234),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_228),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_242),
.B(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_240),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_256),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_227),
.Y(n_275)
);

AOI31xp33_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_278),
.A3(n_265),
.B(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_251),
.B(n_248),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_282),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_10),
.B1(n_12),
.B2(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_9),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_10),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_286),
.B(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_285),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_266),
.C(n_10),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_274),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_292),
.C(n_294),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_293),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_291),
.C(n_278),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_298),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_296),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_12),
.C(n_295),
.Y(n_301)
);


endmodule