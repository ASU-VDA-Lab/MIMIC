module fake_jpeg_17338_n_185 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

OR2x2_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_27),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_18),
.B1(n_22),
.B2(n_28),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_45),
.B1(n_48),
.B2(n_55),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_25),
.C(n_30),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_18),
.B1(n_22),
.B2(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_18),
.B1(n_16),
.B2(n_20),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_25),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_25),
.B(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_23),
.B1(n_20),
.B2(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_32),
.A2(n_23),
.B1(n_29),
.B2(n_19),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_21),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_73),
.B1(n_54),
.B2(n_21),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_75),
.Y(n_80)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_15),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_39),
.B1(n_31),
.B2(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_54),
.B1(n_47),
.B2(n_33),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_40),
.B1(n_27),
.B2(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_38),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_49),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_57),
.C(n_43),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_83),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_38),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_62),
.B(n_66),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_69),
.B1(n_59),
.B2(n_65),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_64),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_92),
.B1(n_97),
.B2(n_70),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_95),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_33),
.B1(n_38),
.B2(n_43),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_38),
.B1(n_43),
.B2(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_107),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_61),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_108),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_92),
.B(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_114),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_67),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_103),
.A3(n_98),
.B1(n_115),
.B2(n_94),
.C1(n_107),
.C2(n_99),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_65),
.Y(n_128)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_113),
.B1(n_108),
.B2(n_74),
.C(n_104),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_91),
.C(n_95),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_126),
.C(n_42),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_84),
.B1(n_85),
.B2(n_76),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_123),
.B(n_124),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_68),
.B1(n_78),
.B2(n_90),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_96),
.B(n_86),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_127),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_73),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_97),
.B(n_71),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_30),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_42),
.B(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_129),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_135),
.Y(n_152)
);

OAI321xp33_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_139),
.A3(n_127),
.B1(n_122),
.B2(n_129),
.C(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_26),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_140),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_144),
.C(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_145),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_51),
.B1(n_1),
.B2(n_2),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_119),
.B1(n_130),
.B2(n_3),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_57),
.C(n_87),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_14),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_137),
.B(n_131),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_148),
.C(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_144),
.C(n_126),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_125),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.C(n_156),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_139),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_164),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_51),
.C(n_57),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_0),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_153),
.B(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_170),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_2),
.B(n_3),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_7),
.C(n_9),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_4),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.C(n_8),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_176),
.B(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_7),
.Y(n_177)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_167),
.B(n_170),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_9),
.B(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_172),
.B(n_10),
.C(n_11),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.C(n_11),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_9),
.C(n_10),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);


endmodule