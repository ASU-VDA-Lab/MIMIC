module fake_aes_3921_n_20 (n_3, n_1, n_2, n_0, n_20);
input n_3;
input n_1;
input n_2;
input n_0;
output n_20;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_4;
wire n_7;
INVx1_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
INVx1_ASAP7_75t_SL g6 ( .A(n_2), .Y(n_6) );
BUFx6f_ASAP7_75t_SL g7 ( .A(n_3), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_4), .B(n_0), .Y(n_8) );
O2A1O1Ixp33_ASAP7_75t_SL g9 ( .A1(n_4), .A2(n_0), .B(n_1), .C(n_2), .Y(n_9) );
AO31x2_ASAP7_75t_L g10 ( .A1(n_5), .A2(n_0), .A3(n_1), .B(n_2), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
NOR3xp33_ASAP7_75t_L g13 ( .A(n_11), .B(n_6), .C(n_9), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_12), .B(n_11), .Y(n_14) );
AOI322xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_12), .A3(n_5), .B1(n_3), .B2(n_1), .C1(n_0), .C2(n_7), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_13), .A2(n_7), .B1(n_10), .B2(n_3), .Y(n_16) );
NAND4xp75_ASAP7_75t_L g17 ( .A(n_15), .B(n_7), .C(n_10), .D(n_3), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_16), .B(n_10), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_10), .B1(n_17), .B2(n_12), .Y(n_19) );
OR2x6_ASAP7_75t_L g20 ( .A(n_19), .B(n_10), .Y(n_20) );
endmodule