module fake_ariane_335_n_1969 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1969);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1969;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_137),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_87),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_38),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_144),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_128),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_85),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_98),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_57),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_136),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_18),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_175),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_44),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_62),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_56),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_148),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_2),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_30),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_76),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_142),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_59),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_57),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_71),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_72),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_32),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_105),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_80),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_41),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_38),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_96),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_43),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_152),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_65),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_28),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_30),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_65),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_18),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_179),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_120),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_165),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_162),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_127),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_68),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_69),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_6),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_147),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_133),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_43),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_33),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_163),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_103),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_29),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_47),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_44),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_185),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_82),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_19),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_184),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_9),
.Y(n_273)
);

BUFx8_ASAP7_75t_SL g274 ( 
.A(n_77),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_140),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_164),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_56),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_94),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_13),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_34),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_63),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_10),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_70),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_62),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_93),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_22),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_167),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_159),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_45),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_129),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_160),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_97),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_83),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_58),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_10),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_37),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_84),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_155),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_192),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_161),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_5),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_11),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_139),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_61),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_15),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_86),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_124),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_130),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_35),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_40),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_78),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_22),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_17),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_131),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_111),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_141),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_172),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_116),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_154),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_123),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_109),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_110),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_2),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_132),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_81),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_25),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_122),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_20),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_126),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_52),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_42),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_58),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_66),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_54),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_50),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_8),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_75),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_121),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_99),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_3),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_37),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_145),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_5),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_108),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_143),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_74),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_47),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_67),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_119),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_31),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_73),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_40),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_54),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_92),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_45),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_102),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_166),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_34),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_24),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_17),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_23),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_6),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_151),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_26),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_28),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_11),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_112),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_169),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_61),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_12),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_101),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_23),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_41),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_59),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_168),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_117),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_33),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_24),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_48),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_63),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_14),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_88),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_297),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_297),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_196),
.B(n_0),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_224),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_274),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_381),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_297),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_297),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_0),
.Y(n_394)
);

BUFx2_ASAP7_75t_SL g395 ( 
.A(n_198),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_250),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_297),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_198),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_255),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_354),
.B(n_1),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_328),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_342),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_371),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_4),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_238),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_240),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_242),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_234),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_244),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_251),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_254),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_265),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_257),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_259),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_262),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_368),
.B(n_7),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_267),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_271),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_336),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_273),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_376),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_305),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_381),
.B(n_7),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_226),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_376),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_277),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_253),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_253),
.B(n_14),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_226),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_279),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_280),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_281),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_194),
.B(n_15),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_285),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_294),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_296),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_287),
.B(n_343),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_287),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_304),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_312),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_231),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_313),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_343),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_246),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_308),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_246),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_258),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_331),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_197),
.B(n_16),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_315),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_333),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_206),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_198),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_258),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_200),
.B(n_16),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_329),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_199),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_203),
.B(n_19),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_207),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_206),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_226),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_208),
.B(n_20),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_221),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_270),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_270),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_318),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_318),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_209),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_207),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_454),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_386),
.A2(n_216),
.B(n_215),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_365),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_391),
.B(n_301),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_223),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_228),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_459),
.B(n_252),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_454),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_454),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_232),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_399),
.B(n_320),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_395),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_460),
.B(n_233),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_429),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_420),
.B(n_367),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_467),
.B(n_252),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_434),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_467),
.B(n_227),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_239),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_397),
.A2(n_276),
.B(n_261),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_473),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_477),
.B(n_282),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_397),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_478),
.B(n_286),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_446),
.A2(n_330),
.B(n_320),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_478),
.B(n_289),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_479),
.B(n_227),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_398),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_479),
.B(n_299),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_480),
.B(n_470),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_480),
.B(n_207),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_450),
.B(n_260),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_481),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_402),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_402),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_403),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_404),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_405),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_405),
.B(n_300),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_406),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_406),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_416),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_416),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_468),
.B(n_302),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_418),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_413),
.B(n_314),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

CKINVDCx8_ASAP7_75t_R g552 ( 
.A(n_389),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_431),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_433),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_433),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_412),
.B(n_260),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_440),
.B(n_284),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_440),
.B(n_284),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_500),
.B(n_414),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_488),
.B(n_419),
.C(n_415),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_500),
.B(n_399),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_547),
.A2(n_394),
.B1(n_408),
.B2(n_388),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_489),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_489),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_441),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_482),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_531),
.B(n_466),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_488),
.B(n_424),
.C(n_421),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_521),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_531),
.B(n_559),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_521),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_514),
.B(n_466),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_514),
.B(n_425),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

BUFx8_ASAP7_75t_SL g582 ( 
.A(n_517),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_499),
.B(n_427),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_550),
.B(n_472),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_485),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_497),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_485),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_521),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_494),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_509),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_521),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_531),
.B(n_559),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_552),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

INVxp33_ASAP7_75t_L g599 ( 
.A(n_487),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_560),
.B(n_472),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_501),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_518),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_539),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_494),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_494),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_515),
.B(n_248),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_503),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_539),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_550),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_539),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_517),
.A2(n_442),
.B1(n_437),
.B2(n_474),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_482),
.Y(n_612)
);

BUFx10_ASAP7_75t_L g613 ( 
.A(n_515),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_560),
.B(n_428),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_560),
.B(n_430),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_534),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_499),
.B(n_439),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_518),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_503),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_482),
.B(n_443),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_484),
.B(n_516),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_518),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_510),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_497),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_518),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_499),
.B(n_444),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_545),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_506),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_497),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_545),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_547),
.B(n_445),
.Y(n_631)
);

INVx4_ASAP7_75t_SL g632 ( 
.A(n_486),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_499),
.A2(n_475),
.B1(n_471),
.B2(n_462),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_494),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_497),
.B(n_451),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_530),
.B(n_448),
.C(n_447),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_545),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_518),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_494),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_556),
.B(n_449),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_545),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_556),
.B(n_452),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_545),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_510),
.A2(n_426),
.B1(n_423),
.B2(n_435),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_506),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_534),
.B(n_453),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_526),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_510),
.A2(n_298),
.B1(n_229),
.B2(n_225),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_552),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_511),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_556),
.B(n_455),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_508),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_530),
.B(n_461),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_534),
.B(n_390),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_556),
.B(n_464),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_511),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_529),
.Y(n_657)
);

BUFx4f_ASAP7_75t_L g658 ( 
.A(n_484),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_509),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_529),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_508),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_556),
.B(n_330),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_508),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_552),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_533),
.B(n_396),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_508),
.B(n_349),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_532),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_526),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_526),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_533),
.B(n_407),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_508),
.B(n_409),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g672 ( 
.A(n_490),
.B(n_237),
.C(n_235),
.Y(n_672)
);

BUFx4f_ASAP7_75t_L g673 ( 
.A(n_484),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_520),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_532),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_520),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_536),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_520),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_507),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_R g680 ( 
.A(n_484),
.B(n_410),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_536),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_510),
.B(n_317),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_510),
.B(n_525),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_535),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_533),
.A2(n_400),
.B1(n_411),
.B2(n_458),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_509),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_525),
.A2(n_369),
.B1(n_339),
.B2(n_338),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_533),
.B(n_332),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_525),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_535),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_541),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_525),
.B(n_327),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_525),
.B(n_533),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_535),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_541),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_193),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_543),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_490),
.B(n_212),
.C(n_209),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_492),
.A2(n_339),
.B1(n_338),
.B2(n_346),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_543),
.Y(n_700)
);

INVx6_ASAP7_75t_L g701 ( 
.A(n_520),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_492),
.B(n_451),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_544),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_523),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_544),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_528),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_498),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_487),
.B(n_283),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_546),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_538),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_498),
.B(n_340),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_509),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_546),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_647),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_666),
.A2(n_516),
.B1(n_484),
.B2(n_522),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_707),
.B(n_502),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_653),
.B(n_502),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_583),
.B(n_507),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_596),
.B(n_512),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_583),
.B(n_507),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_647),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_588),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_587),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_596),
.B(n_422),
.Y(n_724)
);

OAI221xp5_ASAP7_75t_L g725 ( 
.A1(n_633),
.A2(n_363),
.B1(n_268),
.B2(n_372),
.C(n_266),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_582),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_668),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_631),
.B(n_512),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_576),
.B(n_595),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_565),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_620),
.B(n_519),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_563),
.B(n_519),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_614),
.B(n_522),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_615),
.B(n_524),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_617),
.B(n_523),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_613),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_579),
.B(n_524),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_616),
.B(n_432),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_613),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_616),
.B(n_463),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_585),
.B(n_469),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_668),
.Y(n_742)
);

INVxp33_ASAP7_75t_L g743 ( 
.A(n_708),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_566),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_669),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_569),
.B(n_527),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_669),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_R g748 ( 
.A(n_654),
.B(n_212),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_609),
.B(n_523),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_569),
.B(n_527),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_609),
.B(n_193),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_570),
.B(n_542),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_666),
.A2(n_516),
.B1(n_557),
.B2(n_548),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_612),
.B(n_542),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_564),
.B(n_217),
.C(n_213),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_609),
.B(n_195),
.Y(n_756)
);

INVxp33_ASAP7_75t_L g757 ( 
.A(n_708),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_600),
.B(n_217),
.C(n_213),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_612),
.A2(n_245),
.B1(n_222),
.B2(n_218),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_684),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_568),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_700),
.B(n_195),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_700),
.B(n_201),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_613),
.B(n_487),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_649),
.B(n_307),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_568),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_711),
.B(n_548),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_602),
.A2(n_516),
.B(n_495),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_700),
.B(n_591),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_679),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_679),
.B(n_219),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_702),
.B(n_551),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_684),
.Y(n_773)
);

BUFx5_ASAP7_75t_L g774 ( 
.A(n_662),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_584),
.B(n_626),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_572),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_702),
.B(n_551),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_572),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_702),
.B(n_557),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_567),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_702),
.B(n_558),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_655),
.B(n_558),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_573),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_649),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_591),
.B(n_201),
.Y(n_785)
);

BUFx5_ASAP7_75t_L g786 ( 
.A(n_662),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_591),
.B(n_202),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_640),
.B(n_202),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_642),
.B(n_219),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_567),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_573),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_664),
.B(n_567),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_604),
.B(n_605),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_604),
.A2(n_335),
.B1(n_230),
.B2(n_220),
.Y(n_795)
);

BUFx6f_ASAP7_75t_SL g796 ( 
.A(n_664),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_567),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_690),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_604),
.B(n_204),
.Y(n_799)
);

BUFx6f_ASAP7_75t_SL g800 ( 
.A(n_662),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_605),
.B(n_204),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_605),
.B(n_205),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_606),
.A2(n_688),
.B(n_598),
.C(n_601),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_634),
.B(n_205),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_581),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_634),
.A2(n_346),
.B1(n_355),
.B2(n_230),
.Y(n_806)
);

BUFx4_ASAP7_75t_L g807 ( 
.A(n_599),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_694),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_634),
.B(n_210),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_639),
.A2(n_358),
.B1(n_220),
.B2(n_335),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_651),
.B(n_636),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_581),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_587),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_598),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_694),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_606),
.A2(n_290),
.B(n_243),
.C(n_241),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_639),
.B(n_210),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_611),
.B(n_337),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_662),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_665),
.B(n_307),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_639),
.B(n_211),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_652),
.B(n_661),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_670),
.B(n_307),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_601),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_652),
.B(n_211),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_680),
.B(n_337),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_624),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_666),
.A2(n_516),
.B1(n_554),
.B2(n_553),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_652),
.B(n_214),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_689),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_661),
.B(n_214),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_562),
.B(n_350),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_661),
.B(n_218),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_646),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_571),
.B(n_350),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_663),
.B(n_222),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_607),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_624),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_710),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_607),
.Y(n_840)
);

INVx8_ASAP7_75t_L g841 ( 
.A(n_662),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_619),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_663),
.B(n_348),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_644),
.B(n_344),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_710),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_623),
.A2(n_348),
.B1(n_352),
.B2(n_357),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_635),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_663),
.B(n_635),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_689),
.B(n_326),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_344),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_671),
.Y(n_851)
);

BUFx6f_ASAP7_75t_SL g852 ( 
.A(n_662),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_682),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_698),
.B(n_380),
.C(n_351),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_658),
.B(n_352),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_662),
.B(n_357),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_561),
.B(n_351),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_692),
.B(n_359),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_623),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_580),
.B(n_353),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_693),
.B(n_359),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_623),
.A2(n_360),
.B1(n_379),
.B2(n_347),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_658),
.B(n_360),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_666),
.A2(n_538),
.B1(n_554),
.B2(n_553),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_602),
.B(n_379),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_619),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_602),
.B(n_538),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_687),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_618),
.B(n_540),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_629),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_628),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_618),
.B(n_540),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_588),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_574),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_574),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_577),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_618),
.B(n_540),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_577),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_623),
.Y(n_879)
);

NAND2x1_ASAP7_75t_L g880 ( 
.A(n_701),
.B(n_486),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_683),
.B(n_353),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_658),
.B(n_341),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_628),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_645),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_728),
.B(n_648),
.Y(n_885)
);

OAI321xp33_ASAP7_75t_L g886 ( 
.A1(n_725),
.A2(n_699),
.A3(n_356),
.B1(n_361),
.B2(n_364),
.C(n_334),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_728),
.B(n_666),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_733),
.B(n_666),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_733),
.B(n_734),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_717),
.A2(n_704),
.B(n_625),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_819),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_719),
.B(n_811),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_732),
.B(n_629),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_714),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_734),
.A2(n_666),
.B1(n_701),
.B2(n_672),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_819),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_735),
.A2(n_704),
.B(n_625),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_741),
.B(n_456),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_735),
.A2(n_625),
.B(n_622),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_731),
.B(n_622),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_731),
.B(n_622),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_867),
.A2(n_674),
.B(n_638),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_752),
.B(n_638),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_869),
.A2(n_674),
.B(n_638),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_737),
.B(n_674),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_872),
.A2(n_678),
.B(n_676),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_752),
.B(n_729),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_774),
.B(n_578),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_716),
.B(n_676),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_768),
.A2(n_673),
.B(n_590),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_730),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_738),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_851),
.B(n_676),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_848),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_853),
.B(n_678),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_740),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_714),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_792),
.B(n_632),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_721),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_877),
.A2(n_678),
.B(n_673),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_774),
.B(n_578),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_868),
.A2(n_701),
.B1(n_696),
.B2(n_660),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_775),
.A2(n_608),
.B(n_590),
.C(n_593),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_749),
.A2(n_673),
.B(n_594),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_746),
.B(n_750),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_749),
.A2(n_594),
.B(n_593),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_847),
.B(n_645),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_775),
.A2(n_610),
.B(n_597),
.C(n_627),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_792),
.B(n_632),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_803),
.A2(n_603),
.B(n_597),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_754),
.B(n_650),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_744),
.A2(n_701),
.B1(n_650),
.B2(n_709),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_834),
.B(n_656),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_811),
.A2(n_603),
.B(n_608),
.C(n_610),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_819),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_879),
.B(n_751),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_789),
.B(n_656),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_855),
.A2(n_630),
.B(n_627),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_761),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_789),
.B(n_657),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_774),
.B(n_630),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_841),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_766),
.A2(n_713),
.B1(n_657),
.B2(n_709),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_841),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_718),
.B(n_456),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_721),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_882),
.A2(n_641),
.B(n_637),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_841),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_855),
.A2(n_863),
.B(n_767),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_863),
.A2(n_641),
.B(n_637),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_784),
.B(n_660),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_751),
.B(n_667),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_830),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_756),
.B(n_667),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_794),
.A2(n_643),
.B(n_706),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_820),
.B(n_823),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_SL g957 ( 
.A(n_726),
.B(n_284),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_727),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_882),
.A2(n_643),
.B(n_713),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_774),
.B(n_659),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_776),
.A2(n_675),
.B1(n_677),
.B2(n_705),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_822),
.A2(n_875),
.B(n_874),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_778),
.A2(n_675),
.B1(n_677),
.B2(n_705),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_783),
.A2(n_703),
.B(n_697),
.C(n_695),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_832),
.A2(n_695),
.B(n_703),
.C(n_697),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_791),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_756),
.B(n_681),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_805),
.A2(n_814),
.B1(n_824),
.B2(n_812),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_758),
.B(n_755),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_762),
.B(n_588),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_722),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_832),
.B(n_383),
.C(n_375),
.Y(n_972)
);

O2A1O1Ixp5_ASAP7_75t_L g973 ( 
.A1(n_782),
.A2(n_691),
.B(n_681),
.C(n_706),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_720),
.B(n_621),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_874),
.A2(n_691),
.B(n_621),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_875),
.A2(n_706),
.B(n_589),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_838),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_727),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_876),
.A2(n_586),
.B(n_575),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_837),
.A2(n_575),
.B1(n_586),
.B2(n_589),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_765),
.B(n_344),
.Y(n_981)
);

AO21x2_ASAP7_75t_L g982 ( 
.A1(n_772),
.A2(n_779),
.B(n_777),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_881),
.B(n_575),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_876),
.A2(n_589),
.B(n_586),
.Y(n_984)
);

NOR2x2_ASAP7_75t_L g985 ( 
.A(n_748),
.B(n_355),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_844),
.A2(n_621),
.B1(n_554),
.B2(n_549),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_835),
.B(n_588),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_881),
.B(n_588),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_878),
.A2(n_659),
.B(n_686),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_840),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_842),
.B(n_659),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_878),
.A2(n_659),
.B(n_686),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_866),
.B(n_659),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_871),
.A2(n_884),
.B1(n_883),
.B2(n_859),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_770),
.B(n_358),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_742),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_835),
.A2(n_378),
.B(n_370),
.C(n_366),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_838),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_769),
.A2(n_712),
.B(n_686),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_774),
.B(n_686),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_780),
.B(n_632),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_858),
.B(n_362),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_724),
.B(n_362),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_769),
.A2(n_712),
.B(n_686),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_849),
.B(n_369),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_745),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_771),
.B(n_373),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_807),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_816),
.A2(n_715),
.B(n_781),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_849),
.B(n_373),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_828),
.A2(n_483),
.B(n_495),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_745),
.A2(n_483),
.B(n_495),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_715),
.A2(n_712),
.B(n_686),
.Y(n_1013)
);

OAI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_857),
.A2(n_377),
.B(n_380),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_762),
.B(n_377),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_865),
.A2(n_712),
.B(n_592),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_850),
.B(n_382),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_764),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_763),
.B(n_382),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_763),
.B(n_384),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_857),
.B(n_384),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_860),
.B(n_592),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_787),
.A2(n_804),
.B(n_799),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_860),
.B(n_592),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_747),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_787),
.A2(n_712),
.B(n_592),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_747),
.A2(n_712),
.B(n_592),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_826),
.B(n_549),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_826),
.B(n_549),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_799),
.A2(n_483),
.B(n_496),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_804),
.A2(n_496),
.B(n_236),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_831),
.A2(n_496),
.B(n_247),
.Y(n_1032)
);

INVx8_ASAP7_75t_L g1033 ( 
.A(n_796),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_831),
.A2(n_310),
.B(n_249),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_827),
.B(n_553),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_760),
.A2(n_349),
.B(n_504),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_833),
.A2(n_309),
.B(n_256),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_760),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_773),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_861),
.B(n_504),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_723),
.B(n_504),
.Y(n_1041)
);

OAI22x1_ASAP7_75t_L g1042 ( 
.A1(n_818),
.A2(n_295),
.B1(n_263),
.B2(n_264),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_773),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_793),
.A2(n_505),
.B(n_513),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_793),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_736),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_722),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_723),
.B(n_505),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_739),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_798),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_813),
.B(n_505),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_785),
.A2(n_293),
.B1(n_321),
.B2(n_537),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_743),
.B(n_757),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_813),
.B(n_513),
.Y(n_1054)
);

INVx5_ASAP7_75t_L g1055 ( 
.A(n_722),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_722),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_833),
.A2(n_880),
.B(n_788),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_801),
.A2(n_319),
.B(n_269),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_802),
.A2(n_321),
.B1(n_293),
.B2(n_537),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_809),
.A2(n_322),
.B(n_272),
.Y(n_1060)
);

NOR2x1p5_ASAP7_75t_L g1061 ( 
.A(n_854),
.B(n_275),
.Y(n_1061)
);

OAI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_759),
.A2(n_323),
.B(n_278),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_798),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_817),
.B(n_513),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_774),
.B(n_786),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_808),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_821),
.A2(n_324),
.B(n_288),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_870),
.B(n_509),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_748),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_825),
.A2(n_843),
.B(n_836),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_829),
.B(n_632),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_870),
.B(n_806),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_L g1073 ( 
.A1(n_808),
.A2(n_486),
.B(n_509),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_815),
.A2(n_311),
.B(n_291),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_815),
.A2(n_385),
.B(n_303),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_1033),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_889),
.B(n_796),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_1033),
.B(n_1008),
.Y(n_1078)
);

NAND3xp33_ASAP7_75t_SL g1079 ( 
.A(n_972),
.B(n_862),
.C(n_846),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_1003),
.B(n_800),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_918),
.B(n_790),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_894),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_907),
.B(n_797),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_912),
.B(n_795),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_911),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_918),
.B(n_873),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_956),
.B(n_810),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_916),
.B(n_839),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_900),
.A2(n_901),
.B(n_903),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_952),
.A2(n_954),
.B(n_967),
.C(n_972),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_929),
.B(n_873),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_942),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_905),
.A2(n_856),
.B(n_873),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_925),
.B(n_839),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1033),
.Y(n_1095)
);

OA22x2_ASAP7_75t_L g1096 ( 
.A1(n_974),
.A2(n_845),
.B1(n_753),
.B2(n_828),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_981),
.B(n_845),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_929),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1019),
.A2(n_852),
.B1(n_800),
.B2(n_786),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_917),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_905),
.A2(n_873),
.B(n_753),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_974),
.B(n_852),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_919),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_971),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1021),
.A2(n_864),
.B(n_25),
.C(n_26),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_890),
.A2(n_864),
.B(n_786),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_893),
.A2(n_786),
.B(n_292),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_885),
.A2(n_786),
.B1(n_555),
.B2(n_537),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1017),
.B(n_786),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_893),
.A2(n_909),
.B(n_887),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_937),
.A2(n_306),
.B(n_374),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_940),
.A2(n_21),
.B(n_27),
.C(n_29),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_1053),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_SL g1114 ( 
.A(n_942),
.B(n_231),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_952),
.A2(n_21),
.B(n_27),
.C(n_31),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1070),
.A2(n_374),
.B(n_231),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1019),
.A2(n_997),
.B(n_1014),
.C(n_969),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_933),
.B(n_32),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_892),
.B(n_35),
.Y(n_1119)
);

OAI22x1_ASAP7_75t_L g1120 ( 
.A1(n_936),
.A2(n_36),
.B1(n_39),
.B2(n_46),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_933),
.B(n_36),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_974),
.B(n_39),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1069),
.B(n_555),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_936),
.B(n_46),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_888),
.A2(n_374),
.B(n_231),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_931),
.B(n_555),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_939),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_953),
.Y(n_1128)
);

AND2x6_ASAP7_75t_SL g1129 ( 
.A(n_995),
.B(n_48),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_942),
.Y(n_1130)
);

O2A1O1Ixp5_ASAP7_75t_L g1131 ( 
.A1(n_949),
.A2(n_1023),
.B(n_970),
.C(n_973),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_945),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_898),
.B(n_509),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_910),
.A2(n_555),
.B(n_537),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_946),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_914),
.A2(n_555),
.B1(n_537),
.B2(n_528),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_1018),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_895),
.B(n_555),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_953),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1001),
.B(n_509),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_914),
.B(n_555),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_957),
.B(n_118),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_913),
.B(n_49),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_954),
.B(n_555),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_985),
.Y(n_1145)
);

BUFx8_ASAP7_75t_SL g1146 ( 
.A(n_1007),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_958),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_967),
.B(n_537),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_978),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_913),
.B(n_537),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_915),
.B(n_49),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_SL g1152 ( 
.A(n_1055),
.B(n_528),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_915),
.B(n_50),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1042),
.A2(n_231),
.B1(n_374),
.B2(n_53),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_966),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_977),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1006),
.Y(n_1157)
);

AO32x2_ASAP7_75t_L g1158 ( 
.A1(n_968),
.A2(n_537),
.A3(n_528),
.B1(n_53),
.B2(n_55),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_990),
.A2(n_528),
.B1(n_374),
.B2(n_486),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1002),
.B(n_51),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_942),
.B(n_528),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1005),
.B(n_51),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_971),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_969),
.A2(n_528),
.B(n_248),
.C(n_60),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_982),
.B(n_528),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_982),
.B(n_248),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_1046),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_977),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_932),
.A2(n_897),
.B(n_920),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_971),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_975),
.A2(n_114),
.B(n_158),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_943),
.A2(n_486),
.B1(n_55),
.B2(n_60),
.Y(n_1172)
);

OR2x6_ASAP7_75t_SL g1173 ( 
.A(n_1010),
.B(n_52),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1072),
.A2(n_248),
.B1(n_486),
.B2(n_67),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1015),
.B(n_64),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_927),
.B(n_64),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_1001),
.B(n_66),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_998),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_886),
.B(n_248),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1016),
.A2(n_899),
.B(n_983),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_924),
.A2(n_248),
.B(n_89),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_951),
.B(n_248),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_971),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_987),
.B(n_248),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_987),
.B(n_79),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_961),
.B(n_90),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_996),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_926),
.A2(n_91),
.B(n_95),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1062),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_1049),
.B(n_113),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_994),
.A2(n_134),
.B1(n_135),
.B2(n_146),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_963),
.B(n_149),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1028),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1020),
.B(n_153),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_965),
.A2(n_156),
.B(n_174),
.C(n_178),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_R g1196 ( 
.A(n_998),
.B(n_181),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1025),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1009),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_948),
.B(n_186),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_934),
.A2(n_189),
.B(n_928),
.C(n_923),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1038),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_SL g1202 ( 
.A(n_948),
.B(n_1055),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1043),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1050),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1039),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_962),
.A2(n_906),
.B(n_902),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_964),
.A2(n_980),
.B(n_973),
.C(n_1075),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1061),
.B(n_986),
.Y(n_1208)
);

OAI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_922),
.A2(n_986),
.B1(n_964),
.B2(n_988),
.C(n_959),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1063),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1066),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1045),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_948),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1029),
.B(n_1047),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_948),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1040),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1012),
.A2(n_1073),
.B(n_1064),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_SL g1218 ( 
.A1(n_1022),
.A2(n_1024),
.B(n_993),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1055),
.B(n_1047),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_891),
.B(n_896),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1036),
.B(n_1055),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1047),
.B(n_1056),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_991),
.B(n_1047),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_904),
.A2(n_1027),
.B(n_941),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1056),
.B(n_1035),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1057),
.A2(n_1013),
.B(n_947),
.C(n_979),
.Y(n_1226)
);

INVx6_ASAP7_75t_L g1227 ( 
.A(n_1056),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_891),
.A2(n_896),
.B1(n_944),
.B2(n_935),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1056),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_908),
.A2(n_921),
.B(n_941),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_984),
.A2(n_930),
.B(n_950),
.C(n_938),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1058),
.A2(n_1067),
.B(n_1060),
.C(n_908),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_935),
.B(n_944),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1041),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1034),
.B(n_1037),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1048),
.B(n_1054),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_921),
.A2(n_1071),
.B(n_976),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1051),
.B(n_1074),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1085),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1237),
.A2(n_1011),
.B(n_1030),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1132),
.B(n_1068),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1166),
.A2(n_1059),
.A3(n_1052),
.B(n_989),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1166),
.A2(n_992),
.A3(n_1026),
.B(n_1032),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1090),
.B(n_1068),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1089),
.A2(n_960),
.B(n_1000),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1087),
.A2(n_1079),
.B(n_1160),
.C(n_1117),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1110),
.A2(n_1180),
.B(n_1134),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1098),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1134),
.A2(n_960),
.B(n_1000),
.Y(n_1249)
);

AOI221x1_ASAP7_75t_L g1250 ( 
.A1(n_1120),
.A2(n_1031),
.B1(n_955),
.B2(n_1044),
.C(n_999),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1098),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1099),
.A2(n_1065),
.B(n_1004),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1093),
.A2(n_1206),
.B(n_1101),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1143),
.A2(n_1065),
.B1(n_1121),
.B2(n_1118),
.Y(n_1254)
);

AO32x2_ASAP7_75t_L g1255 ( 
.A1(n_1172),
.A2(n_1108),
.A3(n_1154),
.B1(n_1136),
.B2(n_1159),
.Y(n_1255)
);

NAND2x1_ASAP7_75t_L g1256 ( 
.A(n_1227),
.B(n_1152),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1165),
.A2(n_1108),
.A3(n_1198),
.B(n_1226),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1175),
.A2(n_1124),
.B(n_1194),
.C(n_1105),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1127),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1155),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1077),
.B(n_1083),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1208),
.A2(n_1096),
.B1(n_1113),
.B2(n_1122),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1207),
.A2(n_1209),
.B(n_1131),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1169),
.A2(n_1224),
.B(n_1185),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1106),
.A2(n_1231),
.B(n_1186),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1165),
.A2(n_1116),
.B(n_1184),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1139),
.B(n_1113),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1186),
.A2(n_1192),
.B(n_1136),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1164),
.A2(n_1172),
.B(n_1115),
.C(n_1119),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1181),
.A2(n_1217),
.B(n_1218),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1109),
.A2(n_1174),
.B(n_1097),
.C(n_1192),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1076),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1125),
.A2(n_1230),
.B(n_1138),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1232),
.A2(n_1236),
.B(n_1235),
.Y(n_1274)
);

AOI31xp67_ASAP7_75t_L g1275 ( 
.A1(n_1150),
.A2(n_1191),
.A3(n_1144),
.B(n_1148),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1187),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1238),
.A2(n_1171),
.A3(n_1141),
.B(n_1216),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1088),
.B(n_1128),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1141),
.A2(n_1126),
.B(n_1144),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1100),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1086),
.B(n_1081),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1200),
.A2(n_1148),
.B(n_1153),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1086),
.B(n_1081),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1151),
.A2(n_1176),
.B(n_1162),
.C(n_1214),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1201),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1126),
.A2(n_1094),
.B(n_1107),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1103),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1188),
.A2(n_1225),
.B(n_1223),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1111),
.A2(n_1195),
.B(n_1233),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1084),
.B(n_1177),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1135),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1202),
.A2(n_1114),
.B(n_1234),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1112),
.B(n_1189),
.C(n_1179),
.Y(n_1293)
);

AOI31xp67_ASAP7_75t_L g1294 ( 
.A1(n_1096),
.A2(n_1182),
.A3(n_1199),
.B(n_1228),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1147),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1202),
.A2(n_1114),
.B(n_1183),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1221),
.A2(n_1123),
.B(n_1219),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1190),
.A2(n_1193),
.B(n_1133),
.C(n_1203),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1204),
.A2(n_1210),
.B(n_1211),
.Y(n_1299)
);

AOI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1159),
.A2(n_1222),
.B(n_1229),
.Y(n_1300)
);

OAI21xp33_ASAP7_75t_L g1301 ( 
.A1(n_1142),
.A2(n_1080),
.B(n_1177),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1146),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1167),
.B(n_1177),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1193),
.A2(n_1156),
.B(n_1178),
.C(n_1168),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1220),
.A2(n_1161),
.B(n_1102),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1149),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1145),
.B(n_1173),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1104),
.B(n_1170),
.C(n_1163),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1157),
.A2(n_1197),
.B(n_1205),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1161),
.A2(n_1220),
.B(n_1212),
.Y(n_1310)
);

NOR2x1_ASAP7_75t_L g1311 ( 
.A(n_1137),
.B(n_1078),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_1091),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1102),
.A2(n_1163),
.B(n_1170),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1158),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1078),
.A2(n_1091),
.B(n_1092),
.C(n_1215),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1095),
.Y(n_1316)
);

AOI211xp5_ASAP7_75t_L g1317 ( 
.A1(n_1129),
.A2(n_1158),
.B(n_1196),
.C(n_1104),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1102),
.A2(n_1140),
.B(n_1104),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1078),
.A2(n_1140),
.B1(n_1227),
.B2(n_1213),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1158),
.A2(n_1227),
.B1(n_1163),
.B2(n_1170),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1130),
.A2(n_889),
.B(n_907),
.C(n_1090),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1130),
.A2(n_1237),
.B(n_1169),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1076),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1090),
.B(n_889),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1166),
.A2(n_1165),
.A3(n_1108),
.B(n_1198),
.Y(n_1325)
);

AOI221x1_ASAP7_75t_L g1326 ( 
.A1(n_1090),
.A2(n_972),
.B1(n_1120),
.B2(n_1172),
.C(n_1164),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1098),
.B(n_1086),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1132),
.B(n_889),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1090),
.A2(n_889),
.B1(n_907),
.B2(n_1143),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1117),
.A2(n_889),
.B(n_1090),
.C(n_728),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1085),
.Y(n_1335)
);

AO21x1_ASAP7_75t_L g1336 ( 
.A1(n_1117),
.A2(n_1143),
.B(n_1124),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1166),
.A2(n_1165),
.A3(n_1108),
.B(n_1198),
.Y(n_1337)
);

AOI221x1_ASAP7_75t_L g1338 ( 
.A1(n_1090),
.A2(n_972),
.B1(n_1120),
.B2(n_1172),
.C(n_1164),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1166),
.A2(n_1165),
.A3(n_1108),
.B(n_1198),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1079),
.A2(n_850),
.B1(n_826),
.B2(n_741),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1342)
);

INVx3_ASAP7_75t_SL g1343 ( 
.A(n_1095),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1090),
.A2(n_972),
.B1(n_585),
.B2(n_725),
.C(n_611),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1139),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1090),
.A2(n_889),
.B1(n_907),
.B2(n_1143),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1085),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1090),
.B(n_889),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1077),
.B(n_585),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1090),
.A2(n_889),
.B1(n_907),
.B2(n_1143),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1166),
.A2(n_1165),
.A3(n_1108),
.B(n_1198),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1117),
.A2(n_889),
.B(n_1090),
.C(n_728),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1132),
.B(n_889),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1090),
.B(n_889),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1077),
.B(n_889),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1085),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1076),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1098),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1166),
.A2(n_1165),
.A3(n_1108),
.B(n_1198),
.Y(n_1363)
);

AOI221x1_ASAP7_75t_L g1364 ( 
.A1(n_1090),
.A2(n_972),
.B1(n_1120),
.B2(n_1172),
.C(n_1164),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1132),
.Y(n_1366)
);

CKINVDCx11_ASAP7_75t_R g1367 ( 
.A(n_1167),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1077),
.B(n_889),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1077),
.B(n_585),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1132),
.B(n_889),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1090),
.A2(n_889),
.B(n_1101),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1167),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1166),
.A2(n_1165),
.A3(n_1108),
.B(n_1198),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1076),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1090),
.A2(n_889),
.B(n_1101),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1139),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1090),
.A2(n_889),
.B(n_585),
.C(n_956),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1090),
.A2(n_889),
.B(n_1101),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1082),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1077),
.B(n_585),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1095),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1077),
.B(n_596),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1117),
.A2(n_889),
.B(n_1090),
.C(n_728),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1098),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1132),
.B(n_889),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1132),
.B(n_720),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1237),
.A2(n_1169),
.B(n_1181),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_SL g1395 ( 
.A1(n_1090),
.A2(n_889),
.B(n_907),
.C(n_901),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1180),
.A2(n_1169),
.B(n_1217),
.Y(n_1396)
);

CKINVDCx8_ASAP7_75t_R g1397 ( 
.A(n_1095),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1085),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1089),
.A2(n_889),
.B(n_907),
.Y(n_1400)
);

AOI221x1_ASAP7_75t_L g1401 ( 
.A1(n_1090),
.A2(n_972),
.B1(n_1120),
.B2(n_1172),
.C(n_1164),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1085),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1180),
.A2(n_1169),
.B(n_1217),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1331),
.A2(n_1346),
.B1(n_1354),
.B2(n_1324),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1272),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1323),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1344),
.A2(n_1336),
.B1(n_1341),
.B2(n_1262),
.Y(n_1407)
);

BUFx4_ASAP7_75t_R g1408 ( 
.A(n_1316),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1331),
.A2(n_1346),
.B1(n_1354),
.B2(n_1350),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1361),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1251),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1251),
.Y(n_1412)
);

CKINVDCx6p67_ASAP7_75t_R g1413 ( 
.A(n_1367),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1397),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1239),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1370),
.A2(n_1387),
.B1(n_1324),
.B2(n_1349),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1301),
.A2(n_1358),
.B1(n_1349),
.B2(n_1393),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1358),
.A2(n_1254),
.B1(n_1317),
.B2(n_1293),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1267),
.Y(n_1419)
);

INVx11_ASAP7_75t_L g1420 ( 
.A(n_1343),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1301),
.A2(n_1254),
.B1(n_1290),
.B2(n_1359),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1281),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1327),
.Y(n_1423)
);

CKINVDCx6p67_ASAP7_75t_R g1424 ( 
.A(n_1377),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1259),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1317),
.A2(n_1293),
.B1(n_1372),
.B2(n_1378),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1369),
.A2(n_1385),
.B1(n_1295),
.B2(n_1291),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1260),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1335),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1388),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1280),
.A2(n_1287),
.B1(n_1306),
.B2(n_1261),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1333),
.A2(n_1356),
.B1(n_1390),
.B2(n_1258),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1347),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1329),
.A2(n_1371),
.B1(n_1392),
.B2(n_1357),
.Y(n_1434)
);

CKINVDCx14_ASAP7_75t_R g1435 ( 
.A(n_1373),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1372),
.A2(n_1378),
.B1(n_1383),
.B2(n_1320),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1383),
.B(n_1246),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1268),
.A2(n_1382),
.B1(n_1271),
.B2(n_1400),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1302),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1278),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1328),
.A2(n_1353),
.B1(n_1348),
.B2(n_1398),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1309),
.A2(n_1314),
.B1(n_1299),
.B2(n_1282),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1303),
.A2(n_1389),
.B1(n_1241),
.B2(n_1307),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_SL g1444 ( 
.A(n_1388),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1362),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1299),
.A2(n_1282),
.B1(n_1285),
.B2(n_1276),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1320),
.A2(n_1263),
.B1(n_1364),
.B2(n_1401),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1362),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1330),
.B(n_1332),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1360),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1345),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1283),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1399),
.A2(n_1402),
.B1(n_1263),
.B2(n_1283),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1380),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1391),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1334),
.A2(n_1374),
.B1(n_1365),
.B2(n_1342),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1304),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1381),
.A2(n_1269),
.B1(n_1284),
.B2(n_1244),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1391),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1244),
.A2(n_1292),
.B1(n_1326),
.B2(n_1338),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1255),
.A2(n_1265),
.B1(n_1294),
.B2(n_1312),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1319),
.A2(n_1297),
.B1(n_1310),
.B2(n_1255),
.Y(n_1462)
);

INVx2_ASAP7_75t_R g1463 ( 
.A(n_1300),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1296),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1310),
.A2(n_1255),
.B1(n_1305),
.B2(n_1286),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1391),
.A2(n_1248),
.B1(n_1274),
.B2(n_1308),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1248),
.A2(n_1308),
.B1(n_1250),
.B2(n_1313),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1279),
.A2(n_1298),
.B1(n_1247),
.B2(n_1256),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1289),
.A2(n_1249),
.B1(n_1245),
.B2(n_1264),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1395),
.A2(n_1266),
.B1(n_1273),
.B2(n_1321),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1266),
.A2(n_1273),
.B1(n_1288),
.B2(n_1253),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1315),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1318),
.B(n_1257),
.Y(n_1473)
);

CKINVDCx11_ASAP7_75t_R g1474 ( 
.A(n_1275),
.Y(n_1474)
);

BUFx8_ASAP7_75t_SL g1475 ( 
.A(n_1396),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1252),
.A2(n_1403),
.B1(n_1257),
.B2(n_1277),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1257),
.A2(n_1277),
.B1(n_1355),
.B2(n_1325),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1270),
.A2(n_1322),
.B1(n_1240),
.B2(n_1352),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1325),
.B(n_1363),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1243),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1339),
.A2(n_1386),
.B1(n_1384),
.B2(n_1379),
.Y(n_1481)
);

CKINVDCx11_ASAP7_75t_R g1482 ( 
.A(n_1325),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1337),
.B(n_1363),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1351),
.A2(n_1394),
.B1(n_1375),
.B2(n_1368),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1337),
.Y(n_1485)
);

INVx8_ASAP7_75t_L g1486 ( 
.A(n_1243),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1337),
.B(n_1340),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1340),
.A2(n_1355),
.B1(n_1363),
.B2(n_1376),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1340),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1243),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1355),
.Y(n_1491)
);

OAI21xp33_ASAP7_75t_L g1492 ( 
.A1(n_1376),
.A2(n_585),
.B(n_1258),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1376),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1242),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1242),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1344),
.A2(n_1003),
.B1(n_889),
.B2(n_1326),
.Y(n_1496)
);

BUFx10_ASAP7_75t_L g1497 ( 
.A(n_1303),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1327),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1367),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1367),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1327),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1366),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1239),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1344),
.A2(n_1003),
.B1(n_889),
.B2(n_1326),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1344),
.A2(n_1003),
.B1(n_889),
.B2(n_1326),
.Y(n_1505)
);

BUFx10_ASAP7_75t_L g1506 ( 
.A(n_1303),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1239),
.Y(n_1507)
);

OAI22x1_ASAP7_75t_L g1508 ( 
.A1(n_1350),
.A2(n_487),
.B1(n_1387),
.B2(n_1370),
.Y(n_1508)
);

BUFx8_ASAP7_75t_L g1509 ( 
.A(n_1373),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1327),
.Y(n_1510)
);

INVx6_ASAP7_75t_L g1511 ( 
.A(n_1251),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1331),
.A2(n_889),
.B1(n_1354),
.B2(n_1346),
.Y(n_1512)
);

BUFx4_ASAP7_75t_SL g1513 ( 
.A(n_1316),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1331),
.A2(n_889),
.B1(n_1354),
.B2(n_1346),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1344),
.A2(n_826),
.B1(n_487),
.B2(n_972),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1246),
.A2(n_1356),
.B(n_1333),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1344),
.A2(n_826),
.B1(n_487),
.B2(n_972),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1267),
.B(n_1132),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1344),
.A2(n_826),
.B1(n_487),
.B2(n_972),
.Y(n_1519)
);

CKINVDCx6p67_ASAP7_75t_R g1520 ( 
.A(n_1367),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1239),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1239),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1331),
.A2(n_889),
.B1(n_1354),
.B2(n_1346),
.Y(n_1523)
);

CKINVDCx6p67_ASAP7_75t_R g1524 ( 
.A(n_1367),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1239),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1239),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1344),
.A2(n_826),
.B1(n_487),
.B2(n_972),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1350),
.A2(n_1387),
.B1(n_1370),
.B2(n_1154),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1366),
.Y(n_1529)
);

BUFx10_ASAP7_75t_L g1530 ( 
.A(n_1303),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1344),
.A2(n_826),
.B1(n_487),
.B2(n_972),
.Y(n_1531)
);

INVx6_ASAP7_75t_L g1532 ( 
.A(n_1251),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1367),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_R g1534 ( 
.A1(n_1350),
.A2(n_818),
.B1(n_408),
.B2(n_388),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1272),
.Y(n_1535)
);

OAI21xp33_ASAP7_75t_L g1536 ( 
.A1(n_1258),
.A2(n_585),
.B(n_564),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1239),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1239),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1367),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1331),
.A2(n_1154),
.B1(n_411),
.B2(n_400),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1267),
.B(n_1132),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1344),
.A2(n_826),
.B1(n_487),
.B2(n_972),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1331),
.A2(n_889),
.B1(n_1354),
.B2(n_1346),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1311),
.B(n_1267),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1344),
.A2(n_826),
.B1(n_487),
.B2(n_972),
.Y(n_1545)
);

INVx6_ASAP7_75t_L g1546 ( 
.A(n_1251),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1331),
.A2(n_1154),
.B1(n_411),
.B2(n_400),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1493),
.Y(n_1548)
);

OR2x6_ASAP7_75t_L g1549 ( 
.A(n_1486),
.B(n_1473),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1479),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1434),
.B(n_1440),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1440),
.B(n_1416),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1483),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1479),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1487),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1487),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1512),
.A2(n_1523),
.B(n_1514),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1405),
.Y(n_1558)
);

AO21x2_ASAP7_75t_L g1559 ( 
.A1(n_1477),
.A2(n_1488),
.B(n_1492),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1485),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1436),
.B(n_1415),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1475),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1480),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1425),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1490),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1428),
.Y(n_1566)
);

CKINVDCx11_ASAP7_75t_R g1567 ( 
.A(n_1499),
.Y(n_1567)
);

AO21x1_ASAP7_75t_SL g1568 ( 
.A1(n_1437),
.A2(n_1516),
.B(n_1460),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1429),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1441),
.A2(n_1484),
.B(n_1481),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1433),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1502),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1512),
.A2(n_1523),
.B(n_1514),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1450),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1503),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1515),
.A2(n_1527),
.B1(n_1545),
.B2(n_1542),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1507),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1486),
.B(n_1491),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1521),
.Y(n_1580)
);

INVxp33_ASAP7_75t_L g1581 ( 
.A(n_1518),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1409),
.A2(n_1528),
.B1(n_1543),
.B2(n_1418),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1522),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1441),
.A2(n_1471),
.B(n_1476),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1490),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1525),
.B(n_1526),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1419),
.B(n_1437),
.Y(n_1587)
);

AOI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1449),
.A2(n_1438),
.B(n_1476),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1537),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1538),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1447),
.B(n_1426),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1489),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1454),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1491),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1494),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1410),
.B(n_1535),
.Y(n_1596)
);

BUFx4f_ASAP7_75t_SL g1597 ( 
.A(n_1500),
.Y(n_1597)
);

AO21x2_ASAP7_75t_L g1598 ( 
.A1(n_1488),
.A2(n_1449),
.B(n_1469),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1544),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1529),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1424),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1457),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1536),
.A2(n_1543),
.B1(n_1404),
.B2(n_1496),
.C(n_1504),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1464),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1495),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1442),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1547),
.A2(n_1540),
.B(n_1407),
.C(n_1531),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1404),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1482),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1474),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1517),
.A2(n_1519),
.B1(n_1508),
.B2(n_1534),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1435),
.B(n_1414),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1541),
.Y(n_1613)
);

AO21x2_ASAP7_75t_L g1614 ( 
.A1(n_1468),
.A2(n_1438),
.B(n_1467),
.Y(n_1614)
);

BUFx2_ASAP7_75t_SL g1615 ( 
.A(n_1444),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1446),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1458),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1458),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1468),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1516),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1465),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1417),
.B(n_1461),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1463),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1421),
.B(n_1462),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1432),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1478),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1423),
.B(n_1510),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1505),
.A2(n_1432),
.B1(n_1451),
.B2(n_1453),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1470),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1456),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1466),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1423),
.B(n_1510),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1427),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1455),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1443),
.B(n_1501),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1498),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1430),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1408),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1430),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1431),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1455),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1497),
.B(n_1530),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1411),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1406),
.A2(n_1472),
.B(n_1412),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1411),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1497),
.B(n_1530),
.Y(n_1646)
);

OA21x2_ASAP7_75t_L g1647 ( 
.A1(n_1445),
.A2(n_1546),
.B(n_1532),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1448),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1459),
.Y(n_1649)
);

INVx3_ASAP7_75t_SL g1650 ( 
.A(n_1511),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1506),
.Y(n_1651)
);

OAI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_1524),
.B2(n_1520),
.Y(n_1652)
);

AO32x2_ASAP7_75t_L g1653 ( 
.A1(n_1573),
.A2(n_1509),
.A3(n_1513),
.B1(n_1413),
.B2(n_1452),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1564),
.Y(n_1654)
);

A2O1A1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1607),
.A2(n_1452),
.B(n_1533),
.C(n_1439),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1613),
.B(n_1539),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1581),
.B(n_1509),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1549),
.B(n_1420),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1582),
.A2(n_1611),
.B1(n_1628),
.B2(n_1603),
.C(n_1577),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1584),
.A2(n_1571),
.B(n_1626),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1591),
.A2(n_1622),
.B(n_1574),
.C(n_1557),
.Y(n_1661)
);

AO21x2_ASAP7_75t_L g1662 ( 
.A1(n_1629),
.A2(n_1621),
.B(n_1623),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1591),
.A2(n_1620),
.B1(n_1624),
.B2(n_1625),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1617),
.A2(n_1618),
.B1(n_1561),
.B2(n_1608),
.C(n_1630),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1608),
.B(n_1617),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1618),
.B(n_1630),
.C(n_1619),
.Y(n_1666)
);

BUFx4f_ASAP7_75t_SL g1667 ( 
.A(n_1638),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1614),
.A2(n_1598),
.B(n_1619),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1567),
.Y(n_1669)
);

AND4x1_ASAP7_75t_L g1670 ( 
.A(n_1612),
.B(n_1596),
.C(n_1646),
.D(n_1642),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1573),
.B(n_1600),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1638),
.A2(n_1587),
.B1(n_1552),
.B2(n_1561),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1624),
.A2(n_1622),
.B1(n_1629),
.B2(n_1614),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1587),
.B(n_1638),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1549),
.B(n_1638),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1604),
.B(n_1550),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1610),
.A2(n_1562),
.B(n_1621),
.C(n_1602),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1604),
.B(n_1550),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1598),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1586),
.B(n_1563),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1623),
.A2(n_1606),
.B(n_1616),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1631),
.A2(n_1551),
.B1(n_1610),
.B2(n_1626),
.C(n_1562),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1616),
.A2(n_1614),
.B1(n_1631),
.B2(n_1606),
.C(n_1610),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1586),
.B(n_1632),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1610),
.A2(n_1593),
.B1(n_1635),
.B2(n_1651),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1555),
.B(n_1566),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1647),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1584),
.A2(n_1571),
.B(n_1588),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1646),
.B(n_1627),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1569),
.A2(n_1589),
.B1(n_1572),
.B2(n_1590),
.C(n_1583),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1569),
.B(n_1572),
.Y(n_1691)
);

NAND4xp25_ASAP7_75t_L g1692 ( 
.A(n_1575),
.B(n_1590),
.C(n_1578),
.D(n_1580),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1637),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1576),
.A2(n_1589),
.B1(n_1583),
.B2(n_1580),
.C(n_1578),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1597),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1559),
.A2(n_1579),
.B(n_1588),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1634),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1568),
.A2(n_1635),
.B(n_1605),
.C(n_1640),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1651),
.A2(n_1558),
.B1(n_1652),
.B2(n_1637),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1640),
.A2(n_1609),
.B(n_1633),
.C(n_1599),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1639),
.A2(n_1615),
.B1(n_1601),
.B2(n_1650),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1648),
.Y(n_1702)
);

AO32x2_ASAP7_75t_L g1703 ( 
.A1(n_1553),
.A2(n_1556),
.A3(n_1554),
.B1(n_1633),
.B2(n_1559),
.Y(n_1703)
);

AND2x2_ASAP7_75t_SL g1704 ( 
.A(n_1644),
.B(n_1595),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1645),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1560),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1676),
.B(n_1559),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1706),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1659),
.A2(n_1644),
.B1(n_1592),
.B2(n_1560),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1706),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1661),
.B(n_1636),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1684),
.B(n_1680),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1676),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1654),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1678),
.B(n_1548),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1688),
.B(n_1594),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1687),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1686),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1691),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1678),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1664),
.B(n_1636),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1659),
.A2(n_1644),
.B1(n_1553),
.B2(n_1570),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1660),
.B(n_1585),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1665),
.B(n_1641),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1675),
.B(n_1565),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1703),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1670),
.B(n_1692),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1672),
.B(n_1643),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1679),
.Y(n_1730)
);

INVxp33_ASAP7_75t_SL g1731 ( 
.A(n_1669),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1660),
.B(n_1565),
.Y(n_1732)
);

OAI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1655),
.A2(n_1664),
.B1(n_1673),
.B2(n_1663),
.C(n_1683),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1690),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1671),
.Y(n_1735)
);

OAI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1733),
.A2(n_1683),
.B1(n_1698),
.B2(n_1682),
.C(n_1666),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1713),
.B(n_1668),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1712),
.B(n_1674),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1733),
.A2(n_1698),
.B1(n_1682),
.B2(n_1700),
.C(n_1677),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1710),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1712),
.B(n_1689),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1708),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1708),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1707),
.B(n_1697),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1707),
.B(n_1702),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1713),
.B(n_1685),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_L g1747 ( 
.A(n_1734),
.B(n_1730),
.C(n_1728),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1714),
.Y(n_1748)
);

AOI211xp5_ASAP7_75t_L g1749 ( 
.A1(n_1728),
.A2(n_1734),
.B(n_1711),
.C(n_1722),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1732),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1721),
.B(n_1662),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1734),
.A2(n_1722),
.B(n_1711),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1709),
.A2(n_1696),
.B(n_1700),
.C(n_1699),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1732),
.Y(n_1754)
);

INVx5_ASAP7_75t_SL g1755 ( 
.A(n_1726),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_L g1756 ( 
.A(n_1715),
.B(n_1658),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1709),
.A2(n_1662),
.B1(n_1644),
.B2(n_1681),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1721),
.B(n_1681),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1718),
.B(n_1690),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1729),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1717),
.B(n_1704),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1716),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_L g1763 ( 
.A(n_1730),
.B(n_1694),
.C(n_1696),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1748),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1745),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1750),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1737),
.B(n_1715),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1745),
.Y(n_1768)
);

NOR4xp25_ASAP7_75t_SL g1769 ( 
.A(n_1736),
.B(n_1705),
.C(n_1653),
.D(n_1649),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1748),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1743),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1750),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1731),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1715),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1755),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1761),
.B(n_1719),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1759),
.B(n_1719),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1759),
.B(n_1725),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1760),
.B(n_1720),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1743),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1750),
.B(n_1724),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1742),
.B(n_1720),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1740),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1754),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1744),
.B(n_1725),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1743),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1744),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1762),
.B(n_1724),
.Y(n_1788)
);

INVxp67_ASAP7_75t_SL g1789 ( 
.A(n_1763),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1789),
.B(n_1749),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1764),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1764),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1764),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1770),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1775),
.B(n_1756),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1789),
.B(n_1777),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1770),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1770),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1771),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1773),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1775),
.B(n_1756),
.Y(n_1801)
);

INVxp67_ASAP7_75t_SL g1802 ( 
.A(n_1773),
.Y(n_1802)
);

OAI31xp67_ASAP7_75t_L g1803 ( 
.A1(n_1783),
.A2(n_1762),
.A3(n_1747),
.B(n_1731),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1771),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1769),
.A2(n_1736),
.B1(n_1749),
.B2(n_1747),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1771),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1775),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1775),
.B(n_1741),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1780),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1775),
.B(n_1741),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1780),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1775),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1783),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1781),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1778),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1780),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1786),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1777),
.B(n_1695),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1765),
.B(n_1741),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1778),
.B(n_1744),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1781),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1786),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1765),
.B(n_1738),
.Y(n_1823)
);

INVxp33_ASAP7_75t_L g1824 ( 
.A(n_1778),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1768),
.B(n_1738),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1787),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_L g1828 ( 
.A(n_1783),
.B(n_1656),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1785),
.Y(n_1829)
);

AND4x1_ASAP7_75t_L g1830 ( 
.A(n_1769),
.B(n_1752),
.C(n_1763),
.D(n_1729),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1768),
.B(n_1738),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1787),
.B(n_1752),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1776),
.B(n_1735),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1790),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1815),
.B(n_1779),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1814),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1814),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1800),
.B(n_1779),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1813),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1796),
.B(n_1767),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1802),
.B(n_1746),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1830),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1808),
.B(n_1776),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1808),
.B(n_1776),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1829),
.B(n_1767),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1805),
.B(n_1746),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1829),
.B(n_1767),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1791),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1824),
.B(n_1774),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1813),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1821),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1791),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1792),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1833),
.B(n_1827),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1807),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1820),
.B(n_1774),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1792),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1833),
.B(n_1774),
.Y(n_1859)
);

INVxp67_ASAP7_75t_SL g1860 ( 
.A(n_1828),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1833),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1833),
.B(n_1782),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1807),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1810),
.B(n_1788),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1810),
.B(n_1788),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1818),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1812),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1827),
.B(n_1782),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1793),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1819),
.B(n_1788),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1793),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1849),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1843),
.A2(n_1739),
.B1(n_1753),
.B2(n_1757),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1844),
.B(n_1819),
.Y(n_1874)
);

O2A1O1Ixp5_ASAP7_75t_L g1875 ( 
.A1(n_1847),
.A2(n_1803),
.B(n_1831),
.C(n_1801),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1849),
.Y(n_1876)
);

NAND4xp25_ASAP7_75t_L g1877 ( 
.A(n_1839),
.B(n_1803),
.C(n_1831),
.D(n_1801),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1860),
.A2(n_1769),
.B(n_1739),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1861),
.Y(n_1879)
);

AND2x2_ASAP7_75t_SL g1880 ( 
.A(n_1840),
.B(n_1795),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1835),
.A2(n_1861),
.B1(n_1859),
.B2(n_1862),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1835),
.B(n_1823),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1842),
.B(n_1840),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1853),
.Y(n_1884)
);

AOI332xp33_ASAP7_75t_L g1885 ( 
.A1(n_1841),
.A2(n_1797),
.A3(n_1798),
.B1(n_1794),
.B2(n_1825),
.B3(n_1817),
.C1(n_1822),
.C2(n_1799),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1844),
.B(n_1823),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1866),
.A2(n_1832),
.B1(n_1826),
.B2(n_1746),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_SL g1888 ( 
.A1(n_1859),
.A2(n_1753),
.B1(n_1795),
.B2(n_1727),
.Y(n_1888)
);

NOR3x1_ASAP7_75t_L g1889 ( 
.A(n_1850),
.B(n_1812),
.C(n_1820),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1845),
.B(n_1826),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1864),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1853),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1854),
.Y(n_1893)
);

OAI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1862),
.A2(n_1751),
.B1(n_1821),
.B2(n_1758),
.Y(n_1894)
);

NOR2xp67_ASAP7_75t_SL g1895 ( 
.A(n_1851),
.B(n_1693),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1845),
.B(n_1832),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1855),
.A2(n_1866),
.B(n_1836),
.C(n_1841),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1879),
.B(n_1855),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1891),
.Y(n_1899)
);

OAI21xp33_ASAP7_75t_L g1900 ( 
.A1(n_1888),
.A2(n_1850),
.B(n_1846),
.Y(n_1900)
);

AOI21xp33_ASAP7_75t_SL g1901 ( 
.A1(n_1880),
.A2(n_1848),
.B(n_1856),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1879),
.B(n_1857),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1882),
.B(n_1881),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1892),
.Y(n_1904)
);

AOI32xp33_ASAP7_75t_L g1905 ( 
.A1(n_1887),
.A2(n_1836),
.A3(n_1846),
.B1(n_1870),
.B2(n_1865),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1873),
.A2(n_1848),
.B1(n_1857),
.B2(n_1867),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1874),
.B(n_1870),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1892),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1891),
.B(n_1864),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1874),
.B(n_1865),
.Y(n_1910)
);

OAI32xp33_ASAP7_75t_L g1911 ( 
.A1(n_1877),
.A2(n_1868),
.A3(n_1869),
.B1(n_1871),
.B2(n_1854),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1893),
.Y(n_1912)
);

AOI21xp33_ASAP7_75t_L g1913 ( 
.A1(n_1897),
.A2(n_1838),
.B(n_1837),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1878),
.A2(n_1867),
.B1(n_1856),
.B2(n_1863),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1893),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1880),
.A2(n_1852),
.B1(n_1838),
.B2(n_1837),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1872),
.Y(n_1917)
);

AO221x1_ASAP7_75t_L g1918 ( 
.A1(n_1885),
.A2(n_1837),
.B1(n_1852),
.B2(n_1838),
.C(n_1858),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1907),
.B(n_1883),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1902),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1910),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1918),
.B(n_1886),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1909),
.Y(n_1923)
);

OAI21xp33_ASAP7_75t_L g1924 ( 
.A1(n_1900),
.A2(n_1890),
.B(n_1886),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1899),
.Y(n_1925)
);

AOI21xp33_ASAP7_75t_L g1926 ( 
.A1(n_1914),
.A2(n_1884),
.B(n_1876),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1898),
.B(n_1890),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1904),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1901),
.B(n_1896),
.Y(n_1929)
);

OAI211xp5_ASAP7_75t_L g1930 ( 
.A1(n_1922),
.A2(n_1911),
.B(n_1916),
.C(n_1903),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1927),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1927),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1919),
.B(n_1906),
.Y(n_1933)
);

NAND3xp33_ASAP7_75t_L g1934 ( 
.A(n_1926),
.B(n_1914),
.C(n_1906),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1922),
.A2(n_1913),
.B1(n_1895),
.B2(n_1852),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1920),
.B(n_1905),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1928),
.B(n_1908),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1924),
.A2(n_1875),
.B(n_1917),
.Y(n_1938)
);

NAND3xp33_ASAP7_75t_L g1939 ( 
.A(n_1934),
.B(n_1925),
.C(n_1923),
.Y(n_1939)
);

OAI21xp5_ASAP7_75t_SL g1940 ( 
.A1(n_1930),
.A2(n_1929),
.B(n_1921),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1933),
.A2(n_1929),
.B(n_1915),
.Y(n_1941)
);

AOI221xp5_ASAP7_75t_L g1942 ( 
.A1(n_1935),
.A2(n_1912),
.B1(n_1894),
.B2(n_1869),
.C(n_1871),
.Y(n_1942)
);

OAI211xp5_ASAP7_75t_L g1943 ( 
.A1(n_1938),
.A2(n_1889),
.B(n_1896),
.C(n_1863),
.Y(n_1943)
);

NAND4xp25_ASAP7_75t_SL g1944 ( 
.A(n_1943),
.B(n_1932),
.C(n_1941),
.D(n_1939),
.Y(n_1944)
);

NOR3xp33_ASAP7_75t_L g1945 ( 
.A(n_1940),
.B(n_1936),
.C(n_1931),
.Y(n_1945)
);

AOI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1942),
.A2(n_1858),
.B1(n_1895),
.B2(n_1937),
.C(n_1868),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1940),
.A2(n_1657),
.B1(n_1781),
.B2(n_1794),
.Y(n_1947)
);

AOI221xp5_ASAP7_75t_L g1948 ( 
.A1(n_1940),
.A2(n_1797),
.B1(n_1798),
.B2(n_1822),
.C(n_1817),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1943),
.B(n_1799),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1945),
.B(n_1834),
.Y(n_1950)
);

XNOR2xp5_ASAP7_75t_L g1951 ( 
.A(n_1946),
.B(n_1701),
.Y(n_1951)
);

NOR2x1_ASAP7_75t_L g1952 ( 
.A(n_1944),
.B(n_1804),
.Y(n_1952)
);

XOR2xp5_ASAP7_75t_L g1953 ( 
.A(n_1947),
.B(n_1723),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1949),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1950),
.B(n_1804),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1952),
.B(n_1948),
.Y(n_1956)
);

NAND4xp75_ASAP7_75t_L g1957 ( 
.A(n_1954),
.B(n_1834),
.C(n_1653),
.D(n_1816),
.Y(n_1957)
);

AOI22x1_ASAP7_75t_L g1958 ( 
.A1(n_1955),
.A2(n_1951),
.B1(n_1956),
.B2(n_1953),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1958),
.A2(n_1957),
.B1(n_1825),
.B2(n_1816),
.Y(n_1959)
);

OAI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1959),
.A2(n_1811),
.B1(n_1809),
.B2(n_1806),
.Y(n_1960)
);

NAND2x1_ASAP7_75t_L g1961 ( 
.A(n_1959),
.B(n_1806),
.Y(n_1961)
);

AO22x2_ASAP7_75t_L g1962 ( 
.A1(n_1960),
.A2(n_1811),
.B1(n_1809),
.B2(n_1772),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1961),
.A2(n_1653),
.B1(n_1667),
.B2(n_1781),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1963),
.A2(n_1766),
.B1(n_1772),
.B2(n_1784),
.Y(n_1964)
);

NAND3x1_ASAP7_75t_SL g1965 ( 
.A(n_1964),
.B(n_1962),
.C(n_1653),
.Y(n_1965)
);

XNOR2xp5_ASAP7_75t_L g1966 ( 
.A(n_1965),
.B(n_1658),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1966),
.Y(n_1967)
);

OAI221xp5_ASAP7_75t_R g1968 ( 
.A1(n_1967),
.A2(n_1757),
.B1(n_1667),
.B2(n_1785),
.C(n_1740),
.Y(n_1968)
);

AOI211xp5_ASAP7_75t_L g1969 ( 
.A1(n_1968),
.A2(n_1772),
.B(n_1784),
.C(n_1766),
.Y(n_1969)
);


endmodule