module fake_jpeg_17812_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_59),
.Y(n_63)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_52),
.B1(n_51),
.B2(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_52),
.B1(n_55),
.B2(n_62),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_53),
.B1(n_47),
.B2(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_76),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_47),
.B1(n_49),
.B2(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_41),
.B1(n_15),
.B2(n_16),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_49),
.B1(n_41),
.B2(n_2),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_81),
.B1(n_86),
.B2(n_5),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_50),
.B(n_58),
.C(n_44),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_5),
.B(n_6),
.Y(n_95)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_89),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_50),
.B1(n_44),
.B2(n_4),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_92),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_2),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_4),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_93),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_88),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_109),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_14),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_32),
.A3(n_19),
.B1(n_20),
.B2(n_22),
.C(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_34),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_82),
.B(n_101),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_116),
.A2(n_105),
.B1(n_104),
.B2(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_114),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_103),
.A3(n_104),
.B1(n_97),
.B2(n_9),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_122),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_27),
.B(n_28),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_29),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_30),
.B(n_31),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_35),
.B(n_36),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_37),
.Y(n_131)
);


endmodule