module real_jpeg_1924_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_0),
.Y(n_115)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_1),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_35),
.B1(n_37),
.B2(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_55),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_2),
.A2(n_55),
.B1(n_66),
.B2(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_4),
.A2(n_35),
.B1(n_37),
.B2(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_47),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_4),
.A2(n_47),
.B1(n_66),
.B2(n_69),
.Y(n_171)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_147),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_147),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_66),
.B1(n_69),
.B2(n_147),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_7),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_35),
.B1(n_37),
.B2(n_80),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_80),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_7),
.A2(n_66),
.B1(n_69),
.B2(n_80),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_35),
.B1(n_37),
.B2(n_88),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_88),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_66),
.B1(n_69),
.B2(n_88),
.Y(n_192)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_10),
.A2(n_35),
.B1(n_37),
.B2(n_178),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_178),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_10),
.A2(n_66),
.B1(n_69),
.B2(n_178),
.Y(n_263)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_13),
.B(n_56),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_13),
.B(n_29),
.C(n_31),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_13),
.B(n_28),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_13),
.B(n_63),
.C(n_66),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_13),
.B(n_115),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_13),
.B(n_70),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_213),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g344 ( 
.A(n_14),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_14),
.B(n_346),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_15),
.A2(n_35),
.B1(n_37),
.B2(n_125),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_125),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_15),
.A2(n_66),
.B1(n_69),
.B2(n_125),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_16),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_40),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_16),
.A2(n_40),
.B1(n_66),
.B2(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_16),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_344),
.B(n_345),
.Y(n_19)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_339),
.B(n_342),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_331),
.B(n_335),
.Y(n_21)
);

AOI21x1_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_93),
.B(n_330),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_81),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_24),
.B(n_81),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_59),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_25)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_27),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_28),
.B(n_175),
.Y(n_279)
);

AO22x1_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_30),
.A2(n_31),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_31),
.B(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_35),
.B(n_203),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_35),
.B(n_51),
.Y(n_227)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g225 ( 
.A1(n_37),
.A2(n_45),
.A3(n_50),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_41),
.B(n_57),
.C(n_59),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_54),
.B2(n_56),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_49),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_45),
.A2(n_78),
.B(n_213),
.C(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_45),
.B(n_213),
.Y(n_214)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_48),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_48),
.A2(n_56),
.B1(n_146),
.B2(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_48),
.A2(n_54),
.B1(n_56),
.B2(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_48),
.A2(n_56),
.B(n_333),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_78),
.B1(n_79),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_49),
.A2(n_87),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_49),
.B(n_124),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_49),
.A2(n_122),
.B(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_73),
.C(n_77),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_73),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_86),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_105)
);

OAI21x1_ASAP7_75t_R g60 ( 
.A1(n_61),
.A2(n_70),
.B(n_71),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_61),
.A2(n_70),
.B1(n_120),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_61),
.A2(n_70),
.B1(n_141),
.B2(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_61),
.A2(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_61),
.B(n_199),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_72),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_101),
.B1(n_102),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_65),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_65),
.A2(n_220),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_65),
.A2(n_101),
.B1(n_196),
.B2(n_246),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_66),
.B(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_70),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_76),
.B1(n_92),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_74),
.A2(n_76),
.B1(n_99),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_74),
.A2(n_76),
.B1(n_186),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_74),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_74),
.A2(n_217),
.B(n_279),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_76),
.A2(n_143),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_76),
.A2(n_174),
.B(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_78),
.A2(n_145),
.B(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_86),
.B1(n_104),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_154),
.B(n_327),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_150),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_126),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_96),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_96),
.B(n_126),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_96),
.B(n_151),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_103),
.CI(n_107),
.CON(n_96),
.SN(n_96)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_101),
.A2(n_198),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_121),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_109),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_111),
.B1(n_121),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_110),
.A2(n_111),
.B1(n_118),
.B2(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_115),
.B(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_112),
.A2(n_115),
.B1(n_138),
.B2(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_112),
.A2(n_213),
.B(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_113),
.A2(n_114),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_113),
.B(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_113),
.A2(n_114),
.B1(n_193),
.B2(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_113),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_113),
.A2(n_114),
.B1(n_238),
.B2(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_114),
.A2(n_192),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_114),
.B(n_207),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_115),
.A2(n_206),
.B(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_118),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_133),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_142),
.C(n_144),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_135),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_136),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_144),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_149),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_150),
.A2(n_328),
.B(n_329),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_179),
.B(n_326),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_156),
.B(n_159),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_160),
.B(n_163),
.Y(n_324)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_165),
.B(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.C(n_176),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_166),
.A2(n_167),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_168),
.B(n_170),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_169),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_176),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_177),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_321),
.B(n_325),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_290),
.B(n_318),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_232),
.B(n_289),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_208),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_183),
.B(n_208),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.C(n_200),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_184),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_188),
.C(n_191),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_194),
.B(n_200),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_222),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_209),
.B(n_223),
.C(n_231),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_221),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_210),
.B(n_216),
.C(n_218),
.Y(n_303)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_224),
.B(n_229),
.Y(n_294)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_284),
.B(n_288),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_273),
.B(n_283),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_255),
.B(n_272),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_249),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_249),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_241),
.B1(n_247),
.B2(n_248),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_244),
.C(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_266),
.B(n_271),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_264),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_305),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_304),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_304),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_302),
.C(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_296),
.C(n_300),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_317),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_317),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_311),
.C(n_313),
.Y(n_322)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_332),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_337),
.B(n_341),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);


endmodule