module real_aes_6701_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g475 ( .A1(n_0), .A2(n_179), .B(n_476), .C(n_479), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_1), .B(n_470), .Y(n_481) );
INVx1_ASAP7_75t_L g118 ( .A(n_2), .Y(n_118) );
AOI22xp33_ASAP7_75t_SL g105 ( .A1(n_3), .A2(n_106), .B1(n_767), .B2(n_777), .Y(n_105) );
INVx1_ASAP7_75t_L g228 ( .A(n_4), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_5), .B(n_167), .Y(n_504) );
XNOR2xp5_ASAP7_75t_SL g763 ( .A(n_6), .B(n_103), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_7), .A2(n_454), .B(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_8), .A2(n_11), .B1(n_437), .B2(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_8), .Y(n_759) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_9), .A2(n_184), .B(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_10), .A2(n_41), .B1(n_140), .B2(n_152), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_11), .A2(n_124), .B1(n_125), .B2(n_437), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_11), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_12), .B(n_184), .Y(n_217) );
AND2x6_ASAP7_75t_L g155 ( .A(n_13), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_14), .A2(n_155), .B(n_457), .C(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_15), .B(n_42), .Y(n_119) );
INVx1_ASAP7_75t_L g772 ( .A(n_15), .Y(n_772) );
INVx1_ASAP7_75t_L g136 ( .A(n_16), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_17), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g222 ( .A(n_18), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_19), .B(n_167), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_20), .B(n_182), .Y(n_200) );
AO32x2_ASAP7_75t_L g176 ( .A1(n_21), .A2(n_177), .A3(n_181), .B1(n_183), .B2(n_184), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_22), .A2(n_60), .B1(n_743), .B2(n_744), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_22), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_23), .B(n_140), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_24), .B(n_182), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_25), .A2(n_58), .B1(n_140), .B2(n_152), .Y(n_180) );
AOI22xp33_ASAP7_75t_SL g193 ( .A1(n_26), .A2(n_85), .B1(n_140), .B2(n_144), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_27), .B(n_140), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_28), .A2(n_183), .B(n_457), .C(n_459), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_29), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_30), .A2(n_183), .B(n_457), .C(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_31), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_32), .B(n_132), .Y(n_242) );
AOI222xp33_ASAP7_75t_L g120 ( .A1(n_33), .A2(n_121), .B1(n_736), .B2(n_737), .C1(n_746), .C2(n_749), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_34), .A2(n_454), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_35), .B(n_132), .Y(n_174) );
INVx2_ASAP7_75t_L g142 ( .A(n_36), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_37), .A2(n_488), .B(n_489), .C(n_493), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_38), .B(n_140), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_39), .B(n_132), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_40), .B(n_147), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_42), .B(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_43), .B(n_453), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_44), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_45), .B(n_167), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_46), .B(n_454), .Y(n_534) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_47), .A2(n_738), .B1(n_739), .B2(n_745), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_47), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_48), .A2(n_488), .B(n_493), .C(n_515), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_49), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_49), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_50), .B(n_140), .Y(n_210) );
INVx1_ASAP7_75t_L g477 ( .A(n_51), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_52), .A2(n_94), .B1(n_152), .B2(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g516 ( .A(n_53), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_54), .B(n_140), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_55), .B(n_140), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_56), .B(n_454), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_57), .B(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_59), .A2(n_64), .B1(n_140), .B2(n_144), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_60), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_61), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_62), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_63), .B(n_140), .Y(n_241) );
INVx1_ASAP7_75t_L g156 ( .A(n_65), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_66), .B(n_454), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_67), .B(n_470), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_68), .A2(n_215), .B(n_225), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_69), .B(n_140), .Y(n_229) );
INVx1_ASAP7_75t_L g135 ( .A(n_70), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_71), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_72), .B(n_167), .Y(n_491) );
AO32x2_ASAP7_75t_L g189 ( .A1(n_73), .A2(n_183), .A3(n_184), .B1(n_190), .B2(n_194), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_74), .B(n_168), .Y(n_547) );
INVx1_ASAP7_75t_L g240 ( .A(n_75), .Y(n_240) );
INVx1_ASAP7_75t_L g165 ( .A(n_76), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_77), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_78), .B(n_461), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_79), .A2(n_457), .B(n_493), .C(n_502), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_80), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_80), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_81), .B(n_144), .Y(n_166) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_82), .Y(n_525) );
INVx1_ASAP7_75t_L g776 ( .A(n_83), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_84), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_86), .B(n_152), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_87), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_88), .B(n_144), .Y(n_171) );
INVx2_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_90), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_91), .B(n_154), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_92), .B(n_144), .Y(n_211) );
OR2x2_ASAP7_75t_L g115 ( .A(n_93), .B(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g440 ( .A(n_93), .B(n_117), .Y(n_440) );
INVx2_ASAP7_75t_L g735 ( .A(n_93), .Y(n_735) );
NAND3xp33_ASAP7_75t_SL g773 ( .A(n_93), .B(n_118), .C(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_95), .A2(n_104), .B1(n_144), .B2(n_145), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_96), .B(n_454), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_97), .Y(n_490) );
INVxp67_ASAP7_75t_L g528 ( .A(n_98), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_99), .B(n_144), .Y(n_238) );
INVx1_ASAP7_75t_L g503 ( .A(n_100), .Y(n_503) );
INVx1_ASAP7_75t_L g543 ( .A(n_101), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_102), .B(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g518 ( .A(n_103), .B(n_132), .Y(n_518) );
AOI22x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_110), .B1(n_120), .B2(n_751), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_111), .A2(n_752), .B(n_765), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g766 ( .A(n_115), .Y(n_766) );
NOR2x2_ASAP7_75t_L g748 ( .A(n_116), .B(n_735), .Y(n_748) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g734 ( .A(n_117), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
OAI22x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_438), .B1(n_441), .B2(n_732), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_123), .A2(n_442), .B1(n_732), .B2(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_124), .A2(n_125), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_359), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_278), .C(n_293), .D(n_319), .E(n_341), .Y(n_126) );
NOR2xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_258), .Y(n_127) );
OAI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_195), .B1(n_231), .B2(n_247), .C(n_248), .Y(n_128) );
NOR2xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_185), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_130), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g435 ( .A(n_130), .Y(n_435) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_158), .Y(n_130) );
INVx1_ASAP7_75t_L g275 ( .A(n_131), .Y(n_275) );
AND2x2_ASAP7_75t_L g277 ( .A(n_131), .B(n_176), .Y(n_277) );
AND2x2_ASAP7_75t_L g287 ( .A(n_131), .B(n_175), .Y(n_287) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_131), .Y(n_305) );
INVx1_ASAP7_75t_L g315 ( .A(n_131), .Y(n_315) );
OR2x2_ASAP7_75t_L g353 ( .A(n_131), .B(n_252), .Y(n_353) );
INVx2_ASAP7_75t_L g403 ( .A(n_131), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_131), .B(n_251), .Y(n_420) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_137), .B(n_157), .Y(n_131) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_132), .A2(n_162), .B(n_174), .Y(n_161) );
INVx2_ASAP7_75t_L g194 ( .A(n_132), .Y(n_194) );
INVx1_ASAP7_75t_L g467 ( .A(n_132), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_132), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_132), .A2(n_513), .B(n_514), .Y(n_512) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_L g182 ( .A(n_133), .B(n_134), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_149), .B(n_155), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_146), .Y(n_138) );
INVx3_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_140), .Y(n_505) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
BUFx3_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
AND2x6_ASAP7_75t_L g457 ( .A(n_141), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
INVx1_ASAP7_75t_L g216 ( .A(n_142), .Y(n_216) );
INVx2_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx3_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
AND2x2_ASAP7_75t_L g455 ( .A(n_148), .B(n_216), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_148), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_153), .Y(n_149) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_153), .A2(n_227), .B(n_240), .C(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_154), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_177) );
OAI22xp5_ASAP7_75t_SL g190 ( .A1(n_154), .A2(n_168), .B1(n_191), .B2(n_193), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_154), .A2(n_179), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx4_ASAP7_75t_L g478 ( .A(n_154), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g162 ( .A1(n_155), .A2(n_163), .B(n_169), .Y(n_162) );
BUFx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_155), .A2(n_209), .B(n_212), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_155), .A2(n_221), .B(n_226), .Y(n_220) );
AND2x4_ASAP7_75t_L g454 ( .A(n_155), .B(n_455), .Y(n_454) );
INVx4_ASAP7_75t_SL g480 ( .A(n_155), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_155), .B(n_455), .Y(n_544) );
NOR2xp67_ASAP7_75t_L g158 ( .A(n_159), .B(n_175), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_160), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_160), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_160), .B(n_275), .Y(n_335) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
INVx2_ASAP7_75t_L g252 ( .A(n_161), .Y(n_252) );
OR2x2_ASAP7_75t_L g314 ( .A(n_161), .B(n_315), .Y(n_314) );
O2A1O1Ixp5_ASAP7_75t_SL g163 ( .A1(n_164), .A2(n_165), .B(n_166), .C(n_167), .Y(n_163) );
INVx2_ASAP7_75t_L g179 ( .A(n_167), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_167), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_167), .A2(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_167), .B(n_528), .Y(n_527) );
INVx5_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_172), .Y(n_169) );
INVx1_ASAP7_75t_L g225 ( .A(n_172), .Y(n_225) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g461 ( .A(n_173), .Y(n_461) );
AND2x2_ASAP7_75t_L g253 ( .A(n_175), .B(n_189), .Y(n_253) );
AND2x2_ASAP7_75t_L g270 ( .A(n_175), .B(n_250), .Y(n_270) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g188 ( .A(n_176), .B(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g273 ( .A(n_176), .Y(n_273) );
AND2x2_ASAP7_75t_L g402 ( .A(n_176), .B(n_403), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_179), .A2(n_213), .B(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_179), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
INVx2_ASAP7_75t_L g219 ( .A(n_181), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_181), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_182), .Y(n_184) );
NAND3xp33_ASAP7_75t_L g201 ( .A(n_183), .B(n_202), .C(n_205), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_183), .A2(n_236), .B(n_239), .Y(n_235) );
INVx4_ASAP7_75t_L g205 ( .A(n_184), .Y(n_205) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_184), .A2(n_208), .B(n_217), .Y(n_207) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_184), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_184), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g247 ( .A(n_185), .Y(n_247) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
AND2x2_ASAP7_75t_L g365 ( .A(n_186), .B(n_253), .Y(n_365) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g366 ( .A(n_187), .B(n_277), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_188), .A2(n_334), .B(n_336), .C(n_338), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_188), .B(n_334), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_188), .A2(n_264), .B1(n_407), .B2(n_408), .C(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g250 ( .A(n_189), .Y(n_250) );
INVx1_ASAP7_75t_L g286 ( .A(n_189), .Y(n_286) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_189), .Y(n_295) );
INVx2_ASAP7_75t_L g479 ( .A(n_192), .Y(n_479) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_192), .Y(n_492) );
INVx1_ASAP7_75t_L g464 ( .A(n_194), .Y(n_464) );
INVx1_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
AND2x2_ASAP7_75t_L g312 ( .A(n_197), .B(n_257), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_197), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_198), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g404 ( .A(n_198), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g436 ( .A(n_198), .Y(n_436) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g266 ( .A(n_199), .Y(n_266) );
AND2x2_ASAP7_75t_L g292 ( .A(n_199), .B(n_246), .Y(n_292) );
NOR2x1_ASAP7_75t_L g301 ( .A(n_199), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g308 ( .A(n_199), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
AO21x1_ASAP7_75t_L g243 ( .A1(n_202), .A2(n_205), .B(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g470 ( .A(n_205), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_205), .B(n_495), .Y(n_494) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_205), .A2(n_500), .B(n_507), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_205), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_205), .A2(n_542), .B(n_549), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_206), .B(n_348), .Y(n_383) );
INVx1_ASAP7_75t_SL g387 ( .A(n_206), .Y(n_387) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_218), .Y(n_206) );
INVx3_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
AND2x2_ASAP7_75t_L g257 ( .A(n_207), .B(n_234), .Y(n_257) );
AND2x2_ASAP7_75t_L g279 ( .A(n_207), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g324 ( .A(n_207), .B(n_318), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_207), .B(n_256), .Y(n_405) );
INVx2_ASAP7_75t_L g227 ( .A(n_215), .Y(n_227) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g245 ( .A(n_218), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g256 ( .A(n_218), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_218), .B(n_234), .Y(n_281) );
AND2x2_ASAP7_75t_L g317 ( .A(n_218), .B(n_318), .Y(n_317) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_230), .Y(n_218) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_219), .A2(n_235), .B(n_242), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .C(n_225), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_223), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_223), .A2(n_547), .B(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_225), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_227), .A2(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_245), .Y(n_232) );
INVx1_ASAP7_75t_L g297 ( .A(n_233), .Y(n_297) );
AND2x2_ASAP7_75t_L g339 ( .A(n_233), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_233), .B(n_260), .Y(n_345) );
AOI21xp5_ASAP7_75t_SL g419 ( .A1(n_233), .A2(n_251), .B(n_274), .Y(n_419) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_243), .Y(n_233) );
OR2x2_ASAP7_75t_L g262 ( .A(n_234), .B(n_243), .Y(n_262) );
AND2x2_ASAP7_75t_L g309 ( .A(n_234), .B(n_246), .Y(n_309) );
INVx2_ASAP7_75t_L g318 ( .A(n_234), .Y(n_318) );
INVx1_ASAP7_75t_L g424 ( .A(n_234), .Y(n_424) );
AND2x2_ASAP7_75t_L g348 ( .A(n_243), .B(n_318), .Y(n_348) );
INVx1_ASAP7_75t_L g373 ( .A(n_243), .Y(n_373) );
AND2x2_ASAP7_75t_L g282 ( .A(n_245), .B(n_266), .Y(n_282) );
AND2x2_ASAP7_75t_L g294 ( .A(n_245), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_SL g412 ( .A(n_245), .Y(n_412) );
INVx2_ASAP7_75t_L g302 ( .A(n_246), .Y(n_302) );
AND2x2_ASAP7_75t_L g340 ( .A(n_246), .B(n_256), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_246), .B(n_424), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_253), .B(n_254), .Y(n_248) );
AND2x2_ASAP7_75t_L g355 ( .A(n_249), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g409 ( .A(n_249), .Y(n_409) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g329 ( .A(n_250), .Y(n_329) );
BUFx2_ASAP7_75t_L g428 ( .A(n_250), .Y(n_428) );
BUFx2_ASAP7_75t_L g299 ( .A(n_251), .Y(n_299) );
AND2x2_ASAP7_75t_L g401 ( .A(n_251), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g384 ( .A(n_252), .Y(n_384) );
AND2x4_ASAP7_75t_L g311 ( .A(n_253), .B(n_274), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_253), .B(n_335), .Y(n_347) );
AOI32xp33_ASAP7_75t_L g271 ( .A1(n_254), .A2(n_272), .A3(n_274), .B1(n_276), .B2(n_277), .Y(n_271) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx3_ASAP7_75t_L g260 ( .A(n_255), .Y(n_260) );
OR2x2_ASAP7_75t_L g396 ( .A(n_255), .B(n_352), .Y(n_396) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g265 ( .A(n_256), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g372 ( .A(n_256), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g264 ( .A(n_257), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g276 ( .A(n_257), .B(n_266), .Y(n_276) );
INVx1_ASAP7_75t_L g397 ( .A(n_257), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_257), .B(n_372), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_263), .B(n_267), .C(n_271), .Y(n_258) );
OAI322xp33_ASAP7_75t_L g367 ( .A1(n_259), .A2(n_304), .A3(n_368), .B1(n_370), .B2(n_374), .C1(n_375), .C2(n_379), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVxp67_ASAP7_75t_L g332 ( .A(n_260), .Y(n_332) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g386 ( .A(n_262), .B(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_262), .B(n_302), .Y(n_433) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
OR2x2_ASAP7_75t_L g411 ( .A(n_266), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_269), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g320 ( .A(n_270), .B(n_299), .Y(n_320) );
AND2x2_ASAP7_75t_L g391 ( .A(n_270), .B(n_304), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_270), .B(n_378), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_272), .A2(n_279), .B1(n_282), .B2(n_283), .C(n_288), .Y(n_278) );
OR2x2_ASAP7_75t_L g289 ( .A(n_272), .B(n_285), .Y(n_289) );
AND2x2_ASAP7_75t_L g377 ( .A(n_272), .B(n_378), .Y(n_377) );
AOI32xp33_ASAP7_75t_L g416 ( .A1(n_272), .A2(n_302), .A3(n_417), .B1(n_418), .B2(n_421), .Y(n_416) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND3xp33_ASAP7_75t_L g350 ( .A(n_273), .B(n_309), .C(n_332), .Y(n_350) );
AND2x2_ASAP7_75t_L g376 ( .A(n_273), .B(n_369), .Y(n_376) );
INVxp67_ASAP7_75t_L g356 ( .A(n_274), .Y(n_356) );
BUFx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_277), .B(n_329), .Y(n_385) );
INVx2_ASAP7_75t_L g395 ( .A(n_277), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_277), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g364 ( .A(n_280), .Y(n_364) );
OR2x2_ASAP7_75t_L g290 ( .A(n_281), .B(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_283), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_286), .Y(n_369) );
AND2x2_ASAP7_75t_L g328 ( .A(n_287), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g374 ( .A(n_287), .Y(n_374) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_287), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AOI21xp33_ASAP7_75t_SL g313 ( .A1(n_289), .A2(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g407 ( .A(n_292), .B(n_317), .Y(n_407) );
AOI211xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_296), .B(n_306), .C(n_313), .Y(n_293) );
AND2x2_ASAP7_75t_L g337 ( .A(n_295), .B(n_305), .Y(n_337) );
INVx2_ASAP7_75t_L g352 ( .A(n_295), .Y(n_352) );
OR2x2_ASAP7_75t_L g390 ( .A(n_295), .B(n_353), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_295), .B(n_433), .Y(n_432) );
AOI211xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_298), .B(n_300), .C(n_303), .Y(n_296) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_299), .B(n_337), .Y(n_336) );
OAI211xp5_ASAP7_75t_L g418 ( .A1(n_300), .A2(n_395), .B(n_419), .C(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_301), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g358 ( .A(n_302), .B(n_348), .Y(n_358) );
INVx1_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_307), .B(n_310), .Y(n_306) );
INVxp33_ASAP7_75t_L g414 ( .A(n_308), .Y(n_414) );
AND2x2_ASAP7_75t_L g393 ( .A(n_309), .B(n_372), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_314), .A2(n_376), .B(n_377), .Y(n_375) );
OAI322xp33_ASAP7_75t_L g394 ( .A1(n_316), .A2(n_395), .A3(n_396), .B1(n_397), .B2(n_398), .C1(n_400), .C2(n_404), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B1(n_326), .B2(n_330), .C(n_333), .Y(n_319) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g371 ( .A(n_324), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g415 ( .A(n_328), .Y(n_415) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_331), .B(n_351), .Y(n_417) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g380 ( .A(n_340), .B(n_348), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B1(n_346), .B2(n_348), .C(n_349), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_344), .A2(n_361), .B1(n_365), .B2(n_366), .C(n_367), .Y(n_360) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_348), .B(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_354), .B2(n_357), .Y(n_349) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx2_ASAP7_75t_SL g378 ( .A(n_353), .Y(n_378) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND5xp2_ASAP7_75t_L g359 ( .A(n_360), .B(n_381), .C(n_406), .D(n_416), .E(n_426), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_362), .B(n_364), .Y(n_361) );
NOR4xp25_ASAP7_75t_L g434 ( .A(n_363), .B(n_369), .C(n_435), .D(n_436), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_366), .A2(n_427), .B1(n_429), .B2(n_431), .C(n_434), .Y(n_426) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g425 ( .A(n_372), .Y(n_425) );
OAI322xp33_ASAP7_75t_L g382 ( .A1(n_376), .A2(n_383), .A3(n_384), .B1(n_385), .B2(n_386), .C1(n_388), .C2(n_392), .Y(n_382) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_394), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g427 ( .A(n_402), .B(n_428), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g750 ( .A(n_439), .Y(n_750) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_443), .B(n_687), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_622), .Y(n_443) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_445), .B(n_567), .C(n_591), .D(n_614), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_509), .B1(n_539), .B2(n_551), .C(n_554), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_482), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_448), .A2(n_468), .B1(n_510), .B2(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_448), .B(n_483), .Y(n_625) );
AND2x2_ASAP7_75t_L g644 ( .A(n_448), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_448), .B(n_628), .Y(n_714) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_468), .Y(n_448) );
AND2x2_ASAP7_75t_L g582 ( .A(n_449), .B(n_483), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_449), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g605 ( .A(n_449), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_449), .B(n_469), .Y(n_610) );
INVx2_ASAP7_75t_L g642 ( .A(n_449), .Y(n_642) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_449), .Y(n_686) );
AND2x2_ASAP7_75t_L g703 ( .A(n_449), .B(n_580), .Y(n_703) );
INVx5_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g621 ( .A(n_450), .B(n_580), .Y(n_621) );
AND2x4_ASAP7_75t_L g635 ( .A(n_450), .B(n_468), .Y(n_635) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_450), .Y(n_639) );
AND2x2_ASAP7_75t_L g659 ( .A(n_450), .B(n_574), .Y(n_659) );
AND2x2_ASAP7_75t_L g709 ( .A(n_450), .B(n_484), .Y(n_709) );
AND2x2_ASAP7_75t_L g719 ( .A(n_450), .B(n_469), .Y(n_719) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_465), .Y(n_450) );
AOI21xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_456), .B(n_464), .Y(n_451) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx5_ASAP7_75t_L g474 ( .A(n_457), .Y(n_474) );
INVx2_ASAP7_75t_L g463 ( .A(n_461), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_463), .A2(n_490), .B(n_491), .C(n_492), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_463), .A2(n_492), .B(n_516), .C(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x2_ASAP7_75t_L g575 ( .A(n_468), .B(n_483), .Y(n_575) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_468), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_468), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g665 ( .A(n_468), .Y(n_665) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g553 ( .A(n_469), .B(n_498), .Y(n_553) );
AND2x2_ASAP7_75t_L g580 ( .A(n_469), .B(n_499), .Y(n_580) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_481), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_474), .B(n_475), .C(n_480), .Y(n_472) );
INVx2_ASAP7_75t_L g488 ( .A(n_474), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_474), .A2(n_480), .B(n_525), .C(n_526), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g493 ( .A(n_480), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_482), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_496), .Y(n_482) );
OR2x2_ASAP7_75t_L g606 ( .A(n_483), .B(n_497), .Y(n_606) );
AND2x2_ASAP7_75t_L g643 ( .A(n_483), .B(n_553), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_483), .B(n_574), .Y(n_654) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_483), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_483), .B(n_610), .Y(n_727) );
INVx5_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g552 ( .A(n_484), .Y(n_552) );
AND2x2_ASAP7_75t_L g561 ( .A(n_484), .B(n_497), .Y(n_561) );
AND2x2_ASAP7_75t_L g677 ( .A(n_484), .B(n_572), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_484), .B(n_610), .Y(n_699) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_497), .Y(n_645) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_498), .Y(n_597) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g574 ( .A(n_499), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_510), .B(n_587), .Y(n_706) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_511), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g558 ( .A(n_511), .B(n_559), .Y(n_558) );
INVx5_ASAP7_75t_SL g566 ( .A(n_511), .Y(n_566) );
OR2x2_ASAP7_75t_L g589 ( .A(n_511), .B(n_559), .Y(n_589) );
OR2x2_ASAP7_75t_L g599 ( .A(n_511), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g662 ( .A(n_511), .B(n_521), .Y(n_662) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_511), .B(n_520), .Y(n_700) );
NOR4xp25_ASAP7_75t_L g721 ( .A(n_511), .B(n_642), .C(n_722), .D(n_723), .Y(n_721) );
AND2x2_ASAP7_75t_L g731 ( .A(n_511), .B(n_563), .Y(n_731) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g556 ( .A(n_520), .B(n_552), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_520), .B(n_558), .Y(n_725) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
OR2x2_ASAP7_75t_L g565 ( .A(n_521), .B(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g572 ( .A(n_521), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_521), .B(n_541), .Y(n_584) );
INVxp67_ASAP7_75t_L g587 ( .A(n_521), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_521), .B(n_559), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_521), .B(n_531), .Y(n_653) );
AND2x2_ASAP7_75t_L g668 ( .A(n_521), .B(n_563), .Y(n_668) );
OR2x2_ASAP7_75t_L g697 ( .A(n_521), .B(n_531), .Y(n_697) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_529), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_530), .B(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_530), .B(n_566), .Y(n_705) );
OR2x2_ASAP7_75t_L g726 ( .A(n_530), .B(n_603), .Y(n_726) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g540 ( .A(n_531), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g563 ( .A(n_531), .B(n_559), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_531), .B(n_541), .Y(n_578) );
AND2x2_ASAP7_75t_L g648 ( .A(n_531), .B(n_572), .Y(n_648) );
AND2x2_ASAP7_75t_L g682 ( .A(n_531), .B(n_566), .Y(n_682) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_532), .B(n_566), .Y(n_585) );
AND2x2_ASAP7_75t_L g613 ( .A(n_532), .B(n_541), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_539), .B(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_540), .A2(n_628), .B1(n_664), .B2(n_681), .C(n_683), .Y(n_680) );
INVx5_ASAP7_75t_SL g559 ( .A(n_541), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B(n_545), .Y(n_542) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OAI33xp33_ASAP7_75t_L g579 ( .A1(n_552), .A2(n_580), .A3(n_581), .B1(n_583), .B2(n_586), .B3(n_590), .Y(n_579) );
OR2x2_ASAP7_75t_L g595 ( .A(n_552), .B(n_596), .Y(n_595) );
AOI322xp5_ASAP7_75t_L g704 ( .A1(n_552), .A2(n_621), .A3(n_628), .B1(n_705), .B2(n_706), .C1(n_707), .C2(n_710), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_552), .B(n_580), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_SL g728 ( .A1(n_552), .A2(n_580), .B(n_729), .C(n_731), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_553), .A2(n_568), .B1(n_573), .B2(n_576), .C(n_579), .Y(n_567) );
INVx1_ASAP7_75t_L g660 ( .A(n_553), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_553), .B(n_709), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_557), .B1(n_560), .B2(n_562), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g637 ( .A(n_558), .B(n_572), .Y(n_637) );
AND2x2_ASAP7_75t_L g695 ( .A(n_558), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g603 ( .A(n_559), .B(n_566), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_559), .B(n_572), .Y(n_631) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_561), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_561), .B(n_639), .Y(n_693) );
OAI321xp33_ASAP7_75t_L g712 ( .A1(n_561), .A2(n_634), .A3(n_713), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g679 ( .A(n_562), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_563), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g618 ( .A(n_563), .B(n_566), .Y(n_618) );
AOI321xp33_ASAP7_75t_L g676 ( .A1(n_563), .A2(n_580), .A3(n_677), .B1(n_678), .B2(n_679), .C(n_680), .Y(n_676) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g593 ( .A(n_565), .B(n_578), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_566), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_566), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_566), .B(n_652), .Y(n_689) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g612 ( .A(n_570), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g577 ( .A(n_571), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g685 ( .A(n_572), .Y(n_685) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_575), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g608 ( .A(n_580), .Y(n_608) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_582), .B(n_617), .Y(n_666) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OR2x2_ASAP7_75t_L g630 ( .A(n_585), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g675 ( .A(n_585), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_586), .A2(n_633), .B1(n_636), .B2(n_638), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g730 ( .A(n_589), .B(n_653), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B1(n_598), .B2(n_604), .C(n_607), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g628 ( .A(n_597), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_SL g674 ( .A(n_600), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_602), .B(n_652), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_602), .A2(n_670), .B(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g715 ( .A(n_603), .B(n_697), .Y(n_715) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g617 ( .A(n_606), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B(n_611), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g661 ( .A(n_613), .B(n_662), .Y(n_661) );
INVxp67_ASAP7_75t_L g723 ( .A(n_613), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .B(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_617), .B(n_635), .Y(n_671) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g692 ( .A(n_621), .Y(n_692) );
NAND5xp2_ASAP7_75t_L g622 ( .A(n_623), .B(n_640), .C(n_649), .D(n_669), .E(n_676), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B(n_629), .C(n_632), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g664 ( .A(n_628), .Y(n_664) );
CKINVDCx16_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_636), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g678 ( .A(n_638), .Y(n_678) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_644), .B(n_646), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_641), .A2(n_695), .B1(n_698), .B2(n_700), .C(n_701), .Y(n_694) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AOI321xp33_ASAP7_75t_L g649 ( .A1(n_642), .A2(n_650), .A3(n_654), .B1(n_655), .B2(n_661), .C(n_663), .Y(n_649) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g720 ( .A(n_654), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_656), .B(n_660), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g672 ( .A(n_657), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NOR2xp67_ASAP7_75t_SL g684 ( .A(n_658), .B(n_665), .Y(n_684) );
AOI321xp33_ASAP7_75t_SL g716 ( .A1(n_661), .A2(n_717), .A3(n_718), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_666), .C(n_667), .Y(n_663) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_674), .B(n_682), .Y(n_711) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .C(n_686), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_712), .C(n_724), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_690), .B(n_694), .C(n_704), .Y(n_688) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_692), .B(n_693), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_693), .A2(n_725), .B1(n_726), .B2(n_727), .C(n_728), .Y(n_724) );
INVx1_ASAP7_75t_L g713 ( .A(n_695), .Y(n_713) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g717 ( .A(n_715), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
CKINVDCx14_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx14_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp33_ASAP7_75t_SL g752 ( .A1(n_753), .A2(n_754), .B1(n_760), .B2(n_761), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
BUFx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
INVx5_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx9p33_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
BUFx2_ASAP7_75t_L g777 ( .A(n_770), .Y(n_777) );
OR2x4_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
endmodule