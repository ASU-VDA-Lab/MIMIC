module fake_jpeg_18082_n_163 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_2),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_40),
.B1(n_18),
.B2(n_22),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_16),
.B1(n_17),
.B2(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_18),
.B1(n_22),
.B2(n_20),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_38),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_21),
.B1(n_29),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_55),
.B1(n_30),
.B2(n_28),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_25),
.A3(n_15),
.B1(n_24),
.B2(n_16),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_56),
.Y(n_67)
);

AOI22x1_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_29),
.C(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_62),
.Y(n_86)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_26),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_30),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_11),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_35),
.B1(n_33),
.B2(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_9),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_33),
.B(n_4),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_9),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_6),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_53),
.C(n_10),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_53),
.B1(n_12),
.B2(n_14),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_53),
.C(n_7),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_60),
.C(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_90),
.B1(n_84),
.B2(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_80),
.B(n_74),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_64),
.Y(n_113)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.C(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_119),
.B1(n_72),
.B2(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_83),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_98),
.B(n_97),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_84),
.B1(n_94),
.B2(n_92),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_77),
.B1(n_92),
.B2(n_59),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_86),
.B1(n_87),
.B2(n_101),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_86),
.B1(n_89),
.B2(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_114),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_109),
.C(n_122),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_127),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_119),
.B(n_89),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_107),
.B(n_104),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_137),
.Y(n_148)
);

AO221x1_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_106),
.B1(n_115),
.B2(n_66),
.C(n_58),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AO221x1_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_88),
.B1(n_65),
.B2(n_116),
.C(n_71),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_88),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_126),
.B(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_142),
.B(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_145),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_129),
.B(n_123),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_112),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_138),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_148),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_123),
.A3(n_102),
.B1(n_98),
.B2(n_95),
.C1(n_12),
.C2(n_7),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_158),
.B(n_154),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_157),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_141),
.C(n_149),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_158),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);


endmodule