module fake_jpeg_10781_n_447 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_447);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_447;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_54),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_110),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_56),
.Y(n_117)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_78),
.Y(n_123)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_60),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_14),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_90),
.Y(n_121)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_67),
.B(n_69),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_27),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_12),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_70),
.B(n_99),
.Y(n_133)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_71),
.Y(n_164)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_23),
.B(n_12),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_0),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_21),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_17),
.B(n_41),
.C(n_33),
.Y(n_96)
);

NAND2xp67_ASAP7_75t_SL g181 ( 
.A(n_96),
.B(n_21),
.Y(n_181)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_22),
.B(n_0),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_0),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_51),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_104),
.B(n_109),
.Y(n_174)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_107),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_2),
.C(n_4),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_43),
.B(n_39),
.Y(n_146)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_99),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_28),
.B(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_113),
.Y(n_147)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_56),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_116),
.B(n_135),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_44),
.B1(n_41),
.B2(n_33),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_118),
.A2(n_126),
.B1(n_131),
.B2(n_143),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_61),
.B1(n_109),
.B2(n_104),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_44),
.B1(n_25),
.B2(n_17),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_132),
.B(n_160),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_42),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_42),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_136),
.B(n_137),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_32),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_140),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_73),
.A2(n_25),
.B1(n_51),
.B2(n_28),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_80),
.A2(n_43),
.B1(n_39),
.B2(n_34),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_144),
.A2(n_117),
.B1(n_178),
.B2(n_177),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_49),
.C(n_10),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_65),
.B(n_34),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_165),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_85),
.A2(n_31),
.B1(n_29),
.B2(n_6),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_151),
.A2(n_159),
.B1(n_131),
.B2(n_119),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_98),
.A2(n_31),
.B1(n_29),
.B2(n_7),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_90),
.B(n_4),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_96),
.A2(n_79),
.B(n_21),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_5),
.Y(n_165)
);

INVx2_ASAP7_75t_R g167 ( 
.A(n_100),
.Y(n_167)
);

NAND2x1_ASAP7_75t_SL g228 ( 
.A(n_167),
.B(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_7),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_167),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_101),
.B(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_78),
.B(n_9),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_184),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_78),
.B(n_9),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_67),
.B(n_9),
.C(n_10),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_128),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_147),
.A2(n_49),
.B(n_21),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_187),
.A2(n_204),
.B(n_198),
.Y(n_252)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_188),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_189),
.Y(n_293)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_190),
.Y(n_258)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_194),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_196),
.B(n_205),
.Y(n_260)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_228),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_127),
.A2(n_10),
.B1(n_126),
.B2(n_151),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_199),
.A2(n_243),
.B1(n_189),
.B2(n_215),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_201),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_181),
.A2(n_10),
.B1(n_133),
.B2(n_161),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_202),
.A2(n_221),
.B1(n_223),
.B2(n_232),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_121),
.B(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_206),
.Y(n_282)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_121),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_216),
.Y(n_249)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_211),
.B(n_207),
.Y(n_281)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_213),
.Y(n_253)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_214),
.B(n_217),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_141),
.B(n_153),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_218),
.A2(n_220),
.B1(n_189),
.B2(n_215),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_219),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_125),
.B1(n_155),
.B2(n_170),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_173),
.A2(n_145),
.B1(n_166),
.B2(n_169),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_158),
.B(n_166),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_245),
.C(n_239),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_173),
.A2(n_169),
.B1(n_142),
.B2(n_125),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_225),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_157),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_129),
.B(n_142),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_227),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_154),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_234),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_139),
.A2(n_152),
.B1(n_182),
.B2(n_134),
.Y(n_232)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_154),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_118),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_236),
.Y(n_269)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_238),
.Y(n_273)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_114),
.A2(n_139),
.B1(n_170),
.B2(n_182),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_239),
.A2(n_201),
.B(n_197),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_154),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_242),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_241),
.A2(n_247),
.B1(n_222),
.B2(n_242),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_156),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_159),
.A2(n_123),
.B1(n_172),
.B2(n_120),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_119),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_122),
.B(n_120),
.C(n_168),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_114),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_114),
.A2(n_140),
.B1(n_72),
.B2(n_66),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_168),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_254),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_261),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_203),
.A2(n_172),
.B(n_195),
.C(n_209),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_203),
.A2(n_205),
.B(n_204),
.C(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_264),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_214),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_266),
.A2(n_188),
.B1(n_208),
.B2(n_236),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_193),
.B(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_271),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_270),
.B(n_263),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_193),
.B(n_191),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_194),
.C(n_217),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_278),
.C(n_282),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_222),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_199),
.A2(n_235),
.B1(n_227),
.B2(n_230),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_285),
.B1(n_290),
.B2(n_238),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_271),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_210),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_276),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_250),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_220),
.A2(n_218),
.B1(n_200),
.B2(n_237),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_266),
.A2(n_212),
.B1(n_213),
.B2(n_246),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_298),
.A2(n_300),
.B1(n_304),
.B2(n_315),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_251),
.A2(n_285),
.B1(n_252),
.B2(n_284),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_319),
.B1(n_323),
.B2(n_262),
.Y(n_328)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_270),
.A2(n_226),
.B(n_229),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_303),
.A2(n_324),
.B(n_294),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_224),
.B1(n_244),
.B2(n_292),
.Y(n_304)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

INVx13_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_306),
.B(n_307),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_310),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_289),
.Y(n_310)
);

OR2x2_ASAP7_75t_SL g311 ( 
.A(n_255),
.B(n_254),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_314),
.C(n_308),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_268),
.B(n_249),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_292),
.A2(n_286),
.B1(n_264),
.B2(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_249),
.A2(n_261),
.B1(n_260),
.B2(n_269),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_316),
.A2(n_248),
.B1(n_291),
.B2(n_274),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_273),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_267),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_265),
.B1(n_258),
.B2(n_253),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_327),
.C(n_274),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_265),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_326),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_258),
.A2(n_253),
.B1(n_293),
.B2(n_272),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_257),
.B(n_282),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_267),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_253),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_328),
.A2(n_324),
.B1(n_326),
.B2(n_310),
.Y(n_367)
);

A2O1A1O1Ixp25_ASAP7_75t_L g372 ( 
.A1(n_331),
.A2(n_320),
.B(n_302),
.C(n_309),
.D(n_305),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_332),
.B(n_334),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_263),
.C(n_291),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_343),
.C(n_296),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_325),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_336),
.B(n_340),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_256),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_338),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_275),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_275),
.Y(n_341)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_248),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_298),
.A2(n_287),
.B1(n_300),
.B2(n_299),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_346),
.A2(n_349),
.B1(n_319),
.B2(n_323),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_294),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_348),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_312),
.B1(n_304),
.B2(n_316),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g351 ( 
.A(n_315),
.B(n_308),
.Y(n_351)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_349),
.A2(n_312),
.B(n_324),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_339),
.B(n_345),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_318),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_362),
.C(n_364),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_358),
.A2(n_368),
.B1(n_328),
.B2(n_339),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_327),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_329),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_365),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_347),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_346),
.A2(n_311),
.B1(n_303),
.B2(n_301),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_335),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_369),
.B(n_348),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_296),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_373),
.C(n_333),
.Y(n_389)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_372),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_305),
.C(n_321),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_329),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_375),
.Y(n_382)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_350),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_383),
.Y(n_406)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_359),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_381),
.B(n_388),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_351),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_336),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_389),
.C(n_390),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_386),
.A2(n_366),
.B1(n_363),
.B2(n_361),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_387),
.A2(n_363),
.B(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_337),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_391),
.A2(n_375),
.B(n_365),
.Y(n_399)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_360),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_367),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_373),
.C(n_356),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_396),
.Y(n_411)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_397),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_383),
.C(n_384),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_391),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_366),
.C(n_354),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_407),
.C(n_390),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_376),
.A2(n_358),
.B1(n_368),
.B2(n_344),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_403),
.A2(n_404),
.B1(n_405),
.B2(n_387),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_386),
.A2(n_355),
.B1(n_361),
.B2(n_370),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_391),
.A2(n_355),
.B1(n_370),
.B2(n_338),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_341),
.C(n_340),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_406),
.B(n_379),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_406),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_389),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_410),
.B(n_412),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_415),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_393),
.C(n_335),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_418),
.C(n_398),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g416 ( 
.A(n_401),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_417),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_397),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_408),
.A2(n_403),
.B1(n_378),
.B2(n_382),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_420),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_SL g430 ( 
.A(n_421),
.B(n_409),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_423),
.A2(n_424),
.B(n_425),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_407),
.C(n_400),
.Y(n_424)
);

O2A1O1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_415),
.A2(n_399),
.B(n_396),
.C(n_394),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_R g428 ( 
.A(n_426),
.B(n_334),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_429),
.Y(n_435)
);

AOI21x1_ASAP7_75t_L g429 ( 
.A1(n_425),
.A2(n_347),
.B(n_402),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_433),
.B(n_421),
.Y(n_434)
);

INVx13_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_422),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_372),
.B(n_404),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_437),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_427),
.A2(n_423),
.B(n_419),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_436),
.B(n_438),
.C(n_422),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_342),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_439),
.A2(n_381),
.B1(n_353),
.B2(n_342),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_411),
.C(n_432),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_440),
.B(n_411),
.Y(n_442)
);

BUFx24_ASAP7_75t_SL g444 ( 
.A(n_442),
.Y(n_444)
);

AOI322xp5_ASAP7_75t_L g445 ( 
.A1(n_444),
.A2(n_443),
.A3(n_441),
.B1(n_330),
.B2(n_385),
.C1(n_405),
.C2(n_353),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_352),
.B(n_332),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);


endmodule