module fake_jpeg_6616_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_9),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_2),
.C(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_19),
.B1(n_18),
.B2(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_18),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_26),
.B1(n_24),
.B2(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_44),
.B1(n_37),
.B2(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_31),
.B1(n_13),
.B2(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_28),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_39),
.B1(n_42),
.B2(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_38),
.C(n_45),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_55),
.C(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_64),
.B1(n_62),
.B2(n_67),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_64),
.B(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2x1_ASAP7_75t_R g65 ( 
.A(n_52),
.B(n_27),
.Y(n_65)
);

OA21x2_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_36),
.B(n_53),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_48),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_70),
.C(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_54),
.B1(n_55),
.B2(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_73),
.B(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_75),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_54),
.A3(n_44),
.B1(n_51),
.B2(n_13),
.C(n_16),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_62),
.B(n_58),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_51),
.C(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_20),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_14),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_84),
.C(n_14),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_86),
.B1(n_14),
.B2(n_3),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_70),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_75),
.B1(n_68),
.B2(n_8),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_79),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_92),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_14),
.Y(n_92)
);

XNOR2x1_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_2),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_81),
.B(n_87),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g96 ( 
.A(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_98),
.B1(n_89),
.B2(n_4),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_79),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_101),
.C(n_6),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_80),
.B(n_82),
.C(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_104)
);

OAI211xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_105),
.B(n_6),
.C(n_7),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_107),
.B1(n_104),
.B2(n_102),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_7),
.Y(n_110)
);


endmodule