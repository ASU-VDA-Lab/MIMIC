module real_jpeg_28968_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_285, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_285;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_0),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_4),
.B1(n_18),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_23),
.B(n_25),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_35),
.B1(n_41),
.B2(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_3),
.B(n_24),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_5),
.B(n_41),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_3),
.A2(n_58),
.B(n_62),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_40),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_4),
.A2(n_9),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_4),
.A2(n_10),
.B1(n_18),
.B2(n_28),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_8),
.B1(n_18),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_4),
.A2(n_22),
.B(n_35),
.C(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_42),
.Y(n_45)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_50),
.B1(n_61),
.B2(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_41),
.B1(n_43),
.B2(n_50),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_9),
.A2(n_19),
.B1(n_61),
.B2(n_62),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_9),
.A2(n_19),
.B1(n_41),
.B2(n_43),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_28),
.B1(n_41),
.B2(n_43),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_10),
.A2(n_28),
.B1(n_61),
.B2(n_62),
.Y(n_200)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_11),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_277),
.B(n_281),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_65),
.B(n_276),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_29),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_15),
.B(n_29),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_15),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_24),
.B2(n_27),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_32),
.B(n_33),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_20),
.A2(n_24),
.B1(n_34),
.B2(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_20),
.B(n_24),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_SL g26 ( 
.A(n_25),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_25),
.A2(n_35),
.B(n_138),
.C(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_27),
.B(n_280),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_30),
.B(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_30),
.B(n_274),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_36),
.CI(n_46),
.CON(n_30),
.SN(n_30)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_32),
.A2(n_33),
.B(n_49),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_34),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_35),
.A2(n_41),
.B(n_59),
.C(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_35),
.B(n_92),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_35),
.B(n_60),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_40),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_39),
.B(n_77),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_40),
.A2(n_52),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_44),
.B(n_78),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.C(n_53),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_47),
.B(n_81),
.C(n_82),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_47),
.A2(n_80),
.B1(n_96),
.B2(n_121),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_47),
.B(n_121),
.C(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_47),
.A2(n_80),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_51),
.A2(n_53),
.B1(n_255),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_53),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_53),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_56),
.A2(n_60),
.B1(n_101),
.B2(n_108),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_56),
.A2(n_60),
.B1(n_64),
.B2(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_60),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_61),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_89),
.Y(n_88)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_273),
.B(n_275),
.Y(n_65)
);

OAI321xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_247),
.A3(n_266),
.B1(n_271),
.B2(n_272),
.C(n_285),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_229),
.B(n_246),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_210),
.B(n_228),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_131),
.B(n_193),
.C(n_209),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_118),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_71),
.B(n_118),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_93),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_72),
.B(n_94),
.C(n_104),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_82),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_128),
.C(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_74),
.A2(n_81),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_74),
.A2(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_74),
.B(n_235),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_79),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_86),
.A2(n_126),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_86),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_86),
.B(n_176),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_86),
.B(n_153),
.C(n_165),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_89),
.B(n_115),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_88),
.B(n_89),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_88),
.A2(n_92),
.B1(n_113),
.B2(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_103),
.B2(n_104),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_102),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_96),
.A2(n_105),
.B1(n_106),
.B2(n_121),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_97),
.Y(n_254)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_102),
.A2(n_122),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_102),
.A2(n_122),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_102),
.A2(n_122),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_102),
.B(n_253),
.C(n_255),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_102),
.B(n_260),
.C(n_265),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_111),
.B2(n_112),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_105),
.A2(n_106),
.B1(n_160),
.B2(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_105),
.B(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_121),
.C(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_106),
.B(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B(n_110),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.C(n_127),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_119),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_122),
.B(n_203),
.C(n_205),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_127),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_192),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_186),
.B(n_191),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_156),
.B(n_185),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_144),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_153),
.C(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_147),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_152),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_155),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_155),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_153),
.B(n_199),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_180),
.B(n_184),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_167),
.B(n_179),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_162),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_164),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_171),
.B(n_178),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_175),
.B(n_177),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_194),
.B(n_195),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_207),
.B2(n_208),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_202),
.C(n_208),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_207),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_211),
.B(n_212),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_227),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_219),
.C(n_227),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_224),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_224),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_238),
.B(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_244),
.B2(n_245),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_237),
.C(n_245),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_249),
.C(n_256),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_249),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_258),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_257),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_265),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);


endmodule