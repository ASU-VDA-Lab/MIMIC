module real_aes_15465_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_1280;
wire n_394;
wire n_729;
wire n_1323;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1303 ( .A1(n_0), .A2(n_7), .B1(n_1246), .B2(n_1304), .Y(n_1303) );
AOI22xp33_ASAP7_75t_SL g1336 ( .A1(n_0), .A2(n_217), .B1(n_605), .B2(n_1337), .Y(n_1336) );
OAI22xp33_ASAP7_75t_SL g385 ( .A1(n_1), .A2(n_116), .B1(n_386), .B2(n_389), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_1), .A2(n_25), .B1(n_422), .B2(n_423), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_2), .A2(n_26), .B1(n_380), .B2(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_SL g480 ( .A1(n_2), .A2(n_118), .B1(n_401), .B2(n_422), .Y(n_480) );
INVx1_ASAP7_75t_L g608 ( .A(n_3), .Y(n_608) );
INVx1_ASAP7_75t_L g978 ( .A(n_4), .Y(n_978) );
INVx1_ASAP7_75t_L g1206 ( .A(n_5), .Y(n_1206) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_6), .A2(n_232), .B1(n_532), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_6), .A2(n_166), .B1(n_681), .B2(n_683), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_7), .A2(n_225), .B1(n_739), .B2(n_1337), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_8), .Y(n_471) );
INVx1_ASAP7_75t_L g868 ( .A(n_9), .Y(n_868) );
AOI22xp5_ASAP7_75t_SL g1035 ( .A1(n_10), .A2(n_233), .B1(n_1019), .B2(n_1021), .Y(n_1035) );
INVx1_ASAP7_75t_L g589 ( .A(n_11), .Y(n_589) );
AOI21xp33_ASAP7_75t_L g1226 ( .A1(n_12), .A2(n_304), .B(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1276 ( .A(n_12), .Y(n_1276) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_13), .A2(n_214), .B1(n_532), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_13), .A2(n_198), .B1(n_685), .B2(n_686), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_14), .Y(n_436) );
INVx1_ASAP7_75t_L g259 ( .A(n_15), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_15), .B(n_269), .Y(n_334) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_15), .B(n_204), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_15), .B(n_388), .Y(n_1245) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_16), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_17), .A2(n_207), .B1(n_528), .B2(n_532), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_17), .A2(n_61), .B1(n_556), .B2(n_559), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_18), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_19), .Y(n_312) );
INVx1_ASAP7_75t_L g1318 ( .A(n_20), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1328 ( .A1(n_20), .A2(n_40), .B1(n_482), .B2(n_542), .Y(n_1328) );
OAI222xp33_ASAP7_75t_L g496 ( .A1(n_21), .A2(n_193), .B1(n_375), .B2(n_381), .C1(n_497), .C2(n_499), .Y(n_496) );
OAI222xp33_ASAP7_75t_L g539 ( .A1(n_21), .A2(n_133), .B1(n_193), .B2(n_540), .C1(n_542), .C2(n_543), .Y(n_539) );
OAI211xp5_ASAP7_75t_L g884 ( .A1(n_22), .A2(n_794), .B(n_885), .C(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g897 ( .A(n_22), .Y(n_897) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_23), .B(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_L g1017 ( .A(n_23), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_23), .B(n_104), .Y(n_1022) );
INVx1_ASAP7_75t_L g1323 ( .A(n_24), .Y(n_1323) );
OAI22xp33_ASAP7_75t_SL g379 ( .A1(n_25), .A2(n_218), .B1(n_380), .B2(n_382), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_26), .B(n_399), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_27), .A2(n_197), .B1(n_422), .B2(n_610), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_27), .A2(n_245), .B1(n_380), .B2(n_477), .Y(n_622) );
AOI22xp5_ASAP7_75t_SL g1027 ( .A1(n_28), .A2(n_124), .B1(n_1019), .B2(n_1021), .Y(n_1027) );
INVx1_ASAP7_75t_L g905 ( .A(n_29), .Y(n_905) );
INVx1_ASAP7_75t_L g865 ( .A(n_30), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g826 ( .A1(n_31), .A2(n_146), .B1(n_389), .B2(n_476), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g828 ( .A1(n_31), .A2(n_241), .B1(n_422), .B2(n_423), .Y(n_828) );
INVx1_ASAP7_75t_L g514 ( .A(n_32), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_32), .A2(n_207), .B1(n_559), .B2(n_573), .Y(n_572) );
XOR2xp5_ASAP7_75t_L g275 ( .A(n_33), .B(n_276), .Y(n_275) );
AOI22xp5_ASAP7_75t_SL g1039 ( .A1(n_34), .A2(n_228), .B1(n_1002), .B2(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1219 ( .A(n_35), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_35), .A2(n_130), .B1(n_1266), .B2(n_1267), .Y(n_1265) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_36), .Y(n_808) );
XNOR2x2_ASAP7_75t_SL g878 ( .A(n_37), .B(n_879), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g845 ( .A1(n_38), .A2(n_128), .B1(n_380), .B2(n_477), .Y(n_845) );
OAI22xp33_ASAP7_75t_SL g847 ( .A1(n_38), .A2(n_128), .B1(n_422), .B2(n_848), .Y(n_847) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_39), .Y(n_452) );
INVx1_ASAP7_75t_L g1321 ( .A(n_40), .Y(n_1321) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_41), .A2(n_187), .B1(n_380), .B2(n_786), .Y(n_785) );
OAI22xp33_ASAP7_75t_L g789 ( .A1(n_41), .A2(n_98), .B1(n_422), .B2(n_423), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_42), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_43), .Y(n_320) );
INVx1_ASAP7_75t_L g889 ( .A(n_44), .Y(n_889) );
OAI211xp5_ASAP7_75t_L g893 ( .A1(n_44), .A2(n_461), .B(n_894), .C(n_896), .Y(n_893) );
INVx1_ASAP7_75t_L g694 ( .A(n_45), .Y(n_694) );
INVx1_ASAP7_75t_L g968 ( .A(n_46), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g1058 ( .A1(n_47), .A2(n_160), .B1(n_1002), .B2(n_1015), .Y(n_1058) );
INVx1_ASAP7_75t_L g1324 ( .A(n_48), .Y(n_1324) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_49), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_50), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_51), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_52), .A2(n_103), .B1(n_1019), .B2(n_1045), .Y(n_1080) );
AOI22xp5_ASAP7_75t_L g1030 ( .A1(n_53), .A2(n_88), .B1(n_1015), .B2(n_1019), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1059 ( .A1(n_54), .A2(n_162), .B1(n_1019), .B2(n_1040), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_55), .A2(n_136), .B1(n_542), .B2(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_55), .Y(n_712) );
INVx1_ASAP7_75t_L g633 ( .A(n_56), .Y(n_633) );
INVx1_ASAP7_75t_L g843 ( .A(n_57), .Y(n_843) );
OAI211xp5_ASAP7_75t_SL g1193 ( .A1(n_58), .A2(n_1194), .B(n_1199), .C(n_1208), .Y(n_1193) );
INVx1_ASAP7_75t_L g1248 ( .A(n_58), .Y(n_1248) );
INVx1_ASAP7_75t_L g293 ( .A(n_59), .Y(n_293) );
INVx1_ASAP7_75t_L g299 ( .A(n_59), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_60), .A2(n_123), .B1(n_935), .B2(n_937), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_60), .A2(n_123), .B1(n_261), .B2(n_389), .Y(n_961) );
INVx1_ASAP7_75t_L g518 ( .A(n_61), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_62), .Y(n_439) );
XOR2xp5_ASAP7_75t_L g575 ( .A(n_63), .B(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_63), .A2(n_244), .B1(n_1002), .B2(n_1015), .Y(n_1014) );
XOR2x2_ASAP7_75t_L g690 ( .A(n_64), .B(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_65), .A2(n_78), .B1(n_532), .B2(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_65), .A2(n_223), .B1(n_739), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_66), .A2(n_77), .B1(n_1304), .B2(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1335 ( .A(n_66), .Y(n_1335) );
OAI211xp5_ASAP7_75t_L g780 ( .A1(n_67), .A2(n_362), .B(n_781), .C(n_782), .Y(n_780) );
INVx1_ASAP7_75t_L g796 ( .A(n_67), .Y(n_796) );
INVx1_ASAP7_75t_L g253 ( .A(n_68), .Y(n_253) );
INVx2_ASAP7_75t_L g286 ( .A(n_69), .Y(n_286) );
INVx1_ASAP7_75t_L g581 ( .A(n_70), .Y(n_581) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_71), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_71), .A2(n_136), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_72), .A2(n_74), .B1(n_1015), .B2(n_1019), .Y(n_1041) );
INVx1_ASAP7_75t_L g914 ( .A(n_73), .Y(n_914) );
INVx1_ASAP7_75t_L g1314 ( .A(n_75), .Y(n_1314) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_76), .A2(n_98), .B1(n_386), .B2(n_389), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_76), .A2(n_187), .B1(n_399), .B2(n_401), .Y(n_797) );
INVxp67_ASAP7_75t_SL g1339 ( .A(n_77), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_78), .A2(n_86), .B1(n_685), .B2(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g861 ( .A(n_79), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_80), .Y(n_761) );
XOR2xp5_ASAP7_75t_L g487 ( .A(n_81), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g842 ( .A(n_82), .Y(n_842) );
INVx1_ASAP7_75t_L g369 ( .A(n_83), .Y(n_369) );
OAI211xp5_ASAP7_75t_SL g402 ( .A1(n_83), .A2(n_403), .B(n_408), .C(n_418), .Y(n_402) );
INVx1_ASAP7_75t_L g639 ( .A(n_84), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_84), .A2(n_222), .B1(n_295), .B2(n_646), .C(n_648), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_85), .A2(n_144), .B1(n_468), .B2(n_476), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_85), .A2(n_144), .B1(n_399), .B2(n_401), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_86), .A2(n_223), .B1(n_523), .B2(n_725), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_87), .A2(n_170), .B1(n_1002), .B2(n_1021), .Y(n_1029) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_88), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1230 ( .A(n_89), .Y(n_1230) );
INVx1_ASAP7_75t_L g1319 ( .A(n_90), .Y(n_1319) );
AOI221xp5_ASAP7_75t_L g1220 ( .A1(n_91), .A2(n_127), .B1(n_686), .B2(n_745), .C(n_1221), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_91), .A2(n_183), .B1(n_1266), .B2(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g750 ( .A(n_92), .Y(n_750) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_93), .A2(n_245), .B1(n_399), .B2(n_423), .C(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g620 ( .A(n_93), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_94), .A2(n_156), .B1(n_468), .B2(n_476), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g854 ( .A1(n_94), .A2(n_156), .B1(n_399), .B2(n_401), .Y(n_854) );
INVx1_ASAP7_75t_L g974 ( .A(n_95), .Y(n_974) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_96), .Y(n_255) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_96), .B(n_253), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g490 ( .A1(n_97), .A2(n_491), .B(n_492), .C(n_503), .Y(n_490) );
INVx1_ASAP7_75t_L g547 ( .A(n_97), .Y(n_547) );
INVx1_ASAP7_75t_L g583 ( .A(n_99), .Y(n_583) );
INVx1_ASAP7_75t_L g912 ( .A(n_100), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_101), .A2(n_198), .B1(n_494), .B2(n_660), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_101), .A2(n_214), .B1(n_671), .B2(n_673), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_102), .A2(n_145), .B1(n_1002), .B2(n_1015), .Y(n_1043) );
INVx1_ASAP7_75t_L g1005 ( .A(n_104), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_104), .B(n_1017), .Y(n_1020) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_105), .A2(n_167), .B1(n_1002), .B2(n_1015), .Y(n_1036) );
INVx1_ASAP7_75t_L g584 ( .A(n_106), .Y(n_584) );
INVx1_ASAP7_75t_L g702 ( .A(n_107), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_108), .Y(n_810) );
INVx2_ASAP7_75t_L g285 ( .A(n_109), .Y(n_285) );
INVx1_ASAP7_75t_L g329 ( .A(n_109), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_109), .B(n_286), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_110), .Y(n_756) );
INVx1_ASAP7_75t_L g908 ( .A(n_111), .Y(n_908) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_112), .A2(n_234), .B1(n_532), .B2(n_727), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_112), .A2(n_172), .B1(n_554), .B2(n_737), .Y(n_741) );
INVxp67_ASAP7_75t_SL g1224 ( .A(n_113), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_113), .A2(n_127), .B1(n_710), .B2(n_722), .Y(n_1262) );
INVx1_ASAP7_75t_L g859 ( .A(n_114), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_115), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_116), .A2(n_218), .B1(n_399), .B2(n_401), .Y(n_398) );
OAI22xp33_ASAP7_75t_SL g475 ( .A1(n_117), .A2(n_118), .B1(n_476), .B2(n_477), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_117), .A2(n_121), .B1(n_413), .B2(n_414), .Y(n_484) );
INVx1_ASAP7_75t_L g983 ( .A(n_119), .Y(n_983) );
INVx1_ASAP7_75t_L g867 ( .A(n_120), .Y(n_867) );
INVx1_ASAP7_75t_L g473 ( .A(n_121), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_122), .A2(n_211), .B1(n_422), .B2(n_891), .Y(n_890) );
OAI22xp33_ASAP7_75t_L g901 ( .A1(n_122), .A2(n_211), .B1(n_380), .B2(n_389), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_125), .Y(n_823) );
INVx1_ASAP7_75t_L g1079 ( .A(n_126), .Y(n_1079) );
AOI222xp33_ASAP7_75t_L g1187 ( .A1(n_126), .A2(n_1188), .B1(n_1290), .B2(n_1294), .C1(n_1343), .C2(n_1345), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_126), .A2(n_1079), .B1(n_1191), .B2(n_1289), .Y(n_1190) );
INVx1_ASAP7_75t_L g920 ( .A(n_129), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g1228 ( .A1(n_130), .A2(n_183), .B1(n_671), .B2(n_737), .Y(n_1228) );
INVx1_ASAP7_75t_L g502 ( .A(n_131), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_131), .A2(n_203), .B1(n_399), .B2(n_401), .Y(n_544) );
INVx1_ASAP7_75t_L g1210 ( .A(n_132), .Y(n_1210) );
OAI221xp5_ASAP7_75t_L g1252 ( .A1(n_132), .A2(n_185), .B1(n_1253), .B2(n_1259), .C(n_1261), .Y(n_1252) );
INVx1_ASAP7_75t_L g493 ( .A(n_133), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_134), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_135), .A2(n_165), .B1(n_1019), .B2(n_1045), .Y(n_1044) );
BUFx3_ASAP7_75t_L g291 ( .A(n_137), .Y(n_291) );
OAI211xp5_ASAP7_75t_SL g469 ( .A1(n_138), .A2(n_361), .B(n_362), .C(n_470), .Y(n_469) );
OAI211xp5_ASAP7_75t_SL g481 ( .A1(n_138), .A2(n_418), .B(n_482), .C(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g1212 ( .A(n_139), .Y(n_1212) );
INVx1_ASAP7_75t_L g1302 ( .A(n_140), .Y(n_1302) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_141), .Y(n_768) );
INVx1_ASAP7_75t_L g966 ( .A(n_142), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_143), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_146), .A2(n_246), .B1(n_399), .B2(n_401), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_147), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_148), .A2(n_195), .B1(n_1019), .B2(n_1021), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_149), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_150), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_151), .Y(n_509) );
INVx1_ASAP7_75t_L g607 ( .A(n_152), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_153), .Y(n_803) );
XOR2xp5_ASAP7_75t_L g1295 ( .A(n_154), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g971 ( .A(n_155), .Y(n_971) );
INVx1_ASAP7_75t_L g917 ( .A(n_157), .Y(n_917) );
INVx1_ASAP7_75t_L g943 ( .A(n_158), .Y(n_943) );
INVx1_ASAP7_75t_L g921 ( .A(n_159), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_161), .Y(n_302) );
INVx1_ASAP7_75t_L g1315 ( .A(n_163), .Y(n_1315) );
INVx1_ASAP7_75t_L g592 ( .A(n_164), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_166), .A2(n_226), .B1(n_660), .B2(n_662), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_168), .A2(n_181), .B1(n_399), .B2(n_882), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_168), .A2(n_181), .B1(n_386), .B2(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g507 ( .A(n_169), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_169), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g695 ( .A(n_171), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_172), .A2(n_179), .B1(n_722), .B2(n_725), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_173), .B(n_406), .Y(n_606) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_173), .Y(n_615) );
OAI211xp5_ASAP7_75t_SL g938 ( .A1(n_174), .A2(n_418), .B(n_939), .C(n_940), .Y(n_938) );
INVx1_ASAP7_75t_L g956 ( .A(n_174), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_175), .Y(n_324) );
INVx1_ASAP7_75t_L g632 ( .A(n_176), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_177), .Y(n_807) );
OAI211xp5_ASAP7_75t_L g360 ( .A1(n_178), .A2(n_361), .B(n_362), .C(n_368), .Y(n_360) );
INVx1_ASAP7_75t_L g417 ( .A(n_178), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_179), .A2(n_234), .B1(n_554), .B2(n_737), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_180), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_182), .A2(n_238), .B1(n_882), .B2(n_947), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_182), .A2(n_238), .B1(n_958), .B2(n_959), .Y(n_957) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
INVx1_ASAP7_75t_L g1233 ( .A(n_185), .Y(n_1233) );
INVx1_ASAP7_75t_L g638 ( .A(n_186), .Y(n_638) );
INVx1_ASAP7_75t_L g824 ( .A(n_188), .Y(n_824) );
OAI211xp5_ASAP7_75t_L g829 ( .A1(n_188), .A2(n_791), .B(n_794), .C(n_830), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_189), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_190), .Y(n_755) );
INVx1_ASAP7_75t_L g918 ( .A(n_191), .Y(n_918) );
INVx1_ASAP7_75t_L g587 ( .A(n_192), .Y(n_587) );
INVx1_ASAP7_75t_L g864 ( .A(n_194), .Y(n_864) );
OA22x2_ASAP7_75t_L g628 ( .A1(n_196), .A2(n_629), .B1(n_688), .B2(n_689), .Y(n_628) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_196), .Y(n_689) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_197), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_199), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_200), .Y(n_453) );
XOR2xp5_ASAP7_75t_L g431 ( .A(n_201), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g862 ( .A(n_202), .Y(n_862) );
INVx1_ASAP7_75t_L g504 ( .A(n_203), .Y(n_504) );
BUFx3_ASAP7_75t_L g269 ( .A(n_204), .Y(n_269) );
INVx1_ASAP7_75t_L g388 ( .A(n_204), .Y(n_388) );
XOR2x2_ASAP7_75t_L g931 ( .A(n_205), .B(n_932), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_206), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_208), .Y(n_441) );
INVx1_ASAP7_75t_L g580 ( .A(n_209), .Y(n_580) );
OAI211xp5_ASAP7_75t_L g821 ( .A1(n_210), .A2(n_362), .B(n_781), .C(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g831 ( .A(n_210), .Y(n_831) );
INVx1_ASAP7_75t_L g1200 ( .A(n_212), .Y(n_1200) );
INVx1_ASAP7_75t_L g858 ( .A(n_213), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_215), .Y(n_764) );
INVx1_ASAP7_75t_L g980 ( .A(n_216), .Y(n_980) );
INVxp67_ASAP7_75t_SL g1307 ( .A(n_217), .Y(n_1307) );
OAI211xp5_ASAP7_75t_L g839 ( .A1(n_219), .A2(n_362), .B(n_840), .C(n_841), .Y(n_839) );
INVx1_ASAP7_75t_L g851 ( .A(n_219), .Y(n_851) );
INVx1_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
INVx2_ASAP7_75t_L g327 ( .A(n_220), .Y(n_327) );
INVx1_ASAP7_75t_L g567 ( .A(n_220), .Y(n_567) );
INVx1_ASAP7_75t_L g888 ( .A(n_221), .Y(n_888) );
OAI211xp5_ASAP7_75t_L g635 ( .A1(n_222), .A2(n_513), .B(n_636), .C(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g1301 ( .A(n_224), .Y(n_1301) );
INVxp67_ASAP7_75t_SL g1308 ( .A(n_225), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_226), .A2(n_232), .B1(n_676), .B2(n_678), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g1026 ( .A1(n_227), .A2(n_240), .B1(n_1002), .B2(n_1015), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_229), .Y(n_316) );
INVx1_ASAP7_75t_L g1078 ( .A(n_230), .Y(n_1078) );
INVx1_ASAP7_75t_L g591 ( .A(n_231), .Y(n_591) );
INVx1_ASAP7_75t_L g1218 ( .A(n_235), .Y(n_1218) );
INVx1_ASAP7_75t_L g704 ( .A(n_236), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g522 ( .A1(n_237), .A2(n_523), .B(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g552 ( .A(n_237), .Y(n_552) );
INVx1_ASAP7_75t_L g982 ( .A(n_239), .Y(n_982) );
XNOR2xp5_ASAP7_75t_L g798 ( .A(n_240), .B(n_799), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_241), .A2(n_246), .B1(n_380), .B2(n_786), .Y(n_825) );
INVx1_ASAP7_75t_L g945 ( .A(n_242), .Y(n_945) );
OAI211xp5_ASAP7_75t_L g950 ( .A1(n_242), .A2(n_951), .B(n_953), .C(n_954), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g769 ( .A(n_243), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_247), .Y(n_500) );
INVx1_ASAP7_75t_L g784 ( .A(n_248), .Y(n_784) );
OAI211xp5_ASAP7_75t_L g790 ( .A1(n_248), .A2(n_791), .B(n_794), .C(n_795), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_998), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g1293 ( .A(n_251), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_252), .B(n_255), .Y(n_1344) );
INVx1_ASAP7_75t_L g1349 ( .A(n_252), .Y(n_1349) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1351 ( .A(n_255), .B(n_1349), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g394 ( .A(n_258), .B(n_395), .Y(n_394) );
AOI21xp5_ASAP7_75t_SL g489 ( .A1(n_258), .A2(n_490), .B(n_505), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_258), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g358 ( .A(n_259), .B(n_269), .Y(n_358) );
AND2x4_ASAP7_75t_L g526 ( .A(n_259), .B(n_268), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_260), .A2(n_390), .B1(n_632), .B2(n_633), .Y(n_631) );
AND2x4_ASAP7_75t_SL g1291 ( .A(n_260), .B(n_1292), .Y(n_1291) );
AOI22xp33_ASAP7_75t_SL g1322 ( .A1(n_260), .A2(n_390), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
INVx1_ASAP7_75t_L g355 ( .A(n_262), .Y(n_355) );
OR2x6_ASAP7_75t_L g386 ( .A(n_262), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g476 ( .A(n_262), .B(n_387), .Y(n_476) );
BUFx4f_ASAP7_75t_L g508 ( .A(n_262), .Y(n_508) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx4f_ASAP7_75t_L g337 ( .A(n_263), .Y(n_337) );
INVx3_ASAP7_75t_L g381 ( .A(n_263), .Y(n_381) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g342 ( .A(n_265), .Y(n_342) );
INVx2_ASAP7_75t_L g347 ( .A(n_265), .Y(n_347) );
NAND2x1_ASAP7_75t_L g351 ( .A(n_265), .B(n_266), .Y(n_351) );
AND2x2_ASAP7_75t_L g367 ( .A(n_265), .B(n_266), .Y(n_367) );
INVx1_ASAP7_75t_L g378 ( .A(n_265), .Y(n_378) );
AND2x2_ASAP7_75t_L g391 ( .A(n_265), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_266), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g346 ( .A(n_266), .B(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g372 ( .A(n_266), .Y(n_372) );
INVx2_ASAP7_75t_L g392 ( .A(n_266), .Y(n_392) );
INVx1_ASAP7_75t_L g531 ( .A(n_266), .Y(n_531) );
AND2x2_ASAP7_75t_L g533 ( .A(n_266), .B(n_342), .Y(n_533) );
OR2x6_ASAP7_75t_L g380 ( .A(n_267), .B(n_381), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_267), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g364 ( .A(n_268), .Y(n_364) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g371 ( .A(n_269), .Y(n_371) );
AND2x4_ASAP7_75t_L g376 ( .A(n_269), .B(n_377), .Y(n_376) );
XNOR2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_623), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
XNOR2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_486), .Y(n_273) );
XNOR2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_431), .Y(n_274) );
NAND3xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_359), .C(n_397), .Y(n_276) );
NOR2xp33_ASAP7_75t_SL g277 ( .A(n_278), .B(n_331), .Y(n_277) );
OAI33xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_287), .A3(n_301), .B1(n_313), .B2(n_321), .B3(n_325), .Y(n_278) );
OAI33xp33_ASAP7_75t_L g434 ( .A1(n_279), .A2(n_325), .A3(n_435), .B1(n_440), .B2(n_446), .B3(n_451), .Y(n_434) );
OAI33xp33_ASAP7_75t_L g753 ( .A1(n_279), .A2(n_325), .A3(n_754), .B1(n_757), .B2(n_760), .B3(n_765), .Y(n_753) );
OAI33xp33_ASAP7_75t_L g815 ( .A1(n_279), .A2(n_325), .A3(n_816), .B1(n_817), .B2(n_818), .B3(n_819), .Y(n_815) );
OAI33xp33_ASAP7_75t_L g856 ( .A1(n_279), .A2(n_325), .A3(n_857), .B1(n_860), .B2(n_863), .B3(n_866), .Y(n_856) );
BUFx4f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g550 ( .A(n_280), .Y(n_550) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_281), .B(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_281), .Y(n_430) );
INVx1_ASAP7_75t_L g733 ( .A(n_281), .Y(n_733) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g396 ( .A(n_282), .Y(n_396) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g1227 ( .A(n_284), .Y(n_1227) );
NAND2xp33_ASAP7_75t_SL g284 ( .A(n_285), .B(n_286), .Y(n_284) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_285), .Y(n_428) );
AND3x4_ASAP7_75t_L g668 ( .A(n_285), .B(n_406), .C(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g1198 ( .A(n_285), .Y(n_1198) );
INVx3_ASAP7_75t_L g330 ( .A(n_286), .Y(n_330) );
BUFx3_ASAP7_75t_L g406 ( .A(n_286), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B1(n_294), .B2(n_295), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_288), .A2(n_322), .B1(n_336), .B2(n_338), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g321 ( .A1(n_289), .A2(n_322), .B1(n_323), .B2(n_324), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_289), .A2(n_436), .B1(n_437), .B2(n_439), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_289), .A2(n_323), .B1(n_452), .B2(n_453), .Y(n_451) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_289), .A2(n_540), .B1(n_580), .B2(n_581), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_289), .A2(n_295), .B1(n_591), .B2(n_592), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_289), .A2(n_437), .B1(n_755), .B2(n_756), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_289), .A2(n_295), .B1(n_858), .B2(n_859), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g866 ( .A1(n_289), .A2(n_323), .B1(n_867), .B2(n_868), .Y(n_866) );
BUFx4f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x4_ASAP7_75t_L g399 ( .A(n_290), .B(n_400), .Y(n_399) );
OR2x4_ASAP7_75t_L g422 ( .A(n_290), .B(n_330), .Y(n_422) );
INVx2_ASAP7_75t_L g767 ( .A(n_290), .Y(n_767) );
BUFx3_ASAP7_75t_L g967 ( .A(n_290), .Y(n_967) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_291), .Y(n_300) );
INVx2_ASAP7_75t_L g307 ( .A(n_291), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_291), .B(n_299), .Y(n_311) );
AND2x4_ASAP7_75t_L g420 ( .A(n_291), .B(n_412), .Y(n_420) );
INVx1_ASAP7_75t_L g558 ( .A(n_292), .Y(n_558) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVxp67_ASAP7_75t_L g306 ( .A(n_293), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_294), .A2(n_324), .B1(n_344), .B2(n_348), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g816 ( .A1(n_295), .A2(n_766), .B1(n_803), .B2(n_810), .Y(n_816) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx3_ASAP7_75t_L g438 ( .A(n_296), .Y(n_438) );
INVx4_ASAP7_75t_L g541 ( .A(n_296), .Y(n_541) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
BUFx2_ASAP7_75t_L g793 ( .A(n_297), .Y(n_793) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
BUFx2_ASAP7_75t_L g416 ( .A(n_298), .Y(n_416) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g412 ( .A(n_299), .Y(n_412) );
BUFx2_ASAP7_75t_L g407 ( .A(n_300), .Y(n_407) );
INVx2_ASAP7_75t_L g414 ( .A(n_300), .Y(n_414) );
AND2x4_ASAP7_75t_L g562 ( .A(n_300), .B(n_411), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_308), .B2(n_312), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_302), .A2(n_316), .B1(n_344), .B2(n_348), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_303), .A2(n_317), .B1(n_864), .B2(n_865), .Y(n_863) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g586 ( .A(n_304), .Y(n_586) );
INVx2_ASAP7_75t_SL g916 ( .A(n_304), .Y(n_916) );
BUFx8_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_305), .Y(n_315) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_305), .Y(n_425) );
INVx2_ASAP7_75t_L g570 ( .A(n_305), .Y(n_570) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x4_ASAP7_75t_L g557 ( .A(n_307), .B(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_308), .A2(n_761), .B1(n_762), .B2(n_764), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_308), .A2(n_586), .B1(n_861), .B2(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x6_ASAP7_75t_L g401 ( .A(n_310), .B(n_330), .Y(n_401) );
BUFx3_ASAP7_75t_L g979 ( .A(n_310), .Y(n_979) );
BUFx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g319 ( .A(n_311), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_312), .A2(n_320), .B1(n_338), .B2(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_317), .B2(n_320), .Y(n_313) );
INVx2_ASAP7_75t_L g977 ( .A(n_314), .Y(n_977) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_SL g448 ( .A(n_315), .Y(n_448) );
INVx5_ASAP7_75t_L g973 ( .A(n_315), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_317), .A2(n_569), .B1(n_583), .B2(n_584), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_317), .A2(n_916), .B1(n_917), .B2(n_918), .Y(n_915) );
BUFx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_319), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g765 ( .A1(n_323), .A2(n_766), .B1(n_768), .B2(n_769), .Y(n_765) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_323), .A2(n_766), .B1(n_805), .B2(n_811), .Y(n_819) );
INVx2_ASAP7_75t_L g886 ( .A(n_323), .Y(n_886) );
OAI22xp33_ASAP7_75t_L g919 ( .A1(n_323), .A2(n_907), .B1(n_920), .B2(n_921), .Y(n_919) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x4_ASAP7_75t_L g333 ( .A(n_326), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g535 ( .A(n_326), .Y(n_535) );
OR2x6_ASAP7_75t_L g593 ( .A(n_326), .B(n_328), .Y(n_593) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g669 ( .A(n_327), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_327), .B(n_1241), .Y(n_1256) );
INVx3_ASAP7_75t_L g1222 ( .A(n_328), .Y(n_1222) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND3x1_ASAP7_75t_L g565 ( .A(n_329), .B(n_330), .C(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g400 ( .A(n_330), .Y(n_400) );
AND2x4_ASAP7_75t_L g419 ( .A(n_330), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g1197 ( .A(n_330), .B(n_1198), .Y(n_1197) );
OAI33xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .A3(n_343), .B1(n_352), .B2(n_353), .B3(n_356), .Y(n_331) );
OAI33xp33_ASAP7_75t_L g594 ( .A1(n_332), .A2(n_356), .A3(n_595), .B1(n_596), .B2(n_597), .B3(n_600), .Y(n_594) );
OAI33xp33_ASAP7_75t_L g770 ( .A1(n_332), .A2(n_771), .A3(n_772), .B1(n_774), .B2(n_777), .B3(n_778), .Y(n_770) );
OAI33xp33_ASAP7_75t_L g869 ( .A1(n_332), .A2(n_356), .A3(n_870), .B1(n_872), .B2(n_873), .B3(n_874), .Y(n_869) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g455 ( .A(n_333), .Y(n_455) );
INVx4_ASAP7_75t_L g656 ( .A(n_333), .Y(n_656) );
INVx2_ASAP7_75t_L g985 ( .A(n_333), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_336), .A2(n_458), .B1(n_755), .B2(n_768), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_336), .A2(n_338), .B1(n_759), .B2(n_764), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_336), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_336), .A2(n_458), .B1(n_813), .B2(n_814), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g870 ( .A1(n_336), .A2(n_858), .B1(n_867), .B2(n_871), .Y(n_870) );
INVx4_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g989 ( .A(n_337), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_338), .A2(n_443), .B1(n_449), .B2(n_457), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_338), .A2(n_457), .B1(n_580), .B2(n_591), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_338), .A2(n_354), .B1(n_862), .B2(n_865), .Y(n_874) );
INVx4_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g459 ( .A(n_339), .Y(n_459) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_339), .Y(n_511) );
INVx2_ASAP7_75t_SL g804 ( .A(n_339), .Y(n_804) );
INVx1_ASAP7_75t_L g871 ( .A(n_339), .Y(n_871) );
INVx8_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g384 ( .A(n_340), .B(n_371), .Y(n_384) );
OR2x2_ASAP7_75t_L g468 ( .A(n_340), .B(n_364), .Y(n_468) );
BUFx2_ASAP7_75t_L g926 ( .A(n_340), .Y(n_926) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_344), .A2(n_441), .B1(n_447), .B2(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_344), .A2(n_348), .B1(n_861), .B2(n_864), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_344), .A2(n_776), .B1(n_859), .B2(n_868), .Y(n_873) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g598 ( .A(n_345), .Y(n_598) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g463 ( .A(n_346), .Y(n_463) );
INVx2_ASAP7_75t_L g517 ( .A(n_346), .Y(n_517) );
BUFx2_ASAP7_75t_L g775 ( .A(n_346), .Y(n_775) );
BUFx2_ASAP7_75t_L g1275 ( .A(n_346), .Y(n_1275) );
AND2x2_ASAP7_75t_L g530 ( .A(n_347), .B(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_348), .A2(n_758), .B1(n_761), .B2(n_773), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g1272 ( .A1(n_348), .A2(n_1218), .B1(n_1273), .B2(n_1276), .C(n_1277), .Y(n_1272) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g464 ( .A(n_349), .Y(n_464) );
INVx1_ASAP7_75t_L g513 ( .A(n_349), .Y(n_513) );
INVx1_ASAP7_75t_L g781 ( .A(n_349), .Y(n_781) );
INVx2_ASAP7_75t_L g992 ( .A(n_349), .Y(n_992) );
INVx4_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx4f_ASAP7_75t_L g361 ( .A(n_350), .Y(n_361) );
BUFx4f_ASAP7_75t_L g461 ( .A(n_350), .Y(n_461) );
BUFx4f_ASAP7_75t_L g521 ( .A(n_350), .Y(n_521) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_350), .Y(n_599) );
OR2x6_ASAP7_75t_L g1279 ( .A(n_350), .B(n_1280), .Y(n_1279) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g776 ( .A(n_351), .Y(n_776) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI33xp33_ASAP7_75t_L g454 ( .A1(n_356), .A2(n_455), .A3(n_456), .B1(n_460), .B2(n_462), .B3(n_465), .Y(n_454) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI33xp33_ASAP7_75t_L g654 ( .A1(n_357), .A2(n_655), .A3(n_657), .B1(n_659), .B2(n_663), .B3(n_664), .Y(n_654) );
INVx2_ASAP7_75t_L g778 ( .A(n_357), .Y(n_778) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_358), .A2(n_513), .B1(n_514), .B2(n_515), .C(n_518), .Y(n_512) );
AND2x4_ASAP7_75t_L g731 ( .A(n_358), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_358), .B(n_732), .Y(n_1264) );
OAI31xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_379), .A3(n_385), .B(n_393), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_361), .A2(n_463), .B1(n_583), .B2(n_587), .Y(n_596) );
NAND3xp33_ASAP7_75t_SL g613 ( .A(n_362), .B(n_614), .C(n_616), .Y(n_613) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g636 ( .A(n_363), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_363), .A2(n_710), .B(n_712), .C(n_713), .Y(n_709) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x2_ASAP7_75t_L g498 ( .A(n_364), .B(n_372), .Y(n_498) );
AND2x2_ASAP7_75t_L g895 ( .A(n_364), .B(n_495), .Y(n_895) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g711 ( .A(n_366), .Y(n_711) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_367), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_373), .B2(n_374), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g614 ( .A1(n_370), .A2(n_474), .B1(n_494), .B2(n_607), .C1(n_608), .C2(n_615), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_370), .A2(n_888), .B1(n_897), .B2(n_898), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_370), .A2(n_943), .B1(n_955), .B2(n_956), .Y(n_954) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x4_ASAP7_75t_L g472 ( .A(n_371), .B(n_372), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_371), .A2(n_493), .B(n_494), .C(n_496), .Y(n_492) );
INVx1_ASAP7_75t_L g501 ( .A(n_371), .Y(n_501) );
AND2x2_ASAP7_75t_L g618 ( .A(n_371), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g1258 ( .A(n_372), .Y(n_1258) );
AOI32xp33_ASAP7_75t_L g408 ( .A1(n_373), .A2(n_409), .A3(n_413), .B1(n_415), .B2(n_417), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_374), .A2(n_498), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_374), .A2(n_498), .B1(n_783), .B2(n_784), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g1317 ( .A1(n_374), .A2(n_498), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx3_ASAP7_75t_L g474 ( .A(n_376), .Y(n_474) );
INVx2_ASAP7_75t_L g715 ( .A(n_376), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_377), .B(n_1241), .Y(n_1260) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g708 ( .A(n_380), .Y(n_708) );
BUFx3_ASAP7_75t_L g457 ( .A(n_381), .Y(n_457) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_381), .Y(n_601) );
INVx2_ASAP7_75t_SL g925 ( .A(n_381), .Y(n_925) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_383), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g717 ( .A(n_384), .Y(n_717) );
BUFx2_ASAP7_75t_L g786 ( .A(n_384), .Y(n_786) );
BUFx2_ASAP7_75t_L g958 ( .A(n_386), .Y(n_958) );
AND2x4_ASAP7_75t_L g390 ( .A(n_387), .B(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
INVx4_ASAP7_75t_L g477 ( .A(n_390), .Y(n_477) );
INVx3_ASAP7_75t_SL g491 ( .A(n_390), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_390), .A2(n_694), .B1(n_695), .B2(n_708), .Y(n_707) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_391), .Y(n_524) );
BUFx3_ASAP7_75t_L g724 ( .A(n_391), .Y(n_724) );
OAI31xp33_ASAP7_75t_L g779 ( .A1(n_393), .A2(n_780), .A3(n_785), .B(n_787), .Y(n_779) );
OAI31xp33_ASAP7_75t_L g820 ( .A1(n_393), .A2(n_821), .A3(n_825), .B(n_826), .Y(n_820) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_394), .A2(n_467), .A3(n_469), .B(n_475), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_394), .A2(n_613), .B(n_622), .Y(n_612) );
INVx1_ASAP7_75t_L g641 ( .A(n_394), .Y(n_641) );
BUFx2_ASAP7_75t_SL g718 ( .A(n_394), .Y(n_718) );
BUFx3_ASAP7_75t_L g962 ( .A(n_394), .Y(n_962) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_396), .B(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1283 ( .A(n_396), .Y(n_1283) );
OAI31xp33_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_402), .A3(n_421), .B(n_426), .Y(n_397) );
INVx2_ASAP7_75t_SL g703 ( .A(n_399), .Y(n_703) );
BUFx3_ASAP7_75t_L g947 ( .A(n_399), .Y(n_947) );
BUFx2_ASAP7_75t_L g1332 ( .A(n_399), .Y(n_1332) );
AND2x2_ASAP7_75t_L g424 ( .A(n_400), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g651 ( .A(n_400), .B(n_425), .Y(n_651) );
INVx2_ASAP7_75t_L g611 ( .A(n_401), .Y(n_611) );
INVx1_ASAP7_75t_L g705 ( .A(n_401), .Y(n_705) );
INVx1_ASAP7_75t_L g883 ( .A(n_401), .Y(n_883) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_404), .A2(n_415), .B1(n_842), .B2(n_851), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_404), .A2(n_647), .B1(n_888), .B2(n_889), .Y(n_887) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
AND2x2_ASAP7_75t_L g415 ( .A(n_405), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g485 ( .A(n_405), .B(n_407), .Y(n_485) );
AND2x4_ASAP7_75t_L g647 ( .A(n_405), .B(n_416), .Y(n_647) );
AND2x2_ASAP7_75t_L g942 ( .A(n_405), .B(n_407), .Y(n_942) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g409 ( .A(n_406), .B(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_409), .A2(n_471), .B1(n_484), .B2(n_485), .Y(n_483) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_410), .B(n_1197), .Y(n_1211) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x6_ASAP7_75t_L g1209 ( .A(n_413), .B(n_1197), .Y(n_1209) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
INVxp67_ASAP7_75t_L g543 ( .A(n_415), .Y(n_543) );
AOI222xp33_ASAP7_75t_L g604 ( .A1(n_415), .A2(n_485), .B1(n_605), .B2(n_606), .C1(n_607), .C2(n_608), .Y(n_604) );
INVx1_ASAP7_75t_L g700 ( .A(n_415), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_415), .A2(n_485), .B1(n_783), .B2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_415), .A2(n_485), .B1(n_823), .B2(n_831), .Y(n_830) );
CKINVDCx8_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g538 ( .A(n_419), .B(n_539), .C(n_544), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_419), .B(n_644), .C(n_645), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_419), .A2(n_697), .B(n_698), .C(n_699), .Y(n_696) );
CKINVDCx8_ASAP7_75t_R g794 ( .A(n_419), .Y(n_794) );
AOI211xp5_ASAP7_75t_L g1326 ( .A1(n_419), .A2(n_1319), .B(n_1327), .C(n_1328), .Y(n_1326) );
BUFx2_ASAP7_75t_L g559 ( .A(n_420), .Y(n_559) );
BUFx2_ASAP7_75t_L g605 ( .A(n_420), .Y(n_605) );
INVx2_ASAP7_75t_L g674 ( .A(n_420), .Y(n_674) );
BUFx2_ASAP7_75t_L g686 ( .A(n_420), .Y(n_686) );
BUFx2_ASAP7_75t_L g698 ( .A(n_420), .Y(n_698) );
BUFx3_ASAP7_75t_L g739 ( .A(n_420), .Y(n_739) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_420), .B(n_1232), .Y(n_1234) );
INVx1_ASAP7_75t_L g546 ( .A(n_422), .Y(n_546) );
INVx2_ASAP7_75t_SL g650 ( .A(n_422), .Y(n_650) );
INVx2_ASAP7_75t_SL g936 ( .A(n_422), .Y(n_936) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_424), .A2(n_500), .B1(n_546), .B2(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g442 ( .A(n_425), .Y(n_442) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_425), .Y(n_554) );
INVx2_ASAP7_75t_L g677 ( .A(n_425), .Y(n_677) );
INVx1_ASAP7_75t_L g682 ( .A(n_425), .Y(n_682) );
OAI31xp33_ASAP7_75t_SL g478 ( .A1(n_426), .A2(n_479), .A3(n_480), .B(n_481), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_426), .A2(n_603), .B(n_609), .Y(n_602) );
OAI31xp33_ASAP7_75t_SL g788 ( .A1(n_426), .A2(n_789), .A3(n_790), .B(n_797), .Y(n_788) );
OAI31xp33_ASAP7_75t_SL g827 ( .A1(n_426), .A2(n_828), .A3(n_829), .B(n_832), .Y(n_827) );
OAI31xp33_ASAP7_75t_L g846 ( .A1(n_426), .A2(n_847), .A3(n_849), .B(n_854), .Y(n_846) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
AND2x2_ASAP7_75t_SL g548 ( .A(n_427), .B(n_429), .Y(n_548) );
AND2x2_ASAP7_75t_L g653 ( .A(n_427), .B(n_429), .Y(n_653) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_466), .C(n_478), .Y(n_432) );
NOR2xp33_ASAP7_75t_SL g433 ( .A(n_434), .B(n_454), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_436), .A2(n_452), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g969 ( .A(n_438), .Y(n_969) );
INVx2_ASAP7_75t_L g1225 ( .A(n_438), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_439), .A2(n_453), .B1(n_463), .B2(n_464), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_442), .A2(n_444), .B1(n_758), .B2(n_759), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_442), .A2(n_444), .B1(n_807), .B2(n_813), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_442), .A2(n_450), .B1(n_1302), .B2(n_1339), .C(n_1340), .Y(n_1338) );
OAI221xp5_ASAP7_75t_L g1217 ( .A1(n_444), .A2(n_973), .B1(n_1218), .B2(n_1219), .C(n_1220), .Y(n_1217) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g450 ( .A(n_445), .Y(n_450) );
CKINVDCx8_ASAP7_75t_R g571 ( .A(n_445), .Y(n_571) );
INVx3_ASAP7_75t_L g588 ( .A(n_445), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_449), .B2(n_450), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_448), .A2(n_588), .B1(n_808), .B2(n_814), .Y(n_818) );
OAI33xp33_ASAP7_75t_L g801 ( .A1(n_455), .A2(n_778), .A3(n_802), .B1(n_806), .B2(n_809), .B3(n_812), .Y(n_801) );
BUFx6f_ASAP7_75t_L g1271 ( .A(n_455), .Y(n_1271) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_458), .A2(n_584), .B1(n_589), .B2(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g1300 ( .A1(n_461), .A2(n_598), .B1(n_1301), .B2(n_1302), .C(n_1303), .Y(n_1300) );
INVx1_ASAP7_75t_L g621 ( .A(n_468), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g714 ( .A(n_472), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_472), .A2(n_474), .B1(n_842), .B2(n_843), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_474), .A2(n_498), .B1(n_823), .B2(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_485), .B(n_638), .Y(n_648) );
XOR2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_575), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_534), .B(n_536), .Y(n_488) );
BUFx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_495), .Y(n_662) );
BUFx3_ASAP7_75t_L g725 ( .A(n_495), .Y(n_725) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_512), .B(n_519), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_506) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_509), .A2(n_520), .B1(n_569), .B2(n_571), .C(n_572), .Y(n_568) );
INVx5_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx6_ASAP7_75t_L g990 ( .A(n_511), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_515), .A2(n_971), .B1(n_978), .B2(n_992), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_515), .A2(n_781), .B1(n_968), .B2(n_983), .Y(n_993) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g773 ( .A(n_517), .Y(n_773) );
OAI211xp5_ASAP7_75t_SL g519 ( .A1(n_520), .A2(n_521), .B(n_522), .C(n_527), .Y(n_519) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g661 ( .A(n_524), .Y(n_661) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_524), .B(n_1245), .Y(n_1288) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g727 ( .A(n_529), .Y(n_727) );
INVx2_ASAP7_75t_L g1304 ( .A(n_529), .Y(n_1304) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_530), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_530), .B(n_1241), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_530), .B(n_1245), .Y(n_1284) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g1247 ( .A(n_533), .Y(n_1247) );
BUFx3_ASAP7_75t_L g1267 ( .A(n_533), .Y(n_1267) );
BUFx6f_ASAP7_75t_L g1278 ( .A(n_533), .Y(n_1278) );
OAI21xp5_ASAP7_75t_L g1192 ( .A1(n_534), .A2(n_1193), .B(n_1216), .Y(n_1192) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_548), .B(n_549), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_538), .B(n_545), .Y(n_537) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g939 ( .A(n_541), .Y(n_939) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_548), .A2(n_692), .B1(n_706), .B2(n_718), .C(n_719), .Y(n_691) );
BUFx2_ASAP7_75t_L g948 ( .A(n_548), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B1(n_563), .B2(n_568), .Y(n_549) );
OAI33xp33_ASAP7_75t_L g578 ( .A1(n_550), .A2(n_579), .A3(n_582), .B1(n_585), .B2(n_590), .B3(n_593), .Y(n_578) );
OAI33xp33_ASAP7_75t_L g903 ( .A1(n_550), .A2(n_593), .A3(n_904), .B1(n_911), .B2(n_915), .B3(n_919), .Y(n_903) );
OAI33xp33_ASAP7_75t_L g964 ( .A1(n_550), .A2(n_563), .A3(n_965), .B1(n_970), .B2(n_975), .B3(n_981), .Y(n_964) );
OAI22xp33_ASAP7_75t_L g1333 ( .A1(n_550), .A2(n_1334), .B1(n_1338), .B2(n_1341), .Y(n_1333) );
OAI211xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B(n_555), .C(n_560), .Y(n_551) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx8_ASAP7_75t_L g574 ( .A(n_557), .Y(n_574) );
BUFx3_ASAP7_75t_L g672 ( .A(n_557), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g1196 ( .A(n_557), .B(n_1197), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_557), .B(n_1232), .Y(n_1231) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx5_ASAP7_75t_L g679 ( .A(n_562), .Y(n_679) );
BUFx12f_ASAP7_75t_L g737 ( .A(n_562), .Y(n_737) );
AND2x4_ASAP7_75t_L g1207 ( .A(n_562), .B(n_1204), .Y(n_1207) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g743 ( .A(n_565), .Y(n_743) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g1238 ( .A(n_567), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_567), .B(n_1245), .Y(n_1244) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx3_ASAP7_75t_L g763 ( .A(n_570), .Y(n_763) );
OR2x6_ASAP7_75t_SL g1202 ( .A(n_570), .B(n_1203), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_571), .A2(n_971), .B1(n_972), .B2(n_974), .Y(n_970) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx8_ASAP7_75t_L g685 ( .A(n_574), .Y(n_685) );
INVx3_ASAP7_75t_L g1337 ( .A(n_574), .Y(n_1337) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_602), .C(n_612), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_594), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_581), .A2(n_592), .B1(n_598), .B2(n_599), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_588), .A2(n_912), .B1(n_913), .B2(n_914), .Y(n_911) );
INVx1_ASAP7_75t_L g687 ( .A(n_593), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_599), .A2(n_773), .B1(n_810), .B2(n_811), .Y(n_809) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_599), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_599), .A2(n_1306), .B1(n_1307), .B2(n_1308), .C(n_1309), .Y(n_1305) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g1330 ( .A1(n_611), .A2(n_1314), .B1(n_1315), .B2(n_1331), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_620), .B2(n_621), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_618), .A2(n_702), .B1(n_704), .B2(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_618), .A2(n_960), .B1(n_1314), .B2(n_1315), .C(n_1316), .Y(n_1313) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_619), .Y(n_658) );
INVx3_ASAP7_75t_L g666 ( .A(n_619), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_834), .B2(n_997), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_747), .B2(n_833), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
XNOR2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_690), .Y(n_627) );
INVx1_ASAP7_75t_L g688 ( .A(n_629), .Y(n_688) );
NAND4xp75_ASAP7_75t_L g629 ( .A(n_630), .B(n_642), .C(n_654), .D(n_667), .Y(n_629) );
AO21x1_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B(n_641), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_632), .A2(n_633), .B1(n_650), .B2(n_651), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_640), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g1316 ( .A(n_636), .B(n_1317), .C(n_1320), .Y(n_1316) );
AOI21xp33_ASAP7_75t_L g1312 ( .A1(n_641), .A2(n_1313), .B(n_1322), .Y(n_1312) );
AO21x1_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_649), .B(n_652), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx6f_ASAP7_75t_L g944 ( .A(n_647), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_650), .A2(n_651), .B1(n_694), .B2(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g848 ( .A(n_651), .Y(n_848) );
INVx2_ASAP7_75t_L g891 ( .A(n_651), .Y(n_891) );
INVx2_ASAP7_75t_L g937 ( .A(n_651), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_651), .A2(n_936), .B1(n_1323), .B2(n_1324), .Y(n_1329) );
AOI31xp33_ASAP7_75t_L g1325 ( .A1(n_652), .A2(n_1326), .A3(n_1329), .B(n_1330), .Y(n_1325) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI31xp33_ASAP7_75t_L g880 ( .A1(n_653), .A2(n_881), .A3(n_884), .B(n_890), .Y(n_880) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_655), .Y(n_728) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
OAI33xp33_ASAP7_75t_L g922 ( .A1(n_656), .A2(n_778), .A3(n_923), .B1(n_927), .B2(n_929), .B3(n_930), .Y(n_922) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_662), .B(n_1321), .Y(n_1320) );
INVx2_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g1266 ( .A(n_666), .Y(n_1266) );
AOI33xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .A3(n_675), .B1(n_680), .B2(n_684), .B3(n_687), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_668), .B(n_736), .C(n_738), .Y(n_735) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g746 ( .A(n_672), .Y(n_746) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g1327 ( .A(n_674), .Y(n_1327) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g1334 ( .A1(n_677), .A2(n_979), .B1(n_1301), .B2(n_1335), .C(n_1336), .Y(n_1334) );
INVx2_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g683 ( .A(n_679), .Y(n_683) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_696), .C(n_701), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .C(n_716), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g898 ( .A(n_715), .Y(n_898) );
INVx2_ASAP7_75t_L g955 ( .A(n_715), .Y(n_955) );
INVxp67_ASAP7_75t_SL g900 ( .A(n_717), .Y(n_900) );
OAI31xp33_ASAP7_75t_SL g838 ( .A1(n_718), .A2(n_839), .A3(n_844), .B(n_845), .Y(n_838) );
OAI31xp33_ASAP7_75t_L g892 ( .A1(n_718), .A2(n_893), .A3(n_899), .B(n_901), .Y(n_892) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_729), .C(n_735), .D(n_740), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_726), .C(n_728), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .C(n_734), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_731), .Y(n_994) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_739), .Y(n_853) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .C(n_744), .Y(n_740) );
BUFx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_L g1342 ( .A(n_743), .Y(n_1342) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g833 ( .A(n_748), .Y(n_833) );
XNOR2x1_ASAP7_75t_L g748 ( .A(n_749), .B(n_798), .Y(n_748) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
AND3x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_779), .C(n_788), .Y(n_751) );
NOR2xp33_ASAP7_75t_SL g752 ( .A(n_753), .B(n_770), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_756), .A2(n_769), .B1(n_775), .B2(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g913 ( .A(n_763), .Y(n_913) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx3_ASAP7_75t_L g907 ( .A(n_767), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_773), .A2(n_776), .B1(n_807), .B2(n_808), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_775), .A2(n_912), .B1(n_917), .B2(n_928), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_775), .A2(n_908), .B1(n_921), .B2(n_928), .Y(n_929) );
BUFx3_ASAP7_75t_L g928 ( .A(n_776), .Y(n_928) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_776), .B(n_1244), .Y(n_1250) );
INVx2_ASAP7_75t_SL g960 ( .A(n_786), .Y(n_960) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_791), .A2(n_967), .B1(n_982), .B2(n_983), .Y(n_981) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g910 ( .A(n_793), .Y(n_910) );
OR2x6_ASAP7_75t_L g1214 ( .A(n_793), .B(n_1215), .Y(n_1214) );
NAND3xp33_ASAP7_75t_L g849 ( .A(n_794), .B(n_850), .C(n_852), .Y(n_849) );
AND3x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_820), .C(n_827), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_815), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_804), .A2(n_914), .B1(n_918), .B2(n_924), .Y(n_930) );
INVx1_ASAP7_75t_L g997 ( .A(n_834), .Y(n_997) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_875), .Y(n_834) );
INVx2_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_846), .C(n_855), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_843), .B(n_853), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_869), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_877), .B1(n_931), .B2(n_996), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NAND3xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_892), .C(n_902), .Y(n_879) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g953 ( .A(n_895), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_922), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_908), .B2(n_909), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_905), .A2(n_920), .B1(n_924), .B2(n_926), .Y(n_923) );
BUFx4f_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g952 ( .A(n_928), .Y(n_952) );
INVx1_ASAP7_75t_L g996 ( .A(n_931), .Y(n_996) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_949), .C(n_963), .Y(n_932) );
OAI31xp33_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_938), .A3(n_946), .B(n_948), .Y(n_933) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_943), .B1(n_944), .B2(n_945), .Y(n_940) );
BUFx3_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
OAI31xp33_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_957), .A3(n_961), .B(n_962), .Y(n_949) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_984), .Y(n_963) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_966), .A2(n_982), .B1(n_987), .B2(n_990), .Y(n_986) );
BUFx3_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_974), .A2(n_980), .B1(n_987), .B2(n_990), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OAI33xp33_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .A3(n_991), .B1(n_993), .B2(n_994), .B3(n_995), .Y(n_984) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx2_ASAP7_75t_SL g988 ( .A(n_989), .Y(n_988) );
OAI21xp5_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1006), .B(n_1187), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_1000), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_1001), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g1076 ( .A1(n_1001), .A2(n_1077), .B1(n_1078), .B2(n_1079), .C(n_1080), .Y(n_1076) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
AND2x6_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1004), .Y(n_1002) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_1003), .B(n_1016), .Y(n_1015) );
AND2x6_ASAP7_75t_L g1019 ( .A(n_1003), .B(n_1020), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_1003), .B(n_1022), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1003), .B(n_1022), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1003), .B(n_1022), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1003), .B(n_1016), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1348 ( .A(n_1004), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_1005), .B(n_1017), .Y(n_1016) );
NOR2xp67_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1125), .Y(n_1006) );
NAND4xp25_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1081), .C(n_1105), .D(n_1119), .Y(n_1007) );
OAI21xp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1066), .B(n_1072), .Y(n_1008) );
OAI321xp33_ASAP7_75t_L g1009 ( .A1(n_1010), .A2(n_1031), .A3(n_1042), .B1(n_1046), .B2(n_1049), .C(n_1052), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1011), .B(n_1083), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1023), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_1012), .B(n_1050), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1012), .B(n_1024), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1012), .B(n_1097), .Y(n_1107) );
NOR2xp33_ASAP7_75t_L g1171 ( .A(n_1012), .B(n_1098), .Y(n_1171) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_1013), .B(n_1071), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1013), .B(n_1025), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1013), .B(n_1098), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1013), .B(n_1134), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1013), .B(n_1098), .Y(n_1157) );
NAND2xp5_ASAP7_75t_SL g1166 ( .A(n_1013), .B(n_1057), .Y(n_1166) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1013), .B(n_1057), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1018), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1014), .B(n_1018), .Y(n_1088) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1028), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1025), .B(n_1051), .Y(n_1050) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1025), .Y(n_1098) );
AOI321xp33_ASAP7_75t_L g1119 ( .A1(n_1025), .A2(n_1082), .A3(n_1115), .B1(n_1120), .B2(n_1122), .C(n_1124), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1025), .B(n_1028), .Y(n_1134) );
NAND2x1p5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1028), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_1028), .B(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1028), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1028), .B(n_1098), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1030), .Y(n_1028) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1032), .B(n_1085), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1037), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_1033), .B(n_1042), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1033), .B(n_1048), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1033), .B(n_1042), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1033), .B(n_1065), .Y(n_1102) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1033), .B(n_1038), .Y(n_1116) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1033), .Y(n_1132) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1033), .Y(n_1155) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_1034), .B(n_1065), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_1037), .B(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1037), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1037), .B(n_1085), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1037), .B(n_1086), .Y(n_1110) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1038), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1041), .Y(n_1038) );
INVx3_ASAP7_75t_L g1048 ( .A(n_1042), .Y(n_1048) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1042), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1044), .Y(n_1042) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
OAI322xp33_ASAP7_75t_L g1150 ( .A1(n_1047), .A2(n_1049), .A3(n_1088), .B1(n_1151), .B2(n_1153), .C1(n_1154), .C2(n_1155), .Y(n_1150) );
CKINVDCx14_ASAP7_75t_R g1139 ( .A(n_1048), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1048), .B(n_1121), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1048), .B(n_1102), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1048), .B(n_1064), .Y(n_1185) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1049), .Y(n_1111) );
AOI21xp33_ASAP7_75t_SL g1112 ( .A1(n_1049), .A2(n_1113), .B(n_1114), .Y(n_1112) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1050), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_1050), .B(n_1088), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1050), .B(n_1152), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1050), .B(n_1166), .Y(n_1165) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1055), .B1(n_1061), .B2(n_1062), .Y(n_1052) );
OAI21xp5_ASAP7_75t_L g1148 ( .A1(n_1053), .A2(n_1096), .B(n_1149), .Y(n_1148) );
CKINVDCx14_ASAP7_75t_R g1053 ( .A(n_1054), .Y(n_1053) );
NOR3xp33_ASAP7_75t_L g1124 ( .A(n_1054), .B(n_1057), .C(n_1095), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1054), .B(n_1060), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1060), .Y(n_1056) );
INVx4_ASAP7_75t_L g1063 ( .A(n_1057), .Y(n_1063) );
INVx4_ASAP7_75t_L g1086 ( .A(n_1057), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1057), .B(n_1107), .Y(n_1106) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1057), .B(n_1157), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1057), .B(n_1116), .Y(n_1174) );
AND2x4_ASAP7_75t_SL g1057 ( .A(n_1058), .B(n_1059), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1061), .B(n_1086), .Y(n_1136) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1062), .Y(n_1069) );
AOI21xp33_ASAP7_75t_L g1135 ( .A1(n_1062), .A2(n_1071), .B(n_1136), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1062), .B(n_1118), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
CKINVDCx5p33_ASAP7_75t_R g1083 ( .A(n_1063), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1149 ( .A(n_1063), .B(n_1070), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1063), .B(n_1087), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1063), .B(n_1171), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1064), .B(n_1068), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_1064), .A2(n_1098), .B1(n_1104), .B2(n_1127), .C(n_1128), .Y(n_1126) );
NOR3xp33_ASAP7_75t_L g1164 ( .A(n_1064), .B(n_1165), .C(n_1167), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_1064), .A2(n_1132), .B1(n_1170), .B2(n_1172), .Y(n_1169) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
AOI21xp33_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1069), .B(n_1070), .Y(n_1066) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1067), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1068), .B(n_1093), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_1068), .A2(n_1106), .B1(n_1108), .B2(n_1109), .C(n_1112), .Y(n_1105) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1068), .Y(n_1176) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1070), .Y(n_1130) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
OAI321xp33_ASAP7_75t_L g1125 ( .A1(n_1073), .A2(n_1074), .A3(n_1126), .B1(n_1137), .B2(n_1140), .C(n_1163), .Y(n_1125) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1076), .B(n_1086), .Y(n_1123) );
O2A1O1Ixp33_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1084), .B(n_1089), .C(n_1090), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1083), .B(n_1101), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1083), .B(n_1120), .Y(n_1145) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1087), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1085), .B(n_1118), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_1086), .Y(n_1085) );
NAND2xp5_ASAP7_75t_SL g1129 ( .A(n_1086), .B(n_1130), .Y(n_1129) );
NAND2x1_ASAP7_75t_L g1142 ( .A(n_1086), .B(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1087), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1088), .B(n_1097), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1088), .B(n_1133), .Y(n_1162) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1089), .Y(n_1167) );
OAI221xp5_ASAP7_75t_L g1090 ( .A1(n_1091), .A2(n_1094), .B1(n_1095), .B2(n_1099), .C(n_1103), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
OAI21xp5_ASAP7_75t_SL g1103 ( .A1(n_1092), .A2(n_1100), .B(n_1104), .Y(n_1103) );
INVxp67_ASAP7_75t_L g1158 ( .A(n_1093), .Y(n_1158) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1094), .B(n_1183), .Y(n_1182) );
OAI32xp33_ASAP7_75t_L g1184 ( .A1(n_1095), .A2(n_1102), .A3(n_1123), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1097), .Y(n_1152) );
NAND3xp33_ASAP7_75t_L g1154 ( .A(n_1097), .B(n_1110), .C(n_1118), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1097), .B(n_1178), .Y(n_1186) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_1102), .Y(n_1101) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_1102), .A2(n_1129), .B1(n_1131), .B2(n_1133), .C(n_1135), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1117), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1116), .B(n_1118), .Y(n_1183) );
OAI21xp33_ASAP7_75t_L g1168 ( .A1(n_1118), .A2(n_1169), .B(n_1173), .Y(n_1168) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_1121), .Y(n_1120) );
OAI322xp33_ASAP7_75t_L g1175 ( .A1(n_1121), .A2(n_1123), .A3(n_1162), .B1(n_1176), .B2(n_1177), .C1(n_1180), .C2(n_1181), .Y(n_1175) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AOI21xp33_ASAP7_75t_L g1137 ( .A1(n_1127), .A2(n_1138), .B(n_1139), .Y(n_1137) );
NOR2xp33_ASAP7_75t_L g1141 ( .A(n_1131), .B(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1134), .B(n_1178), .Y(n_1177) );
CKINVDCx14_ASAP7_75t_R g1147 ( .A(n_1138), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1138), .B(n_1174), .Y(n_1173) );
O2A1O1Ixp33_ASAP7_75t_L g1156 ( .A1(n_1139), .A2(n_1157), .B(n_1158), .C(n_1159), .Y(n_1156) );
NOR5xp2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1144), .C(n_1150), .D(n_1156), .E(n_1160), .Y(n_1140) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1143), .Y(n_1181) );
A2O1A1Ixp33_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1146), .B(n_1147), .C(n_1148), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
NOR5xp2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1168), .C(n_1175), .D(n_1182), .E(n_1184), .Y(n_1163) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1191), .Y(n_1289) );
NAND4xp25_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1235), .C(n_1251), .D(n_1281), .Y(n_1191) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1197), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_1200), .A2(n_1201), .B1(n_1206), .B2(n_1207), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_1200), .A2(n_1230), .B1(n_1282), .B2(n_1285), .Y(n_1281) );
CKINVDCx5p33_ASAP7_75t_R g1201 ( .A(n_1202), .Y(n_1201) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1205), .Y(n_1232) );
AOI222xp33_ASAP7_75t_L g1235 ( .A1(n_1206), .A2(n_1212), .B1(n_1236), .B2(n_1242), .C1(n_1248), .C2(n_1249), .Y(n_1235) );
AOI221xp5_ASAP7_75t_L g1208 ( .A1(n_1209), .A2(n_1210), .B1(n_1211), .B2(n_1212), .C(n_1213), .Y(n_1208) );
CKINVDCx5p33_ASAP7_75t_R g1213 ( .A(n_1214), .Y(n_1213) );
NAND3xp33_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1223), .C(n_1229), .Y(n_1216) );
INVx3_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
OAI211xp5_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1225), .B(n_1226), .C(n_1228), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1231), .B1(n_1233), .B2(n_1234), .Y(n_1229) );
AND2x4_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1239), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
AND2x4_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1246), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
INVx3_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1268), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
NAND2x2_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1257), .Y(n_1254) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1255), .Y(n_1280) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx2_ASAP7_75t_SL g1257 ( .A(n_1258), .Y(n_1257) );
NAND3xp33_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1263), .C(n_1265), .Y(n_1261) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI22xp33_ASAP7_75t_L g1299 ( .A1(n_1264), .A2(n_1271), .B1(n_1300), .B2(n_1305), .Y(n_1299) );
OAI21xp5_ASAP7_75t_L g1268 ( .A1(n_1269), .A2(n_1272), .B(n_1279), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1274), .Y(n_1306) );
INVx4_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1278), .Y(n_1311) );
AND2x4_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1283), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVxp67_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
HB1xp67_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
NOR4xp25_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1312), .C(n_1325), .D(n_1333), .Y(n_1298) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
HB1xp67_ASAP7_75t_SL g1343 ( .A(n_1344), .Y(n_1343) );
INVx2_ASAP7_75t_SL g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
OAI21xp5_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1349), .B(n_1350), .Y(n_1347) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
endmodule