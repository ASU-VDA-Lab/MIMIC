module fake_aes_10054_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_L g3 ( .A(n_0), .B(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_4), .Y(n_5) );
INVx1_ASAP7_75t_SL g6 ( .A(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
OAI221xp5_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_5), .B1(n_3), .B2(n_0), .C(n_1), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
NOR3xp33_ASAP7_75t_L g11 ( .A(n_9), .B(n_8), .C(n_1), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
NAND3xp33_ASAP7_75t_SL g13 ( .A(n_12), .B(n_11), .C(n_8), .Y(n_13) );
endmodule