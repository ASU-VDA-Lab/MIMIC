module real_jpeg_14260_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_3),
.A2(n_36),
.B1(n_43),
.B2(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_48),
.B1(n_55),
.B2(n_57),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_48),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_6),
.A2(n_36),
.B1(n_43),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_55),
.B1(n_57),
.B2(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_61),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_7),
.A2(n_36),
.B1(n_43),
.B2(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_7),
.A2(n_55),
.B1(n_57),
.B2(n_70),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_70),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_55),
.B1(n_57),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_8),
.A2(n_36),
.B1(n_43),
.B2(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_9),
.A2(n_31),
.B1(n_55),
.B2(n_57),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_13),
.B(n_91),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_13),
.B(n_26),
.C(n_80),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_13),
.A2(n_41),
.B1(n_55),
.B2(n_57),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_94),
.B1(n_98),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_13),
.B(n_59),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_14),
.A2(n_36),
.B1(n_43),
.B2(n_68),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_55),
.B1(n_57),
.B2(n_68),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_15),
.A2(n_33),
.B1(n_55),
.B2(n_57),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_105),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_92),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_45),
.B1(n_71),
.B2(n_72),
.Y(n_20)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_22),
.A2(n_23),
.B1(n_34),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_23)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_24),
.B(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_24),
.A2(n_97),
.B(n_124),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_24),
.A2(n_28),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_25),
.A2(n_26),
.B1(n_78),
.B2(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_25),
.B(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_28),
.B(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_30),
.A2(n_98),
.B(n_121),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_34),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.C(n_42),
.Y(n_34)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_43),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_36),
.B(n_41),
.CON(n_159),
.SN(n_159)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_36),
.B(n_53),
.C(n_57),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_37),
.A2(n_67),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.CON(n_37),
.SN(n_37)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_43),
.C(n_44),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_41),
.B(n_98),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_41),
.B(n_101),
.Y(n_202)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_62),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_46),
.B(n_62),
.C(n_71),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_58),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_49),
.B1(n_54),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_49),
.A2(n_54),
.B1(n_88),
.B2(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_60),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_50),
.A2(n_59),
.B1(n_143),
.B2(n_159),
.Y(n_161)
);

AND2x4_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_52),
.A2(n_55),
.B(n_159),
.C(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_57),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_55),
.B(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_65),
.B1(n_69),
.B2(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_92),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_86),
.C(n_89),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_74),
.A2(n_75),
.B1(n_86),
.B2(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_82),
.B(n_83),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_76),
.A2(n_101),
.B1(n_102),
.B2(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_76),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_76),
.A2(n_101),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_76),
.A2(n_101),
.B1(n_164),
.B2(n_189),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_SL g80 ( 
.A(n_78),
.Y(n_80)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_81),
.A2(n_104),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_81),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_100),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_94),
.A2(n_98),
.B1(n_192),
.B2(n_200),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_94),
.A2(n_123),
.B(n_194),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_125),
.B2(n_126),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_229),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_149),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_147),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_134),
.B(n_147),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_140),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_135),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_223),
.B(n_228),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_178),
.B(n_222),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_166),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_152),
.B(n_166),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_161),
.C(n_162),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_153),
.A2(n_154),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_162),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_167),
.B(n_172),
.C(n_176),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_216),
.B(n_221),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_206),
.B(n_215),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_195),
.B(n_205),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_190),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_201),
.B(n_204),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_220)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.Y(n_221)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_227),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);


endmodule