module fake_jpeg_7068_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_38),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_51),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_17),
.B1(n_23),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_23),
.B1(n_32),
.B2(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_23),
.B1(n_17),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_39),
.B1(n_20),
.B2(n_35),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_18),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_23),
.B1(n_17),
.B2(n_32),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_21),
.C(n_29),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_45),
.C(n_22),
.Y(n_80)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_83),
.B(n_96),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_82),
.B1(n_34),
.B2(n_19),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_39),
.B1(n_20),
.B2(n_35),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_27),
.B1(n_33),
.B2(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_19),
.B1(n_27),
.B2(n_28),
.Y(n_82)
);

AND2x4_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_88),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_37),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_22),
.B1(n_27),
.B2(n_34),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_22),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_116),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_37),
.A3(n_54),
.B1(n_58),
.B2(n_61),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_104),
.C(n_127),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_89),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_70),
.B1(n_62),
.B2(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_108),
.B1(n_120),
.B2(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_98),
.B1(n_82),
.B2(n_96),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_64),
.B1(n_47),
.B2(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_52),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_123),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_126),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_47),
.B1(n_48),
.B2(n_30),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_58),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_58),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_117),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_97),
.B1(n_75),
.B2(n_85),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_130),
.B1(n_145),
.B2(n_150),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_85),
.B(n_72),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_14),
.C(n_15),
.Y(n_183)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_140),
.B(n_152),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_77),
.B(n_92),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_151),
.B(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_86),
.B1(n_94),
.B2(n_88),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_134),
.B1(n_139),
.B2(n_147),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_99),
.B1(n_71),
.B2(n_74),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_40),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_73),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_154),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_155),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_86),
.B1(n_74),
.B2(n_73),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_125),
.B(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_99),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_100),
.B(n_71),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_158),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_114),
.C(n_101),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_165),
.C(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_106),
.B1(n_112),
.B2(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_170),
.B1(n_172),
.B2(n_190),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_102),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_163),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_167),
.B(n_168),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_128),
.C(n_133),
.Y(n_165)
);

AO22x1_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_108),
.B1(n_107),
.B2(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_166),
.A2(n_178),
.B1(n_183),
.B2(n_31),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_95),
.B(n_37),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_67),
.C(n_40),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_53),
.B1(n_46),
.B2(n_44),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_24),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_53),
.B1(n_46),
.B2(n_44),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_152),
.Y(n_197)
);

OAI22x1_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_67),
.B1(n_25),
.B2(n_30),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_155),
.B1(n_25),
.B2(n_30),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_25),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_149),
.B(n_157),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_40),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_138),
.Y(n_189)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_130),
.A2(n_53),
.B1(n_46),
.B2(n_44),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_198),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_201),
.C(n_213),
.Y(n_222)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_158),
.B1(n_132),
.B2(n_156),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_206),
.B1(n_212),
.B2(n_220),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_30),
.B1(n_24),
.B2(n_136),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_219),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_163),
.B(n_40),
.CI(n_46),
.CON(n_208),
.SN(n_208)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_187),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_24),
.B1(n_26),
.B2(n_136),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_24),
.B1(n_136),
.B2(n_40),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_162),
.B(n_67),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_24),
.C(n_26),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_218),
.C(n_181),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_26),
.B(n_1),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_3),
.B(n_5),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_8),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_26),
.C(n_2),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_167),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_169),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_237),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_180),
.B(n_173),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_238),
.B(n_244),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_196),
.B(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_231),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_174),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_230),
.B(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_240),
.C(n_218),
.Y(n_257)
);

OAI21x1_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_190),
.B(n_170),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_209),
.B(n_216),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_160),
.B1(n_172),
.B2(n_173),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_244),
.B1(n_221),
.B2(n_231),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_164),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_192),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_239),
.Y(n_258)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_164),
.C(n_4),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_205),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_246),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_245),
.B1(n_194),
.B2(n_199),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_234),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_5),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_213),
.CI(n_201),
.CON(n_250),
.SN(n_250)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_251),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_194),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_260),
.B(n_9),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_224),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_262),
.C(n_267),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_197),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_9),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_215),
.C(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_208),
.B1(n_211),
.B2(n_6),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_246),
.B1(n_221),
.B2(n_242),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_8),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_3),
.C(n_5),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_273),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_228),
.C(n_236),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.C(n_283),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_226),
.C(n_239),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_250),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_258),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_237),
.B1(n_243),
.B2(n_7),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_254),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_6),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_280),
.Y(n_295)
);

FAx1_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_6),
.CI(n_7),
.CON(n_281),
.SN(n_281)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_256),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_259),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_6),
.C(n_7),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_267),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_294),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_290),
.B(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_249),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_250),
.C(n_261),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_297),
.C(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_255),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_283),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_269),
.B1(n_248),
.B2(n_284),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_272),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_306),
.C(n_309),
.Y(n_311)
);

OR2x6_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_281),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_288),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_268),
.B1(n_259),
.B2(n_271),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_268),
.C(n_282),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_9),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_14),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_315),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_287),
.B(n_7),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_319),
.Y(n_320)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_11),
.A3(n_12),
.B1(n_14),
.B2(n_302),
.C1(n_301),
.C2(n_308),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_312),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_304),
.A2(n_305),
.B(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_11),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_12),
.Y(n_321)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_12),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_324),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_311),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_322),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_320),
.B(n_327),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_326),
.Y(n_332)
);


endmodule