module fake_jpeg_2901_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_27),
.C(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_14),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_55),
.Y(n_90)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_12),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_36),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_28),
.Y(n_61)
);

CKINVDCx9p33_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_66),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_68),
.B(n_75),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_83),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_77),
.B1(n_27),
.B2(n_28),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_25),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_72),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_78),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_20),
.B1(n_32),
.B2(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_21),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_101),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_31),
.B(n_19),
.C(n_21),
.Y(n_83)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_17),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_45),
.B(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_34),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_128),
.B1(n_146),
.B2(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_37),
.B1(n_32),
.B2(n_22),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_133),
.B1(n_71),
.B2(n_79),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_28),
.A3(n_31),
.B1(n_30),
.B2(n_37),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_131),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_37),
.B1(n_40),
.B2(n_39),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_128),
.A2(n_141),
.B1(n_118),
.B2(n_132),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_69),
.A2(n_40),
.B1(n_39),
.B2(n_22),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_129),
.A2(n_142),
.B1(n_148),
.B2(n_111),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_28),
.A3(n_27),
.B1(n_35),
.B2(n_39),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_39),
.B1(n_28),
.B2(n_35),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_73),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_145),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_70),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_149),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_96),
.C(n_98),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_153),
.C(n_154),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_86),
.B1(n_85),
.B2(n_106),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_173),
.B1(n_181),
.B2(n_113),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_74),
.C(n_88),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_74),
.C(n_87),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_76),
.C(n_104),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_107),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_174),
.B1(n_183),
.B2(n_185),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_165),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_65),
.B1(n_70),
.B2(n_76),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_65),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_91),
.CI(n_82),
.CON(n_169),
.SN(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_171),
.B(n_151),
.C(n_153),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_82),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_116),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_85),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_177),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_111),
.B1(n_103),
.B2(n_92),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_103),
.B1(n_92),
.B2(n_3),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_2),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_114),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_136),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_124),
.B1(n_114),
.B2(n_145),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_204),
.B1(n_216),
.B2(n_183),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_159),
.A2(n_124),
.B1(n_113),
.B2(n_119),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_213),
.B1(n_149),
.B2(n_181),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_212),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_201),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_116),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_120),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_208),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_136),
.B1(n_120),
.B2(n_117),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_211),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_117),
.B(n_137),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_162),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_137),
.B1(n_7),
.B2(n_8),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_154),
.A2(n_137),
.B(n_7),
.C(n_8),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_182),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_137),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_6),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_156),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_161),
.C(n_150),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_222),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_161),
.C(n_150),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_191),
.B1(n_205),
.B2(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_245),
.B1(n_188),
.B2(n_193),
.Y(n_252)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_213),
.B1(n_191),
.B2(n_187),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_237),
.B(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_218),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_177),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_195),
.B(n_169),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_198),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_156),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_244),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_174),
.B1(n_168),
.B2(n_175),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_254),
.B1(n_262),
.B2(n_239),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_194),
.B1(n_201),
.B2(n_191),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_250),
.Y(n_274)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_201),
.A3(n_210),
.B1(n_199),
.B2(n_203),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_189),
.B(n_186),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_266),
.B1(n_267),
.B2(n_223),
.Y(n_279)
);

AOI221xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_186),
.B1(n_195),
.B2(n_215),
.C(n_219),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_211),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_228),
.A2(n_198),
.B1(n_204),
.B2(n_207),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_225),
.A2(n_208),
.B1(n_214),
.B2(n_212),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_166),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_263),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_239),
.B1(n_221),
.B2(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_276),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_222),
.C(n_220),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_280),
.C(n_255),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_240),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_277),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_224),
.B1(n_246),
.B2(n_223),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_246),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_232),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_286),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_281),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_226),
.C(n_235),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_238),
.B1(n_234),
.B2(n_233),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_236),
.B1(n_231),
.B2(n_229),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_247),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_229),
.B(n_190),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_266),
.B(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_249),
.B(n_209),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_276),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_295),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_301),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_296),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_281),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_282),
.B1(n_283),
.B2(n_272),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_260),
.C(n_259),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_258),
.C(n_257),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_258),
.C(n_257),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_300),
.B(n_253),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_313),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_271),
.B1(n_279),
.B2(n_274),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_307),
.B1(n_311),
.B2(n_305),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_274),
.B(n_285),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g322 ( 
.A1(n_305),
.A2(n_208),
.A3(n_230),
.B1(n_265),
.B2(n_206),
.C(n_176),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_284),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_291),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_291),
.B1(n_272),
.B2(n_301),
.Y(n_311)
);

OAI221xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_282),
.B1(n_298),
.B2(n_299),
.C(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_300),
.C(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_318),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_310),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_292),
.C(n_253),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_315),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_248),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_320),
.B(n_311),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_265),
.B1(n_208),
.B2(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_325),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_308),
.B(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_308),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_319),
.C(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_330),
.B(n_334),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_329),
.B1(n_317),
.B2(n_206),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_325),
.C(n_316),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.Y(n_338)
);

NAND4xp25_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_332),
.C(n_335),
.D(n_168),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_178),
.C(n_9),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_6),
.Y(n_342)
);


endmodule