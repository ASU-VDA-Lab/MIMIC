module fake_jpeg_26593_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_50),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_15),
.B(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_21),
.B1(n_30),
.B2(n_23),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_48),
.B1(n_41),
.B2(n_32),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_22),
.B1(n_19),
.B2(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_24),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_22),
.B1(n_41),
.B2(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_65),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_72),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_33),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_42),
.B(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_80),
.B1(n_30),
.B2(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_32),
.B1(n_25),
.B2(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_25),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_91),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_59),
.B1(n_49),
.B2(n_60),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_90),
.Y(n_107)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_40),
.C(n_51),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_51),
.C(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_99),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_60),
.B1(n_44),
.B2(n_45),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_68),
.B1(n_72),
.B2(n_82),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_42),
.C(n_60),
.Y(n_99)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_96),
.B1(n_97),
.B2(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_115),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_81),
.B1(n_28),
.B2(n_20),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_28),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_119),
.Y(n_124)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_28),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_87),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_113),
.B(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_132),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_114),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_135),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_93),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_89),
.B(n_84),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_91),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_106),
.C(n_99),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_148),
.C(n_150),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_115),
.C(n_11),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_153),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_106),
.C(n_103),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_106),
.B(n_105),
.C(n_89),
.D(n_94),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_27),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_132),
.C(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_11),
.C(n_14),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_2),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_140),
.C(n_139),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_165),
.C(n_151),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_139),
.B(n_130),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_138),
.A3(n_126),
.B1(n_127),
.B2(n_20),
.C1(n_101),
.C2(n_90),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_127),
.B1(n_116),
.B2(n_111),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_166),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_119),
.C(n_20),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_27),
.B1(n_4),
.B2(n_5),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_146),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_152),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_146),
.CI(n_148),
.CON(n_171),
.SN(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_165),
.C(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_152),
.C(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_163),
.C(n_7),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_6),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_173),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_179),
.C(n_184),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_192),
.B(n_193),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_171),
.B1(n_8),
.B2(n_9),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_169),
.C(n_185),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_177),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_7),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_7),
.B(n_8),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_196),
.A2(n_197),
.B(n_10),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_8),
.B(n_9),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_9),
.Y(n_200)
);


endmodule