module fake_ibex_731_n_909 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_909);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_909;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_375;
wire n_340;
wire n_280;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_35),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_71),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_9),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_67),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_97),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_48),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_63),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_43),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_1),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_125),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_39),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_24),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_53),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_22),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_35),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_55),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_168),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_59),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_109),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_26),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_34),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_R g211 ( 
.A(n_128),
.B(n_150),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_81),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_160),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_56),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_122),
.B(n_83),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_38),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_9),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_44),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_39),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_87),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_12),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_100),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_145),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_105),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_3),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_92),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_91),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_58),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_139),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_143),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_136),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_144),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_66),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_36),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_116),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_45),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_18),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_28),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_90),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_80),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_101),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_46),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_74),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_96),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_114),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_118),
.B(n_112),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_149),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_131),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_174),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_130),
.B(n_64),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_133),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_163),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_164),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_40),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_129),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_2),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_17),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_173),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_84),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_85),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_89),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_134),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_72),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_41),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_94),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_77),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_95),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_42),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_82),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_132),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_23),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_75),
.Y(n_288)
);

BUFx8_ASAP7_75t_SL g289 ( 
.A(n_17),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_124),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_73),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_70),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_152),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_76),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_98),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_31),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_0),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_54),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_140),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_4),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_103),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_78),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_24),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_102),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_93),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_19),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_52),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_31),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_18),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_108),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_12),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_201),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_297),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_205),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_201),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_225),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_254),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_0),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_2),
.Y(n_322)
);

BUFx12f_ASAP7_75t_L g323 ( 
.A(n_189),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_205),
.Y(n_324)
);

BUFx8_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_189),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_194),
.B(n_49),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_203),
.B(n_4),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_189),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_246),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_246),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_289),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_5),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_227),
.B(n_6),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_275),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_200),
.B(n_6),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_180),
.A2(n_88),
.B(n_171),
.Y(n_343)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_180),
.A2(n_86),
.B(n_169),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_207),
.B(n_7),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_252),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_193),
.B(n_307),
.Y(n_347)
);

AOI22x1_ASAP7_75t_SL g348 ( 
.A1(n_179),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_10),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_178),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_282),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_222),
.Y(n_353)
);

BUFx8_ASAP7_75t_SL g354 ( 
.A(n_179),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_211),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_247),
.Y(n_357)
);

BUFx8_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_248),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_176),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_273),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g362 ( 
.A(n_215),
.B(n_50),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_273),
.Y(n_363)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_295),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_243),
.B(n_20),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_186),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_264),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_185),
.A2(n_111),
.B(n_166),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_187),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_267),
.B(n_51),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_271),
.B(n_25),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_197),
.A2(n_113),
.B(n_162),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_279),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_197),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_244),
.B(n_249),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_199),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g380 ( 
.A1(n_199),
.A2(n_110),
.B(n_157),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_218),
.A2(n_107),
.B(n_156),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_284),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_218),
.A2(n_106),
.B(n_155),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_284),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_236),
.B(n_25),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_186),
.A2(n_213),
.B1(n_253),
.B2(n_260),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_236),
.A2(n_104),
.B(n_153),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_241),
.B(n_27),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_241),
.B(n_27),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g391 ( 
.A1(n_259),
.A2(n_117),
.B(n_148),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_259),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_284),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_292),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_270),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_270),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_175),
.Y(n_397)
);

OAI22x1_ASAP7_75t_R g398 ( 
.A1(n_229),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_190),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_192),
.Y(n_400)
);

BUFx12f_ASAP7_75t_L g401 ( 
.A(n_177),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_292),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_182),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_188),
.Y(n_404)
);

CKINVDCx11_ASAP7_75t_R g405 ( 
.A(n_304),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_358),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_326),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g409 ( 
.A(n_397),
.B(n_213),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_358),
.B(n_195),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_358),
.B(n_196),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

CKINVDCx6p67_ASAP7_75t_R g415 ( 
.A(n_323),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_316),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_313),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_340),
.B(n_198),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_316),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_394),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_313),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_362),
.A2(n_223),
.B1(n_308),
.B2(n_301),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_316),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_318),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_209),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

INVx6_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_318),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_357),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_318),
.Y(n_435)
);

OAI22xp33_ASAP7_75t_L g436 ( 
.A1(n_366),
.A2(n_304),
.B1(n_310),
.B2(n_309),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_332),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_365),
.B(n_212),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_342),
.B(n_216),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_314),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_342),
.B(n_217),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_362),
.A2(n_253),
.B1(n_260),
.B2(n_265),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_314),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_351),
.B(n_202),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_342),
.B(n_219),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_331),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_341),
.B(n_257),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_338),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_360),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_347),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_356),
.B(n_226),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_338),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_352),
.B(n_220),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_347),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_356),
.B(n_228),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_324),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_352),
.B(n_237),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_404),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_352),
.B(n_242),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_356),
.B(n_233),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_327),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_403),
.B(n_234),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_377),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_403),
.B(n_235),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_320),
.B(n_258),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_346),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_395),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_377),
.B(n_238),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_320),
.B(n_269),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_346),
.Y(n_475)
);

BUFx6f_ASAP7_75t_SL g476 ( 
.A(n_315),
.Y(n_476)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_328),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_331),
.Y(n_478)
);

INVx8_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

OAI22xp33_ASAP7_75t_L g480 ( 
.A1(n_350),
.A2(n_300),
.B1(n_283),
.B2(n_296),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_317),
.B(n_277),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_319),
.B(n_245),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_337),
.B(n_287),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_328),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_328),
.B(n_181),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g487 ( 
.A(n_322),
.B(n_311),
.C(n_256),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_375),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_379),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_337),
.B(n_183),
.Y(n_490)
);

CKINVDCx9p33_ASAP7_75t_R g491 ( 
.A(n_348),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_335),
.B(n_299),
.C(n_288),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_400),
.B(n_263),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g495 ( 
.A1(n_343),
.A2(n_274),
.B(n_268),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_399),
.B(n_184),
.Y(n_497)
);

AND2x2_ASAP7_75t_SL g498 ( 
.A(n_329),
.B(n_262),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_321),
.B(n_191),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_396),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_361),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_353),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_433),
.B(n_359),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_367),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_448),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_462),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_467),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_374),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_467),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_485),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_429),
.B(n_381),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_440),
.B(n_401),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_469),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_451),
.B(n_387),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_427),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_415),
.B(n_355),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_418),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_442),
.B(n_336),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_426),
.A2(n_265),
.B1(n_272),
.B2(n_210),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_339),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_446),
.B(n_325),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_386),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_406),
.B(n_272),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_444),
.A2(n_371),
.B1(n_345),
.B2(n_305),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_477),
.B(n_370),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_419),
.B(n_389),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_432),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_407),
.A2(n_382),
.B(n_373),
.C(n_368),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_455),
.B(n_459),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_502),
.B(n_390),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_461),
.B(n_484),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_469),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_410),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_L g541 ( 
.A(n_487),
.B(n_470),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_483),
.B(n_206),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_483),
.B(n_208),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_452),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_405),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_499),
.B(n_405),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_408),
.B(n_344),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_490),
.B(n_231),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_414),
.B(n_334),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_456),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_413),
.A2(n_204),
.B1(n_214),
.B2(n_280),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_L g553 ( 
.A(n_480),
.B(n_278),
.C(n_294),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_460),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_456),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_479),
.B(n_334),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_493),
.B(n_306),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_453),
.B(n_224),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_458),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_474),
.A2(n_302),
.B1(n_230),
.B2(n_232),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_457),
.B(n_239),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_481),
.A2(n_240),
.B1(n_250),
.B2(n_255),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_486),
.A2(n_382),
.B(n_380),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_411),
.A2(n_261),
.B1(n_266),
.B2(n_276),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_463),
.B(n_281),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_436),
.B(n_409),
.C(n_412),
.Y(n_566)
);

O2A1O1Ixp33_ASAP7_75t_L g567 ( 
.A1(n_436),
.A2(n_378),
.B(n_385),
.C(n_384),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_473),
.B(n_285),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_494),
.B(n_290),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_478),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_476),
.B(n_291),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_449),
.Y(n_572)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_466),
.B(n_378),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_430),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_438),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_421),
.B(n_298),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_431),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_439),
.B(n_388),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_434),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_434),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_479),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_482),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_449),
.A2(n_378),
.B1(n_385),
.B2(n_391),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_488),
.Y(n_584)
);

NAND2x1_ASAP7_75t_L g585 ( 
.A(n_431),
.B(n_388),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_489),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_479),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_505),
.B(n_464),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_577),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_514),
.B(n_465),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_563),
.A2(n_495),
.B(n_465),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_575),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_585),
.A2(n_495),
.B(n_468),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_570),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_511),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_525),
.B(n_537),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_525),
.B(n_492),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_523),
.B(n_354),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_537),
.B(n_496),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_526),
.B(n_476),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_544),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_572),
.B(n_515),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_522),
.B(n_500),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_472),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_506),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_515),
.B(n_354),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_539),
.B(n_536),
.Y(n_608)
);

AO32x1_ASAP7_75t_L g609 ( 
.A1(n_583),
.A2(n_437),
.A3(n_443),
.B1(n_423),
.B2(n_424),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_527),
.B(n_503),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_550),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_530),
.A2(n_422),
.B1(n_443),
.B2(n_364),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_551),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_532),
.B(n_504),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_509),
.B(n_30),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_555),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_535),
.A2(n_393),
.B(n_383),
.C(n_361),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_530),
.A2(n_398),
.B(n_491),
.C(n_450),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_566),
.A2(n_363),
.B1(n_364),
.B2(n_393),
.Y(n_620)
);

AND3x2_ASAP7_75t_L g621 ( 
.A(n_556),
.B(n_491),
.C(n_38),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_553),
.A2(n_364),
.B1(n_383),
.B2(n_393),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_542),
.B(n_37),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_541),
.B(n_37),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_510),
.Y(n_625)
);

INVx11_ASAP7_75t_L g626 ( 
.A(n_571),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_529),
.B(n_41),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_507),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_517),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_520),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_518),
.A2(n_557),
.B1(n_552),
.B2(n_548),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_558),
.A2(n_501),
.B(n_475),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_543),
.B(n_57),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_545),
.B(n_376),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_519),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_531),
.A2(n_521),
.B(n_524),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_528),
.A2(n_533),
.B(n_540),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_582),
.A2(n_372),
.B(n_471),
.C(n_454),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_508),
.B(n_61),
.Y(n_639)
);

AO21x1_ASAP7_75t_L g640 ( 
.A1(n_584),
.A2(n_62),
.B(n_65),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_577),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_517),
.B(n_454),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_561),
.A2(n_445),
.B(n_441),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_546),
.B(n_68),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

OAI22x1_ASAP7_75t_L g646 ( 
.A1(n_564),
.A2(n_560),
.B1(n_568),
.B2(n_576),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_597),
.A2(n_565),
.B(n_586),
.Y(n_647)
);

INVxp67_ASAP7_75t_SL g648 ( 
.A(n_608),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_593),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_631),
.A2(n_512),
.B1(n_568),
.B2(n_559),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_645),
.B(n_569),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_596),
.B(n_516),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_615),
.B(n_538),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_603),
.B(n_562),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_600),
.B(n_538),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_621),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_611),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_611),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_598),
.B(n_604),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_599),
.B(n_554),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_616),
.A2(n_613),
.B1(n_627),
.B2(n_590),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_628),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_605),
.B(n_573),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_623),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_637),
.B(n_601),
.Y(n_665)
);

AO31x2_ASAP7_75t_L g666 ( 
.A1(n_640),
.A2(n_574),
.A3(n_580),
.B(n_579),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_602),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_612),
.Y(n_668)
);

CKINVDCx14_ASAP7_75t_R g669 ( 
.A(n_630),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_626),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_595),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_595),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_607),
.B(n_119),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_618),
.A2(n_638),
.A3(n_643),
.B(n_632),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_634),
.B(n_172),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_614),
.B(n_141),
.Y(n_676)
);

AND2x2_ASAP7_75t_SL g677 ( 
.A(n_639),
.B(n_146),
.Y(n_677)
);

BUFx6f_ASAP7_75t_SL g678 ( 
.A(n_639),
.Y(n_678)
);

OAI22x1_ASAP7_75t_L g679 ( 
.A1(n_622),
.A2(n_147),
.B1(n_620),
.B2(n_624),
.Y(n_679)
);

NOR2xp67_ASAP7_75t_L g680 ( 
.A(n_646),
.B(n_633),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g681 ( 
.A1(n_609),
.A2(n_642),
.B(n_617),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_606),
.A2(n_625),
.B(n_635),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_589),
.B(n_641),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_588),
.B(n_591),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_629),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_597),
.B(n_610),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_597),
.A2(n_537),
.B(n_567),
.C(n_535),
.Y(n_687)
);

AOI21x1_ASAP7_75t_L g688 ( 
.A1(n_592),
.A2(n_563),
.B(n_547),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_597),
.B(n_610),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_597),
.A2(n_578),
.B(n_594),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_611),
.B(n_444),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_597),
.B(n_610),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_597),
.A2(n_578),
.B(n_594),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_597),
.B(n_511),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_597),
.B(n_610),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_597),
.A2(n_608),
.B1(n_600),
.B2(n_426),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_SL g697 ( 
.A1(n_597),
.A2(n_583),
.B(n_485),
.Y(n_697)
);

AOI21x1_ASAP7_75t_L g698 ( 
.A1(n_592),
.A2(n_563),
.B(n_547),
.Y(n_698)
);

OAI21x1_ASAP7_75t_SL g699 ( 
.A1(n_637),
.A2(n_608),
.B(n_600),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_597),
.B(n_511),
.Y(n_700)
);

NOR4xp25_ASAP7_75t_L g701 ( 
.A(n_619),
.B(n_530),
.C(n_426),
.D(n_567),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_597),
.B(n_511),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_597),
.A2(n_537),
.B(n_567),
.C(n_535),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_596),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_596),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_597),
.A2(n_608),
.B1(n_600),
.B2(n_426),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_597),
.B(n_610),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_597),
.A2(n_537),
.B(n_567),
.C(n_535),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_597),
.A2(n_608),
.B1(n_600),
.B2(n_426),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_596),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_597),
.B(n_610),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_596),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_595),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_596),
.Y(n_714)
);

AO31x2_ASAP7_75t_L g715 ( 
.A1(n_640),
.A2(n_534),
.A3(n_592),
.B(n_636),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g716 ( 
.A1(n_597),
.A2(n_610),
.B(n_631),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_597),
.A2(n_578),
.B(n_594),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_611),
.B(n_444),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_597),
.B(n_505),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_595),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_597),
.B(n_610),
.Y(n_721)
);

NAND2x1p5_ASAP7_75t_L g722 ( 
.A(n_595),
.B(n_581),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_686),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_716),
.B(n_692),
.Y(n_724)
);

CKINVDCx11_ASAP7_75t_R g725 ( 
.A(n_705),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_648),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_695),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_707),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_677),
.B(n_658),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_658),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_716),
.A2(n_709),
.B(n_706),
.C(n_696),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_711),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_720),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_678),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_678),
.A2(n_721),
.B1(n_661),
.B2(n_676),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_691),
.A2(n_718),
.B1(n_654),
.B2(n_665),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_647),
.B(n_649),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_R g738 ( 
.A(n_669),
.B(n_713),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_712),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_661),
.A2(n_676),
.B1(n_664),
.B2(n_650),
.Y(n_740)
);

AO31x2_ASAP7_75t_L g741 ( 
.A1(n_690),
.A2(n_693),
.A3(n_717),
.B(n_679),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_691),
.A2(n_718),
.B1(n_650),
.B2(n_700),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_670),
.B(n_657),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_670),
.B(n_657),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_722),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_680),
.A2(n_675),
.B1(n_655),
.B2(n_697),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_694),
.B(n_702),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_714),
.A2(n_653),
.B1(n_704),
.B2(n_710),
.Y(n_748)
);

INVx4_ASAP7_75t_SL g749 ( 
.A(n_685),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_673),
.B(n_701),
.C(n_660),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_671),
.Y(n_751)
);

OAI21x1_ASAP7_75t_SL g752 ( 
.A1(n_682),
.A2(n_683),
.B(n_684),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_652),
.B(n_651),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_672),
.A2(n_719),
.B1(n_662),
.B2(n_667),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_668),
.B(n_663),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_656),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_681),
.A2(n_685),
.B1(n_715),
.B2(n_674),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_666),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_716),
.B(n_686),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_716),
.B(n_706),
.C(n_696),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

AO21x2_ASAP7_75t_L g762 ( 
.A1(n_699),
.A2(n_698),
.B(n_688),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_686),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_657),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_716),
.A2(n_659),
.B(n_648),
.C(n_687),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_686),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_712),
.Y(n_767)
);

NAND2x1p5_ASAP7_75t_L g768 ( 
.A(n_677),
.B(n_658),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_648),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_677),
.B(n_658),
.Y(n_770)
);

INVx6_ASAP7_75t_L g771 ( 
.A(n_658),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_686),
.B(n_689),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_716),
.A2(n_706),
.B1(n_709),
.B2(n_696),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_694),
.B(n_721),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_686),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_686),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_686),
.B(n_689),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_716),
.B(n_686),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_687),
.A2(n_708),
.B(n_703),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_686),
.B(n_721),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_737),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_726),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_725),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_726),
.B(n_749),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_724),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_723),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_772),
.B(n_777),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_759),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_769),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_771),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_730),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_780),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_762),
.Y(n_793)
);

AOI222xp33_ASAP7_75t_L g794 ( 
.A1(n_780),
.A2(n_774),
.B1(n_747),
.B2(n_766),
.C1(n_727),
.C2(n_728),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_735),
.A2(n_742),
.B1(n_740),
.B2(n_736),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_735),
.A2(n_742),
.B1(n_740),
.B2(n_736),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_729),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_778),
.Y(n_798)
);

INVxp33_ASAP7_75t_L g799 ( 
.A(n_738),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_752),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_739),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_729),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_750),
.A2(n_765),
.B(n_731),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_732),
.B(n_763),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_761),
.B(n_776),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_758),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_758),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_779),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_775),
.B(n_748),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_785),
.B(n_757),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_781),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_782),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_788),
.B(n_760),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_784),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_789),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_789),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_788),
.B(n_760),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_784),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_793),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_795),
.A2(n_768),
.B1(n_770),
.B2(n_773),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_800),
.B(n_741),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_819),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_814),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_821),
.B(n_793),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_811),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_815),
.B(n_806),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_820),
.B(n_792),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_810),
.B(n_798),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_815),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_810),
.B(n_806),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_811),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_816),
.B(n_807),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_813),
.B(n_808),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_810),
.B(n_807),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_816),
.B(n_786),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_822),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_833),
.B(n_812),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_824),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_835),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_833),
.B(n_812),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_825),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_828),
.B(n_813),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_829),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_825),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_828),
.B(n_813),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_830),
.B(n_834),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_831),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_830),
.B(n_817),
.Y(n_848)
);

NOR2x1_ASAP7_75t_SL g849 ( 
.A(n_823),
.B(n_814),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_835),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_834),
.B(n_817),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_839),
.B(n_826),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_846),
.B(n_838),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_836),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_841),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_841),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_850),
.B(n_826),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_837),
.B(n_832),
.Y(n_858)
);

NOR2x1_ASAP7_75t_L g859 ( 
.A(n_837),
.B(n_784),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_840),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_844),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_838),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_846),
.B(n_824),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_838),
.B(n_824),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_858),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_862),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_SL g867 ( 
.A(n_860),
.B(n_770),
.C(n_768),
.Y(n_867)
);

AOI321xp33_ASAP7_75t_L g868 ( 
.A1(n_859),
.A2(n_827),
.A3(n_820),
.B1(n_796),
.B2(n_843),
.C(n_809),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_858),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_857),
.B(n_840),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_852),
.B(n_842),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_853),
.A2(n_838),
.B1(n_845),
.B2(n_818),
.Y(n_872)
);

AOI33xp33_ASAP7_75t_L g873 ( 
.A1(n_853),
.A2(n_748),
.A3(n_767),
.B1(n_804),
.B2(n_787),
.B3(n_753),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_857),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_852),
.B(n_848),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_863),
.B(n_824),
.Y(n_876)
);

AOI221xp5_ASAP7_75t_L g877 ( 
.A1(n_872),
.A2(n_874),
.B1(n_865),
.B2(n_869),
.C(n_871),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_870),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_867),
.Y(n_879)
);

OAI221xp5_ASAP7_75t_L g880 ( 
.A1(n_868),
.A2(n_862),
.B1(n_851),
.B2(n_861),
.C(n_803),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_876),
.A2(n_864),
.B1(n_863),
.B2(n_862),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_875),
.B(n_854),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_866),
.A2(n_799),
.B(n_794),
.C(n_801),
.Y(n_883)
);

AOI21xp33_ASAP7_75t_L g884 ( 
.A1(n_879),
.A2(n_756),
.B(n_734),
.Y(n_884)
);

OAI221xp5_ASAP7_75t_SL g885 ( 
.A1(n_877),
.A2(n_873),
.B1(n_866),
.B2(n_864),
.C(n_876),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_883),
.B(n_783),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_878),
.B(n_880),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_SL g888 ( 
.A(n_881),
.B(n_873),
.C(n_802),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_882),
.B(n_855),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_889),
.Y(n_890)
);

NAND2xp33_ASAP7_75t_L g891 ( 
.A(n_887),
.B(n_734),
.Y(n_891)
);

XNOR2x1_ASAP7_75t_L g892 ( 
.A(n_886),
.B(n_866),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_888),
.Y(n_893)
);

AOI211xp5_ASAP7_75t_L g894 ( 
.A1(n_893),
.A2(n_885),
.B(n_884),
.C(n_746),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_891),
.A2(n_849),
.B(n_802),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_890),
.Y(n_896)
);

AOI211x1_ASAP7_75t_L g897 ( 
.A1(n_891),
.A2(n_855),
.B(n_856),
.C(n_847),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_894),
.B(n_892),
.Y(n_898)
);

OAI211xp5_ASAP7_75t_SL g899 ( 
.A1(n_896),
.A2(n_767),
.B(n_754),
.C(n_764),
.Y(n_899)
);

XNOR2xp5_ASAP7_75t_L g900 ( 
.A(n_898),
.B(n_895),
.Y(n_900)
);

AND2x2_ASAP7_75t_SL g901 ( 
.A(n_899),
.B(n_743),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_901),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_902),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_903),
.B(n_900),
.C(n_902),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_904),
.A2(n_901),
.B1(n_744),
.B2(n_743),
.Y(n_905)
);

OAI322xp33_ASAP7_75t_L g906 ( 
.A1(n_905),
.A2(n_897),
.A3(n_745),
.B1(n_755),
.B2(n_764),
.C1(n_790),
.C2(n_805),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_906),
.A2(n_744),
.B(n_733),
.Y(n_907)
);

OR2x6_ASAP7_75t_L g908 ( 
.A(n_907),
.B(n_751),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_908),
.A2(n_771),
.B1(n_797),
.B2(n_791),
.Y(n_909)
);


endmodule