module fake_jpeg_7747_n_170 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_3),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_27),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx6p67_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_13),
.B1(n_23),
.B2(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_17),
.B1(n_22),
.B2(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_53),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_63),
.B1(n_24),
.B2(n_36),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_0),
.C(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_65),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_26),
.B(n_27),
.C(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_12),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_58),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_15),
.B(n_30),
.C(n_19),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_61),
.B(n_62),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_12),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_0),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_76),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_27),
.C(n_40),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_83),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_0),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_14),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_17),
.B(n_14),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_65),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_46),
.B1(n_56),
.B2(n_40),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_102),
.B1(n_69),
.B2(n_82),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_32),
.B1(n_59),
.B2(n_29),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_66),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_108),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_44),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_77),
.Y(n_115)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_69),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_77),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_83),
.B(n_84),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_118),
.B1(n_100),
.B2(n_108),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_84),
.B(n_44),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_93),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_124),
.B1(n_90),
.B2(n_92),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_105),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_95),
.C(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_76),
.B1(n_75),
.B2(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.C(n_136),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_109),
.C(n_70),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_130),
.B1(n_121),
.B2(n_114),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_114),
.B(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_106),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_28),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_88),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_110),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_112),
.C(n_86),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_141),
.B1(n_143),
.B2(n_136),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_64),
.B(n_57),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_116),
.B1(n_118),
.B2(n_111),
.Y(n_141)
);

AOI211xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_123),
.B(n_120),
.C(n_75),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_147),
.C(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_73),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_151),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_140),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_120),
.B(n_134),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_28),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_14),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_57),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_146),
.B(n_143),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_3),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_159),
.B1(n_4),
.B2(n_5),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_147),
.B1(n_29),
.B2(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

OAI221xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_14),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_4),
.B(n_8),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_166),
.B(n_161),
.C(n_159),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_167),
.B1(n_9),
.B2(n_8),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_169),
.Y(n_170)
);


endmodule