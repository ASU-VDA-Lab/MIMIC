module fake_jpeg_28057_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_69),
.Y(n_80)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_49),
.B1(n_41),
.B2(n_60),
.Y(n_92)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_50),
.B1(n_61),
.B2(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_58),
.B1(n_47),
.B2(n_46),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_57),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_82),
.Y(n_96)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_89),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_53),
.B1(n_60),
.B2(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_93),
.Y(n_108)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_43),
.B1(n_49),
.B2(n_45),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_41),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_106),
.A2(n_70),
.B1(n_96),
.B2(n_80),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_114),
.B1(n_9),
.B2(n_10),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_86),
.B1(n_93),
.B2(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_117),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_102),
.C(n_81),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_5),
.C(n_6),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_75),
.B1(n_81),
.B2(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_4),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_97),
.B1(n_98),
.B2(n_3),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_103),
.B(n_101),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_19),
.B(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_0),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_132),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_129),
.B(n_32),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_27),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_128),
.C(n_29),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_30),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_16),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_5),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_133),
.B1(n_17),
.B2(n_18),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_137),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_136),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_134),
.C(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_138),
.C(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_145),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_143),
.C(n_119),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_140),
.A3(n_141),
.B1(n_121),
.B2(n_129),
.C1(n_120),
.C2(n_139),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

AOI321xp33_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_140),
.A3(n_33),
.B1(n_35),
.B2(n_36),
.C(n_37),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_153),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);


endmodule