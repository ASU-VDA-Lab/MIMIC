module real_aes_4930_n_13 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_13);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_13;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_16;
wire n_37;
wire n_35;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_0), .Y(n_24) );
AOI322xp5_ASAP7_75t_SL g13 ( .A1(n_1), .A2(n_6), .A3(n_14), .B1(n_15), .B2(n_25), .C1(n_32), .C2(n_37), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_2), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g31 ( .A(n_2), .B(n_5), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_3), .B(n_18), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_4), .B(n_17), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_4), .Y(n_30) );
NOR4xp25_ASAP7_75t_SL g40 ( .A(n_4), .B(n_23), .C(n_24), .D(n_41), .Y(n_40) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_5), .Y(n_14) );
NAND3xp33_ASAP7_75t_SL g18 ( .A(n_7), .B(n_19), .C(n_20), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g22 ( .A(n_8), .B(n_9), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g27 ( .A(n_8), .B(n_28), .C(n_29), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_9), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_10), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_11), .Y(n_20) );
BUFx8_ASAP7_75t_SL g36 ( .A(n_12), .Y(n_36) );
NAND2xp33_ASAP7_75t_R g39 ( .A(n_14), .B(n_40), .Y(n_39) );
NOR4xp25_ASAP7_75t_SL g15 ( .A(n_16), .B(n_21), .C(n_23), .D(n_24), .Y(n_15) );
NAND3xp33_ASAP7_75t_SL g29 ( .A(n_17), .B(n_24), .C(n_30), .Y(n_29) );
NAND2xp33_ASAP7_75t_R g41 ( .A(n_17), .B(n_22), .Y(n_41) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_26), .Y(n_25) );
NAND2xp33_ASAP7_75t_R g26 ( .A(n_27), .B(n_31), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g34 ( .A(n_35), .Y(n_34) );
CKINVDCx20_ASAP7_75t_R g35 ( .A(n_36), .Y(n_35) );
HB1xp67_ASAP7_75t_L g37 ( .A(n_38), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g38 ( .A(n_39), .Y(n_38) );
endmodule