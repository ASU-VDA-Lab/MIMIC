module real_jpeg_20940_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g11 ( 
.A1(n_1),
.A2(n_2),
.B1(n_12),
.B2(n_13),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_15),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_4),
.B1(n_13),
.B2(n_19),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g27 ( 
.A1(n_1),
.A2(n_2),
.B(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_5),
.B1(n_12),
.B2(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_2),
.B(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_5),
.B1(n_32),
.B2(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_5),
.B1(n_19),
.B2(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_12),
.B(n_19),
.C(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_37),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_24),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_20),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_17),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_10),
.B(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_36),
.B1(n_41),
.B2(n_46),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_14),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_12),
.B(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_35),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_47),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);


endmodule