module real_jpeg_18975_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_1),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_1),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_1),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_1),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_1),
.B(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_3),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_3),
.Y(n_313)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_3),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_4),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_4),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_5),
.B(n_104),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_5),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_5),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_5),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_5),
.B(n_450),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_5),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_5),
.B(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_5),
.B(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_6),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_6),
.B(n_88),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_6),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_6),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_6),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_6),
.B(n_424),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_6),
.B(n_508),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_7),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_7),
.B(n_64),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_7),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_7),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_7),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_7),
.B(n_219),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_8),
.Y(n_101)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g457 ( 
.A(n_8),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_9),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_9),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_9),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_9),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_9),
.A2(n_10),
.B1(n_287),
.B2(n_292),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_10),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_10),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g306 ( 
.A(n_10),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_10),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_10),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_10),
.B(n_498),
.Y(n_497)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_11),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_11),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_12),
.B(n_120),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_12),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g308 ( 
.A(n_12),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g311 ( 
.A(n_12),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_12),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_12),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_12),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_12),
.B(n_457),
.Y(n_456)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_13),
.Y(n_320)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_14),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_14),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_14),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_14),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_14),
.B(n_349),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g462 ( 
.A(n_16),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_16),
.Y(n_496)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_17),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_17),
.Y(n_178)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_259),
.B(n_528),
.C(n_535),
.D(n_537),
.Y(n_21)
);

NOR3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_229),
.C(n_249),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_182),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_25),
.A2(n_531),
.B(n_532),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_147),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_26),
.B(n_147),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_109),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_27),
.B(n_110),
.C(n_123),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_77),
.C(n_92),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_29),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_48),
.C(n_62),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_30),
.B(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_32),
.A2(n_40),
.B1(n_113),
.B2(n_117),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_32),
.B(n_41),
.C(n_42),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_32),
.B(n_306),
.C(n_308),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_32),
.A2(n_40),
.B1(n_306),
.B2(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_34),
.Y(n_349)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_35),
.Y(n_482)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_36),
.B(n_95),
.C(n_99),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_36),
.A2(n_41),
.B1(n_99),
.B2(n_100),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_36),
.B(n_218),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_36),
.B(n_358),
.Y(n_421)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_40),
.B(n_113),
.C(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_43),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_43),
.B(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_44),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_45),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_46),
.Y(n_346)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_48),
.B(n_62),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_59),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_168)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_52),
.Y(n_309)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_52),
.Y(n_480)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_59),
.A2(n_60),
.B1(n_113),
.B2(n_117),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_60),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_60),
.B(n_113),
.C(n_294),
.Y(n_351)
);

XNOR2x1_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_63),
.B(n_71),
.C(n_75),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_63),
.B(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_63),
.B(n_137),
.C(n_224),
.Y(n_252)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_65),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_71),
.A2(n_76),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_74),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_76),
.B(n_137),
.C(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_77),
.B(n_92),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_87),
.B2(n_91),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_83),
.C(n_87),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_81),
.B(n_171),
.C(n_175),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_81),
.B(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_86),
.Y(n_282)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_87),
.A2(n_91),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_87),
.B(n_225),
.C(n_255),
.Y(n_536)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_105),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g179 ( 
.A1(n_93),
.A2(n_94),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_95),
.A2(n_224),
.B1(n_225),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_95),
.Y(n_255)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_158),
.C(n_162),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_99),
.A2(n_100),
.B1(n_162),
.B2(n_163),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_99),
.B(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_100),
.B(n_428),
.Y(n_464)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_101),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_101),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_102),
.A2(n_252),
.B(n_536),
.Y(n_537)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_104),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_106),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_170),
.C(n_176),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_106),
.A2(n_107),
.B1(n_176),
.B2(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_106),
.B(n_140),
.C(n_143),
.Y(n_234)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_123),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.C(n_122),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_113),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_117),
.B1(n_133),
.B2(n_137),
.Y(n_132)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_117),
.B(n_133),
.C(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_138),
.B2(n_139),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_126),
.B(n_127),
.C(n_138),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_128),
.Y(n_243)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_133),
.A2(n_137),
.B1(n_224),
.B2(n_225),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_133),
.A2(n_137),
.B1(n_198),
.B2(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_136),
.Y(n_307)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_152),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_150),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_169),
.C(n_179),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_154),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_167),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_155),
.B(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_157),
.B(n_167),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_159),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_159),
.B(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_162),
.A2(n_163),
.B1(n_301),
.B2(n_302),
.Y(n_325)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_163),
.B(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_164),
.Y(n_317)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_179),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

OR2x6_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_183),
.B(n_185),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_192),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_186),
.B(n_189),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_192),
.B(n_409),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_205),
.C(n_210),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_193),
.A2(n_194),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_202),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_195),
.B(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_197),
.A2(n_202),
.B1(n_203),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_197),
.Y(n_386)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_198),
.Y(n_341)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_398)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.C(n_224),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_212),
.A2(n_213),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_214),
.A2(n_218),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_214),
.Y(n_357)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_215),
.Y(n_430)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_217),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_218),
.Y(n_358)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_220),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_223),
.Y(n_426)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_226),
.Y(n_378)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

A2O1A1O1Ixp25_ASAP7_75t_L g529 ( 
.A1(n_230),
.A2(n_250),
.B(n_530),
.C(n_533),
.D(n_534),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_248),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_231),
.B(n_248),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_234),
.C(n_247),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_246),
.B2(n_247),
.Y(n_233)
);

CKINVDCx12_ASAP7_75t_R g246 ( 
.A(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_242),
.C(n_244),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_239),
.Y(n_244)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_251),
.B(n_258),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_251),
.Y(n_538)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.CI(n_257),
.CON(n_251),
.SN(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

NAND2x1_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_411),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_388),
.B(n_404),
.C(n_405),
.D(n_410),
.Y(n_260)
);

OAI21x1_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_364),
.B(n_387),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_335),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g527 ( 
.A(n_263),
.B(n_335),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_296),
.C(n_321),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_264),
.B(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_276),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_265),
.B(n_277),
.C(n_293),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.C(n_271),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_266),
.B(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_267),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_419)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_293),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_283),
.B(n_286),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_286),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_296),
.A2(n_297),
.B1(n_321),
.B2(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_310),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_304),
.B2(n_305),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_305),
.C(n_310),
.Y(n_352)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_306),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_311),
.B(n_315),
.C(n_318),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_321),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.C(n_326),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_322),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_325),
.B(n_326),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.C(n_333),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_327),
.B(n_333),
.Y(n_469)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_330),
.B(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_353),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_354),
.C(n_363),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_352),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_347),
.B1(n_348),
.B2(n_350),
.Y(n_343)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_348),
.B(n_351),
.C(n_380),
.Y(n_379)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_350),
.Y(n_380)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_368),
.C(n_369),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_363),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_361),
.C(n_362),
.Y(n_373)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_360),
.Y(n_362)
);

NOR2x1_ASAP7_75t_L g526 ( 
.A(n_364),
.B(n_527),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_366),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_390),
.C(n_391),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_383),
.B2(n_384),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_374)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_375),
.Y(n_381)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_394),
.C(n_395),
.Y(n_393)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_384),
.Y(n_391)
);

NAND4xp25_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_405),
.C(n_412),
.D(n_526),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_392),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_393),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_400),
.B1(n_402),
.B2(n_403),
.Y(n_396)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_397),
.Y(n_402)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_398),
.Y(n_399)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_400),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_402),
.C(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_406),
.B(n_408),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_434),
.B(n_525),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_431),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_414),
.B(n_431),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_418),
.C(n_420),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_415),
.A2(n_416),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_418),
.B(n_420),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.C(n_427),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_421),
.A2(n_422),
.B1(n_423),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_421),
.Y(n_472)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_427),
.B(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_519),
.B(n_524),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_473),
.B(n_518),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_465),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_437),
.B(n_465),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_454),
.C(n_463),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_438),
.A2(n_439),
.B1(n_484),
.B2(n_486),
.Y(n_483)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_449),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_447),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_447),
.C(n_449),
.Y(n_467)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_454),
.A2(n_463),
.B1(n_464),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_476)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_470),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_467),
.B(n_468),
.C(n_470),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_487),
.B(n_517),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_483),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_475),
.B(n_483),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.C(n_481),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_500),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_477),
.A2(n_478),
.B1(n_481),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_481),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_484),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_488),
.A2(n_502),
.B(n_516),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_499),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_489),
.B(n_499),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_497),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_497),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_506),
.B(n_515),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_505),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_504),
.B(n_505),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_510),
.Y(n_506)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_521),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_520),
.B(n_521),
.Y(n_524)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_536),
.Y(n_535)
);


endmodule