module fake_jpeg_10499_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_32),
.B1(n_17),
.B2(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_55),
.B1(n_64),
.B2(n_17),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_31),
.B1(n_27),
.B2(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_100)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_38),
.B1(n_43),
.B2(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_59),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_38),
.B1(n_43),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_83),
.B1(n_33),
.B2(n_28),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_36),
.C(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_86),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_36),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_28),
.B(n_1),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_17),
.B1(n_21),
.B2(n_30),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_19),
.B1(n_21),
.B2(n_30),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_19),
.B1(n_29),
.B2(n_22),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_58),
.B1(n_43),
.B2(n_19),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_84),
.B1(n_100),
.B2(n_33),
.Y(n_114)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_91),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_37),
.C(n_42),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_22),
.B(n_29),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_97),
.B(n_1),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_0),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_0),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_96),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_24),
.B1(n_65),
.B2(n_37),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_42),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_114),
.B1(n_72),
.B2(n_69),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_109),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_40),
.Y(n_109)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_116),
.B1(n_124),
.B2(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_119),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_126),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_73),
.B1(n_74),
.B2(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_87),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_70),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_75),
.C(n_86),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_151),
.C(n_5),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_2),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_137),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_120),
.B(n_104),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_70),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_95),
.B1(n_96),
.B2(n_71),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_141),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_102),
.B(n_101),
.C(n_109),
.D(n_106),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_118),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_148),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_111),
.B1(n_102),
.B2(n_112),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_71),
.B1(n_85),
.B2(n_94),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_85),
.B1(n_97),
.B2(n_82),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_107),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_105),
.A3(n_97),
.B1(n_119),
.B2(n_113),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_104),
.B(n_6),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_153),
.B1(n_134),
.B2(n_147),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_89),
.C(n_90),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_89),
.B1(n_15),
.B2(n_4),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_5),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_131),
.Y(n_187)
);

NAND2x1_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_104),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_161),
.B(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_167),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_3),
.B(n_4),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_166),
.B1(n_158),
.B2(n_169),
.C(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_175),
.B1(n_159),
.B2(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_170),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_104),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_103),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_172),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.C(n_176),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_5),
.C(n_6),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_143),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_6),
.C(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_186),
.B(n_191),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_185),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_148),
.C(n_142),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_164),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_195),
.B1(n_164),
.B2(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_137),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_140),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_173),
.C(n_174),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_145),
.B1(n_129),
.B2(n_151),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_167),
.B(n_155),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_204),
.B(n_210),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_203),
.C(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_206),
.B1(n_8),
.B2(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_8),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

NAND3xp33_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_179),
.C(n_180),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_217),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_200),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_213),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_208),
.A2(n_195),
.A3(n_192),
.B1(n_181),
.B2(n_182),
.C1(n_194),
.C2(n_177),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_219),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_177),
.C(n_138),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_220),
.C(n_201),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_13),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_209),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_11),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_210),
.B(n_12),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_224),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_208),
.B1(n_199),
.B2(n_197),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_204),
.B1(n_213),
.B2(n_220),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_199),
.C(n_197),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_212),
.B(n_11),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_219),
.C(n_13),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_216),
.B1(n_228),
.B2(n_224),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_235),
.B(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_13),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_223),
.Y(n_241)
);

NOR4xp25_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_242),
.C(n_234),
.D(n_232),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_229),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_247),
.B(n_238),
.CI(n_236),
.CON(n_248),
.SN(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_229),
.B1(n_246),
.B2(n_238),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_248),
.Y(n_250)
);


endmodule