module fake_jpeg_25841_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx2_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_17),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_81),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_62),
.B1(n_55),
.B2(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_54),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_58),
.B1(n_64),
.B2(n_53),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_55),
.B1(n_49),
.B2(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_74),
.B1(n_70),
.B2(n_63),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_69),
.B(n_67),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_60),
.B(n_56),
.C(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_102),
.B1(n_90),
.B2(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_105),
.Y(n_111)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_64),
.B1(n_71),
.B2(n_51),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_60),
.B(n_73),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_106),
.B(n_108),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_61),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_61),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_107),
.A2(n_93),
.B1(n_89),
.B2(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_0),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_94),
.B1(n_93),
.B2(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_119),
.B1(n_95),
.B2(n_2),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_118),
.B1(n_97),
.B2(n_96),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_87),
.B(n_24),
.C(n_26),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_20),
.B1(n_46),
.B2(n_45),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_19),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_47),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_101),
.B(n_102),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_130),
.B(n_131),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_128),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_127),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_23),
.C(n_43),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_120),
.C(n_3),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

AND2x4_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_109),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_138),
.B1(n_143),
.B2(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_140),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_111),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_139),
.B(n_142),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_112),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_1),
.B(n_5),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_148),
.B(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_141),
.B1(n_134),
.B2(n_135),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_156),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_148),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_157),
.A3(n_134),
.B1(n_147),
.B2(n_155),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_150),
.B1(n_152),
.B2(n_142),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_35),
.A3(n_34),
.B1(n_33),
.B2(n_31),
.C(n_30),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_28),
.A3(n_27),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_7),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_8),
.B(n_9),
.Y(n_165)
);

OAI31xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_10),
.A3(n_13),
.B(n_14),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_16),
.Y(n_167)
);


endmodule