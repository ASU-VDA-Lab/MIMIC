module fake_jpeg_16754_n_271 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_18),
.B1(n_31),
.B2(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_20),
.B1(n_22),
.B2(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_30),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_27),
.C(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_63),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_60),
.B1(n_61),
.B2(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_19),
.B1(n_21),
.B2(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_32),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_71),
.Y(n_95)
);

OR2x4_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_27),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_55),
.B(n_47),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_16),
.B1(n_24),
.B2(n_25),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_17),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_77),
.B1(n_51),
.B2(n_54),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_33),
.B1(n_38),
.B2(n_35),
.Y(n_77)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_33),
.B1(n_38),
.B2(n_35),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_83),
.B1(n_54),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_38),
.B1(n_16),
.B2(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_24),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_112),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_65),
.B(n_0),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_106),
.B(n_27),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_51),
.B1(n_54),
.B2(n_38),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_70),
.B1(n_89),
.B2(n_77),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_56),
.B1(n_40),
.B2(n_39),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_20),
.B(n_22),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_115),
.B(n_71),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_1),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_40),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_117),
.B(n_128),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_69),
.C(n_80),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_69),
.B1(n_79),
.B2(n_90),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_135),
.B1(n_114),
.B2(n_108),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_86),
.B1(n_56),
.B2(n_80),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_108),
.B1(n_96),
.B2(n_113),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_88),
.C(n_27),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_132),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_92),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_64),
.B1(n_57),
.B2(n_49),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_25),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_2),
.B(n_4),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_4),
.B(n_5),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_155),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_149),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_157),
.B1(n_159),
.B2(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_95),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_123),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_158),
.Y(n_171)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_106),
.B1(n_98),
.B2(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_105),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_104),
.B1(n_64),
.B2(n_57),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_160),
.A2(n_162),
.B(n_138),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_27),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_102),
.B(n_109),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_155),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_116),
.B(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_183),
.B1(n_174),
.B2(n_162),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_120),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_181),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_144),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_177),
.B1(n_180),
.B2(n_185),
.Y(n_194)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_182),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_131),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_151),
.Y(n_192)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_152),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_141),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_121),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_143),
.B1(n_157),
.B2(n_133),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_201),
.B1(n_204),
.B2(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_202),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_168),
.B1(n_176),
.B2(n_117),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_177),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_150),
.C(n_161),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_178),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_156),
.C(n_131),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_124),
.C(n_163),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_159),
.C(n_130),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_126),
.B1(n_160),
.B2(n_119),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_102),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_102),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_73),
.C(n_57),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_166),
.B1(n_164),
.B2(n_182),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_213),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_169),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_219),
.C(n_205),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_167),
.B(n_170),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_221),
.B(n_109),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_166),
.B1(n_180),
.B2(n_177),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_216),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_184),
.B(n_165),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_165),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_195),
.C(n_203),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_226),
.C(n_227),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_186),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_192),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_165),
.C(n_198),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_16),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_25),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_237),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_238),
.B(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_214),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_218),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_210),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_218),
.B1(n_210),
.B2(n_217),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_6),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_243),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_223),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_248),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_24),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_222),
.C(n_229),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_234),
.C(n_16),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_49),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_23),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_8),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_6),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_258),
.A3(n_253),
.B1(n_246),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_247),
.B(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_259),
.B(n_8),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_264),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_9),
.Y(n_265)
);

AOI31xp67_ASAP7_75t_SL g264 ( 
.A1(n_254),
.A2(n_9),
.A3(n_10),
.B(n_12),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_267),
.B(n_262),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_23),
.C(n_14),
.Y(n_267)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_14),
.B(n_15),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_268),
.Y(n_271)
);


endmodule