module fake_jpeg_7336_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_38),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_19),
.B1(n_23),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_49),
.B1(n_15),
.B2(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_33),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_19),
.B1(n_23),
.B2(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_56),
.Y(n_85)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_63),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_25),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_32),
.B(n_1),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_68),
.B(n_77),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_67),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_15),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_16),
.B1(n_20),
.B2(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_78),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_16),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_27),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_61),
.B1(n_69),
.B2(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_68),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_11),
.C(n_12),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_103),
.B(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_72),
.C(n_59),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_91),
.C(n_100),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_106),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_13),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_113),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_97),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_0),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_66),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_87),
.B1(n_98),
.B2(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_87),
.B(n_12),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_66),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_130),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_132),
.C(n_118),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_84),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_24),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_87),
.B1(n_82),
.B2(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_129),
.A2(n_101),
.B1(n_112),
.B2(n_103),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_87),
.C(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_105),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_140),
.C(n_120),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_139),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_143),
.B1(n_137),
.B2(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_102),
.C(n_93),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_132),
.B(n_83),
.CI(n_62),
.CON(n_141),
.SN(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_126),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_144),
.B1(n_131),
.B2(n_95),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_121),
.B(n_127),
.C(n_129),
.D(n_123),
.Y(n_143)
);

OAI321xp33_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_83),
.A3(n_62),
.B1(n_24),
.B2(n_9),
.C(n_10),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_122),
.C(n_140),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_131),
.C(n_121),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_141),
.B1(n_143),
.B2(n_24),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_104),
.C(n_80),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_55),
.B1(n_24),
.B2(n_34),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_158),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_147),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_141),
.B1(n_11),
.B2(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_153),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_157),
.C(n_160),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_166),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_0),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_2),
.C(n_3),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_37),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_2),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_4),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_173),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_167),
.B(n_6),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);


endmodule