module real_jpeg_11123_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_11, n_14, n_344, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_11;
input n_14;
input n_344;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_1),
.A2(n_34),
.B1(n_65),
.B2(n_68),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_12),
.B(n_32),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_3),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_3),
.A2(n_128),
.B(n_154),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_8),
.A2(n_65),
.B1(n_68),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_8),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_107),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_107),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_107),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_65),
.B1(n_68),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_9),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_156),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_156),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_156),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_11),
.A2(n_57),
.B1(n_65),
.B2(n_68),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_277)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_48),
.B(n_60),
.C(n_87),
.D(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_12),
.B(n_46),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_12),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_12),
.A2(n_108),
.B(n_110),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_12),
.A2(n_31),
.B(n_42),
.C(n_144),
.D(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_12),
.B(n_31),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_12),
.B(n_35),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_125),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_13),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_13),
.A2(n_65),
.B1(n_68),
.B2(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_13),
.A2(n_23),
.B1(n_25),
.B2(n_90),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_14),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_22),
.B1(n_65),
.B2(n_68),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_14),
.A2(n_22),
.B1(n_47),
.B2(n_48),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_23),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_15),
.A2(n_55),
.B1(n_65),
.B2(n_68),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_16),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_16),
.A2(n_65),
.B1(n_68),
.B2(n_102),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_102),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_16),
.A2(n_23),
.B1(n_25),
.B2(n_102),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_337),
.B(n_340),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_76),
.B(n_336),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_20),
.B(n_36),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_20),
.B(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_20),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_23),
.A2(n_28),
.B(n_125),
.C(n_187),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_26),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_26),
.B(n_206),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_339)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_27),
.A2(n_30),
.B1(n_220),
.B2(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_27),
.A2(n_205),
.B(n_243),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_286),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_30),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_30),
.A2(n_221),
.B(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_35),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_71),
.C(n_73),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_37),
.A2(n_38),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_311),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_41),
.A2(n_50),
.B1(n_165),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_41),
.A2(n_200),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_46),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_42),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_42),
.A2(n_46),
.B1(n_240),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_42),
.A2(n_46),
.B1(n_258),
.B2(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_44),
.B(n_47),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_45),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_48),
.A2(n_144),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_50),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_50),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_50),
.A2(n_166),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_52),
.A2(n_53),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_58),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_58),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_59),
.A2(n_69),
.B1(n_101),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_59),
.A2(n_142),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_59),
.A2(n_69),
.B1(n_197),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_59),
.A2(n_69),
.B1(n_215),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_59),
.A2(n_69),
.B1(n_234),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_60),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_60),
.A2(n_64),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_68),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_68),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_65),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_109),
.Y(n_108)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_68),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_69),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_69),
.A2(n_103),
.B(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_70),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_71),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_329),
.B(n_335),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_302),
.A3(n_322),
.B1(n_327),
.B2(n_328),
.C(n_344),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_250),
.A3(n_290),
.B1(n_296),
.B2(n_301),
.C(n_345),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_208),
.C(n_247),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_180),
.B(n_207),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_159),
.B(n_179),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_136),
.B(n_158),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_113),
.B(n_135),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_95),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_112),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_108),
.A2(n_109),
.B1(n_155),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_108),
.A2(n_109),
.B1(n_170),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_108),
.A2(n_109),
.B1(n_190),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_108),
.A2(n_109),
.B1(n_213),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_108),
.A2(n_109),
.B(n_232),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_117),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_125),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_122),
.B(n_134),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_120),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_129),
.B(n_133),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_126),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_138),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_149),
.B2(n_157),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_148),
.C(n_157),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_175),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_176),
.C(n_177),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_174),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_171),
.C(n_172),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_182),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_194),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_193),
.C(n_194),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_189),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_209),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_227),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_210),
.B(n_227),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_216),
.CI(n_217),
.CON(n_210),
.SN(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_214),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_245),
.B2(n_246),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_235),
.C(n_246),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_241),
.C(n_244),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_238),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_249),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_268),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_251),
.B(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_261),
.C(n_267),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_252),
.A2(n_253),
.B1(n_261),
.B2(n_295),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_257),
.C(n_259),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_261),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_263),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_281),
.B(n_285),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_264),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_264),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_265),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_288),
.B2(n_289),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_279),
.B2(n_280),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_280),
.C(n_289),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_276),
.B(n_278),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_276),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_278),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_278),
.A2(n_304),
.B1(n_313),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_287),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_283),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_297),
.B(n_300),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_315),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_313),
.C(n_314),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_306),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_317),
.C(n_321),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_309),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_334),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_339),
.B(n_342),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);


endmodule