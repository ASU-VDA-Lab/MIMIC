module real_aes_9730_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_13;
wire n_15;
wire n_9;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
NOR2xp33_ASAP7_75t_R g13 ( .A(n_0), .B(n_5), .Y(n_13) );
NOR3xp33_ASAP7_75t_SL g11 ( .A(n_1), .B(n_6), .C(n_12), .Y(n_11) );
NAND2xp33_ASAP7_75t_R g12 ( .A(n_2), .B(n_13), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
NOR4xp25_ASAP7_75t_SL g9 ( .A(n_4), .B(n_10), .C(n_14), .D(n_15), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_9), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
endmodule