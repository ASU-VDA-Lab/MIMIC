module fake_jpeg_30507_n_302 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_302);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_288;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx13_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_65),
.Y(n_83)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_19),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx2_ASAP7_75t_SL g105 ( 
.A(n_66),
.Y(n_105)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_1),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_31),
.B1(n_30),
.B2(n_37),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_37),
.B1(n_26),
.B2(n_41),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_98),
.B1(n_55),
.B2(n_68),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_104),
.B1(n_108),
.B2(n_39),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_39),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_26),
.B1(n_29),
.B2(n_44),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_49),
.A2(n_40),
.B1(n_31),
.B2(n_26),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_44),
.B1(n_29),
.B2(n_40),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_119),
.B1(n_126),
.B2(n_130),
.Y(n_152)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g156 ( 
.A(n_113),
.Y(n_156)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_124),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_71),
.B1(n_33),
.B2(n_34),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_54),
.B1(n_61),
.B2(n_58),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_140),
.B1(n_56),
.B2(n_109),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_127),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_32),
.B1(n_22),
.B2(n_21),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_132),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_32),
.B1(n_46),
.B2(n_22),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_33),
.B1(n_46),
.B2(n_38),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_133),
.B(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_47),
.C(n_50),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_85),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_135),
.Y(n_148)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_137),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_36),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_35),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_35),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_80),
.C(n_96),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_153),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_98),
.B1(n_78),
.B2(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_120),
.B1(n_102),
.B2(n_92),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_132),
.B(n_142),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_158),
.B(n_143),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_140),
.B(n_39),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_169),
.B(n_174),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_140),
.B1(n_97),
.B2(n_91),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_162),
.B1(n_157),
.B2(n_153),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_170),
.B1(n_175),
.B2(n_147),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_171),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_137),
.B(n_136),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_84),
.B1(n_115),
.B2(n_112),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_137),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_106),
.B1(n_124),
.B2(n_127),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_121),
.B1(n_134),
.B2(n_135),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_35),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_153),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_182),
.B1(n_167),
.B2(n_175),
.Y(n_203)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_162),
.A3(n_158),
.B1(n_157),
.B2(n_66),
.C1(n_40),
.C2(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_192),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_191),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_159),
.B(n_150),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_145),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_196),
.C(n_145),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_147),
.B(n_143),
.C(n_159),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_R g194 ( 
.A(n_169),
.B(n_156),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_174),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_163),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_191),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_201),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_205),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_164),
.B1(n_166),
.B2(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_164),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_204),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_203),
.A2(n_182),
.B1(n_187),
.B2(n_189),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_213),
.Y(n_220)
);

OAI21x1_ASAP7_75t_R g208 ( 
.A1(n_192),
.A2(n_156),
.B(n_146),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_184),
.A3(n_193),
.B1(n_183),
.B2(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_150),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_176),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_187),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_146),
.B(n_114),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_196),
.C(n_188),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_227),
.C(n_228),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_225),
.B1(n_123),
.B2(n_102),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_203),
.B1(n_199),
.B2(n_206),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_179),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_207),
.C(n_201),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_128),
.C(n_156),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_198),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_211),
.B1(n_206),
.B2(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_234),
.A2(n_239),
.B1(n_232),
.B2(n_231),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_204),
.B1(n_208),
.B2(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_222),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_239),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_240),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_217),
.B(n_18),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_242),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_227),
.C(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_247),
.C(n_241),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_156),
.C(n_44),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_229),
.B1(n_235),
.B2(n_4),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_113),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_35),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_44),
.B1(n_67),
.B2(n_19),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_256),
.A2(n_27),
.B1(n_3),
.B2(n_5),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_264),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_257),
.C(n_247),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_263),
.C(n_265),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_68),
.C(n_60),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_16),
.C(n_122),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_266),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_16),
.B1(n_3),
.B2(n_5),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_269),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_244),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_249),
.B(n_244),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_8),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_255),
.B(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_2),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_35),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_6),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_7),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_272),
.B(n_277),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_27),
.B1(n_9),
.B2(n_10),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_273),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_272),
.B(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_291),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_282),
.B(n_290),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_8),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_286),
.B(n_9),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_293),
.B(n_13),
.C(n_14),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.C(n_8),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_299),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_13),
.B1(n_15),
.B2(n_35),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_301),
.B(n_13),
.Y(n_302)
);


endmodule