module fake_jpeg_10119_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_40),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_32),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_20),
.B1(n_29),
.B2(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_27),
.B1(n_32),
.B2(n_30),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_71),
.B1(n_27),
.B2(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_70),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_40),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_38),
.C(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_35),
.A2(n_27),
.B1(n_32),
.B2(n_30),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_43),
.B1(n_62),
.B2(n_61),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_78),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_80),
.B1(n_92),
.B2(n_93),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_41),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_87),
.C(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_43),
.B1(n_37),
.B2(n_34),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_45),
.B(n_22),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_101),
.Y(n_135)
);

OR2x4_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_42),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_102),
.B(n_111),
.Y(n_133)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_33),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_91),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_66),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_109),
.C(n_113),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_107),
.Y(n_137)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_120),
.B1(n_95),
.B2(n_26),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_16),
.B(n_17),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_112),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_67),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_116),
.Y(n_148)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_122),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_28),
.B1(n_24),
.B2(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_98),
.B(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_90),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_73),
.B1(n_88),
.B2(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_131),
.B1(n_151),
.B2(n_139),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_80),
.B1(n_79),
.B2(n_56),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_136),
.B1(n_145),
.B2(n_147),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_69),
.B1(n_63),
.B2(n_64),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_139),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_92),
.B1(n_69),
.B2(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_82),
.C(n_81),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_105),
.C(n_100),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_92),
.B1(n_56),
.B2(n_70),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_104),
.Y(n_167)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_104),
.B(n_28),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_98),
.A2(n_82),
.B1(n_81),
.B2(n_83),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_170),
.B1(n_145),
.B2(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_164),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_123),
.B(n_122),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_162),
.B(n_167),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_102),
.B1(n_83),
.B2(n_101),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_165),
.B1(n_177),
.B2(n_178),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_119),
.B(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_127),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_134),
.B1(n_126),
.B2(n_129),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_172),
.C(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_100),
.C(n_109),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_142),
.B(n_137),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_81),
.B1(n_54),
.B2(n_110),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_171),
.A2(n_174),
.B(n_130),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_93),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_115),
.B(n_33),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_83),
.B1(n_97),
.B2(n_107),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_107),
.B1(n_54),
.B2(n_116),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_37),
.B1(n_28),
.B2(n_24),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_131),
.B1(n_137),
.B2(n_147),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_141),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_191),
.C(n_198),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_199),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_150),
.B1(n_132),
.B2(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_195),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_197),
.Y(n_213)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_170),
.B1(n_179),
.B2(n_165),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_149),
.B1(n_138),
.B2(n_130),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_173),
.B1(n_158),
.B2(n_168),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_194),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_202),
.B1(n_176),
.B2(n_175),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_129),
.C(n_135),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_138),
.B1(n_135),
.B2(n_24),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_72),
.B1(n_37),
.B2(n_29),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_174),
.A2(n_29),
.B(n_26),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_72),
.B1(n_94),
.B2(n_26),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_207),
.A2(n_157),
.B1(n_154),
.B2(n_22),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_209),
.A2(n_222),
.B1(n_223),
.B2(n_229),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_172),
.C(n_163),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_214),
.C(n_224),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_163),
.C(n_164),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_182),
.B(n_167),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_230),
.B1(n_203),
.B2(n_207),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_169),
.C(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_19),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_206),
.A2(n_94),
.B1(n_19),
.B2(n_17),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_196),
.B1(n_202),
.B2(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_16),
.B1(n_15),
.B2(n_21),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_15),
.C(n_1),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_186),
.B1(n_194),
.B2(n_188),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_243),
.B1(n_230),
.B2(n_228),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_189),
.B1(n_184),
.B2(n_183),
.Y(n_236)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_237),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_182),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_185),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_183),
.B1(n_195),
.B2(n_187),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_224),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_249),
.C(n_213),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_203),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_0),
.B(n_1),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_252),
.B(n_2),
.Y(n_270)
);

AOI321xp33_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_233),
.A3(n_218),
.B1(n_208),
.B2(n_231),
.C(n_220),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_252)
);

NAND2x1p5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_21),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_229),
.B(n_208),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_215),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_221),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_0),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_266),
.Y(n_289)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_223),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_262),
.C(n_265),
.Y(n_283)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_269),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_33),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_33),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_65),
.C(n_58),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_271),
.C(n_4),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_244),
.C(n_238),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_2),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_273),
.A2(n_243),
.B1(n_235),
.B2(n_234),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_275),
.A2(n_281),
.B(n_7),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_268),
.B(n_258),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_248),
.B1(n_237),
.B2(n_253),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_251),
.B1(n_246),
.B2(n_241),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_284),
.B1(n_7),
.B2(n_8),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_250),
.B1(n_245),
.B2(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_288),
.Y(n_291)
);

NOR4xp25_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_7),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_4),
.C(n_6),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_7),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_263),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_295),
.Y(n_305)
);

HAxp5_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_283),
.CON(n_304),
.SN(n_304)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_300),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_265),
.B(n_8),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_290),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_276),
.B(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_282),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_8),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_9),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_304),
.A2(n_310),
.B1(n_294),
.B2(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_278),
.B1(n_280),
.B2(n_277),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_288),
.Y(n_312)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_303),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_315),
.A2(n_320),
.B(n_9),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_300),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_321),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_305),
.A2(n_13),
.B(n_10),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_311),
.B(n_307),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_315),
.B(n_316),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_326),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_319),
.A2(n_10),
.B(n_11),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_323),
.B(n_318),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_328),
.B(n_325),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_11),
.B(n_12),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_12),
.B1(n_13),
.B2(n_211),
.Y(n_332)
);


endmodule