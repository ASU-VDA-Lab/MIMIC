module fake_jpeg_27866_n_382 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_38),
.Y(n_100)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_49),
.B(n_31),
.Y(n_98)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_61),
.Y(n_69)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_28),
.A2(n_12),
.B(n_11),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_26),
.B(n_29),
.C(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_26),
.B(n_29),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_30),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_70),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_17),
.B1(n_27),
.B2(n_21),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_66),
.A2(n_34),
.B1(n_25),
.B2(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_27),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_91),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_17),
.B1(n_29),
.B2(n_31),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_84),
.B1(n_61),
.B2(n_51),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_81),
.B(n_82),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_33),
.C(n_30),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_33),
.C(n_38),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_19),
.B1(n_31),
.B2(n_23),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_1),
.Y(n_133)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_22),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_19),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_50),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_105),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_59),
.B1(n_55),
.B2(n_50),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_110),
.B1(n_113),
.B2(n_139),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_60),
.B1(n_55),
.B2(n_40),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_120),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_60),
.B1(n_46),
.B2(n_45),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_123),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_121),
.B1(n_124),
.B2(n_90),
.Y(n_166)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_97),
.Y(n_162)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_18),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_138),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_13),
.B1(n_10),
.B2(n_34),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_63),
.A2(n_10),
.B1(n_34),
.B2(n_33),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_64),
.B(n_34),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_128),
.Y(n_161)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_130),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_74),
.B(n_43),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_133),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_135),
.Y(n_142)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_97),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_65),
.B(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_25),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_71),
.A2(n_34),
.B1(n_25),
.B2(n_4),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_87),
.B(n_77),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_158),
.B(n_118),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_90),
.B1(n_67),
.B2(n_63),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_151),
.A2(n_168),
.B1(n_174),
.B2(n_93),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_67),
.B1(n_85),
.B2(n_94),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_104),
.B1(n_128),
.B2(n_132),
.Y(n_187)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_87),
.B(n_77),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_113),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_109),
.A2(n_72),
.B1(n_94),
.B2(n_85),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_169),
.B1(n_175),
.B2(n_104),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_72),
.B1(n_95),
.B2(n_75),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_120),
.A2(n_75),
.B1(n_25),
.B2(n_73),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx5_ASAP7_75t_SL g171 ( 
.A(n_122),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_116),
.B1(n_122),
.B2(n_102),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_2),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_172),
.B(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_110),
.A2(n_73),
.B1(n_93),
.B2(n_5),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_105),
.A2(n_93),
.B1(n_3),
.B2(n_5),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_182),
.B(n_211),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_179),
.A2(n_208),
.B1(n_210),
.B2(n_153),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_129),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_196),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_112),
.B1(n_103),
.B2(n_127),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_111),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_185),
.Y(n_216)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_198),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_103),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_205),
.B1(n_146),
.B2(n_157),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_188),
.A2(n_212),
.B1(n_164),
.B2(n_153),
.Y(n_247)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_191),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_133),
.B1(n_127),
.B2(n_128),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_202),
.B1(n_207),
.B2(n_156),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_133),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_199),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_137),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_203),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_141),
.B(n_119),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_135),
.B1(n_126),
.B2(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_213),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_148),
.A2(n_93),
.B1(n_3),
.B2(n_6),
.Y(n_207)
);

INVx5_ASAP7_75t_SL g209 ( 
.A(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_157),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_147),
.A2(n_145),
.B1(n_151),
.B2(n_174),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_169),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_150),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_9),
.C(n_3),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_215),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_156),
.B(n_158),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_217),
.A2(n_227),
.B(n_232),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_172),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_222),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_228),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_156),
.B(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_147),
.B1(n_168),
.B2(n_161),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_238),
.B1(n_247),
.B2(n_190),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_205),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_241),
.B1(n_244),
.B2(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_180),
.B(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_235),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_166),
.B(n_141),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_237),
.B(n_213),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_178),
.B(n_181),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_179),
.A2(n_164),
.B1(n_175),
.B2(n_157),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_192),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_200),
.B1(n_193),
.B2(n_177),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_198),
.C(n_197),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_252),
.C(n_265),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_177),
.B1(n_208),
.B2(n_179),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_253),
.B1(n_221),
.B2(n_235),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_196),
.C(n_211),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_190),
.B1(n_204),
.B2(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_264),
.B1(n_266),
.B2(n_268),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_256),
.A2(n_245),
.B(n_225),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_261),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_191),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_189),
.B1(n_159),
.B2(n_8),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_218),
.C(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_189),
.B1(n_159),
.B2(n_8),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_224),
.A2(n_228),
.B1(n_214),
.B2(n_248),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_159),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_230),
.C(n_216),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_222),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_231),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_216),
.B(n_2),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_277),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_9),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_278),
.A2(n_285),
.B(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_223),
.Y(n_287)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_263),
.A2(n_231),
.B(n_240),
.Y(n_288)
);

NAND2x1_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_271),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_273),
.B(n_271),
.Y(n_304)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_241),
.B1(n_219),
.B2(n_239),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_296),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_243),
.B(n_230),
.C(n_244),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_291),
.A2(n_7),
.B1(n_289),
.B2(n_290),
.Y(n_320)
);

BUFx4f_ASAP7_75t_SL g293 ( 
.A(n_254),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_293),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_269),
.Y(n_303)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_262),
.A2(n_250),
.B(n_258),
.C(n_261),
.D(n_265),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_252),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_237),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_300),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_262),
.A2(n_220),
.B(n_246),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_264),
.B1(n_267),
.B2(n_253),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_307),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_304),
.Y(n_336)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_268),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_309),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_283),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_277),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_278),
.B(n_291),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_275),
.B1(n_246),
.B2(n_226),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_246),
.B1(n_226),
.B2(n_9),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_319),
.B1(n_292),
.B2(n_279),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_321),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_299),
.B(n_288),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_326),
.A2(n_332),
.B(n_337),
.Y(n_350)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_281),
.C(n_294),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_303),
.C(n_339),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_280),
.B1(n_291),
.B2(n_295),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_335),
.A2(n_312),
.B1(n_319),
.B2(n_311),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_291),
.B(n_280),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_317),
.B(n_313),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_342),
.C(n_344),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_341),
.A2(n_338),
.B1(n_324),
.B2(n_332),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_307),
.C(n_308),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_322),
.C(n_306),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_310),
.C(n_321),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_346),
.B(n_335),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_304),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_326),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_333),
.Y(n_348)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_324),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_351),
.Y(n_360)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_327),
.B(n_343),
.C(n_350),
.Y(n_354)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_346),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_356),
.A2(n_361),
.B(n_336),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_358),
.A2(n_341),
.B(n_328),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_329),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_362),
.Y(n_369)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_367),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_353),
.B(n_344),
.Y(n_365)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_325),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_370),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_SL g370 ( 
.A(n_357),
.B(n_342),
.Y(n_370)
);

A2O1A1Ixp33_ASAP7_75t_SL g375 ( 
.A1(n_366),
.A2(n_356),
.B(n_354),
.C(n_361),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_375),
.A2(n_355),
.B(n_347),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_373),
.A2(n_369),
.B1(n_368),
.B2(n_357),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_377),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_293),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_378),
.Y(n_380)
);

OAI321xp33_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_371),
.A3(n_374),
.B1(n_340),
.B2(n_312),
.C(n_302),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_302),
.Y(n_382)
);


endmodule