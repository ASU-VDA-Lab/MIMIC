module real_jpeg_30502_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_1),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_1),
.B(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_12),
.B1(n_44),
.B2(n_47),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_2),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_3),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g196 ( 
.A(n_3),
.B(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_6),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_6),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_8),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_8),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_8),
.B(n_47),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_89),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_8),
.B(n_117),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_8),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_8),
.B(n_296),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_8),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

NAND2x1_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_10),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_10),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_10),
.B(n_25),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_10),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

NAND2x1_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_12),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_12),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_12),
.B(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_12),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_12),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_12),
.B(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_13),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_14),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_R g211 ( 
.A(n_14),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_14),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_15),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_15),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_15),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_15),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_15),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_15),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_15),
.B(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_222),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_219),
.Y(n_17)
);

HB1xp67_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_176),
.Y(n_19)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_20),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.C(n_144),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_21),
.B(n_398),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_62),
.B(n_100),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_23),
.B(n_40),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_23),
.B(n_41),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_23)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_27),
.Y(n_267)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_27),
.Y(n_316)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_31),
.B(n_36),
.C(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_36),
.B(n_192),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_36),
.A2(n_37),
.B1(n_192),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_38),
.Y(n_367)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_50),
.B2(n_61),
.Y(n_41)
);

OA21x2_ASAP7_75t_SL g232 ( 
.A1(n_42),
.A2(n_233),
.B(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_43),
.B(n_160),
.C(n_161),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_51),
.Y(n_161)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_56),
.Y(n_352)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_57),
.Y(n_160)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_60),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_62),
.B(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_79),
.C(n_93),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_64),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_66),
.B(n_74),
.C(n_75),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_70),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_72),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_78),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_79),
.B(n_93),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.C(n_88),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_80),
.A2(n_88),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_80),
.Y(n_260)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_83),
.Y(n_299)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_83),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_84),
.B(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_86),
.Y(n_354)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_88),
.Y(n_259)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_92),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_94),
.B(n_98),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_97),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_97),
.B(n_376),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_97),
.B(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_98),
.B(n_107),
.C(n_109),
.Y(n_208)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_99),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_102),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_104),
.B(n_142),
.C(n_143),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_107),
.B(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_107),
.B(n_291),
.Y(n_328)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_108),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_109),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_128),
.B1(n_142),
.B2(n_143),
.Y(n_112)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_124),
.C(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_121),
.Y(n_382)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_128),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.C(n_138),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_131),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_134),
.B1(n_138),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_137),
.Y(n_198)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_145),
.B(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_162),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_158),
.B2(n_159),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_153),
.C(n_157),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_154),
.Y(n_270)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_163),
.B(n_167),
.Y(n_405)
);

XOR2x2_ASAP7_75t_L g404 ( 
.A(n_166),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_173),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_168),
.A2(n_169),
.B1(n_185),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_169),
.Y(n_185)
);

OR2x2_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_202),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_192),
.Y(n_302)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_193),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_218),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_395),
.B(n_412),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_303),
.B(n_394),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_280),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_226),
.B(n_280),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_255),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_227),
.B(n_256),
.C(n_278),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_241),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_229),
.B(n_232),
.C(n_241),
.Y(n_403)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_249),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_242),
.A2(n_243),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_245),
.B1(n_249),
.B2(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_247),
.B(n_310),
.Y(n_374)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_278),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_276),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_276),
.B1(n_277),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_268),
.C(n_271),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_262),
.A2(n_263),
.B1(n_271),
.B2(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_268),
.B(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.C(n_288),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_282),
.B(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_285),
.B(n_288),
.Y(n_392)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_295),
.C(n_300),
.Y(n_288)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_293),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_295),
.A2(n_300),
.B1(n_301),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_388),
.B(n_393),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_343),
.B(n_387),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_329),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_306),
.B(n_329),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_320),
.C(n_328),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_307),
.B(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_317),
.C(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_320),
.A2(n_321),
.B1(n_328),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_322),
.A2(n_325),
.B1(n_326),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_337),
.B1(n_341),
.B2(n_342),
.Y(n_329)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_342),
.C(n_390),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_337),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_358),
.B(n_386),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_355),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_355),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.C(n_353),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_347),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_349),
.B(n_353),
.Y(n_362)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_372),
.B(n_385),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_363),
.Y(n_385)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_364),
.A2(n_365),
.B1(n_368),
.B2(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_379),
.B(n_384),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_383),
.Y(n_384)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_391),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_406),
.Y(n_395)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_400),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.C(n_404),
.Y(n_400)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_401),
.Y(n_411)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_403),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_408),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B(n_416),
.Y(n_413)
);


endmodule