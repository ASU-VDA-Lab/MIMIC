module fake_jpeg_25171_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_7),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_19),
.Y(n_28)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_40),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_25),
.B(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_14),
.Y(n_40)
);

OR2x4_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_24),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_43),
.B(n_30),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_14),
.B1(n_18),
.B2(n_15),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_27),
.B(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_13),
.B1(n_17),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_29),
.B1(n_35),
.B2(n_22),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_27),
.C(n_23),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_30),
.C(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_63),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_56),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_47),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_0),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_22),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_48),
.C(n_46),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_46),
.B(n_35),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_1),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_71),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_70),
.C(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_61),
.B(n_52),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_13),
.B(n_3),
.C(n_4),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_2),
.B(n_3),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_53),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_80),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_79),
.B(n_81),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_56),
.C(n_52),
.Y(n_79)
);

AO221x1_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_49),
.B1(n_51),
.B2(n_60),
.C(n_6),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_82),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_51),
.B(n_10),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_67),
.B1(n_72),
.B2(n_70),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_68),
.B1(n_84),
.B2(n_73),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_88),
.A2(n_77),
.B(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_93),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_73),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_85),
.C(n_87),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_99),
.C(n_5),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_85),
.A3(n_90),
.B1(n_10),
.B2(n_66),
.C1(n_13),
.C2(n_5),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_90),
.Y(n_101)
);

OAI21x1_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_95),
.B(n_92),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_2),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_6),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_105),
.Y(n_107)
);


endmodule