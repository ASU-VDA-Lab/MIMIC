module fake_jpeg_3454_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_46),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_40),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_53),
.B1(n_51),
.B2(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_72),
.B1(n_50),
.B2(n_55),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_54),
.B1(n_43),
.B2(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_45),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_44),
.B(n_48),
.C(n_40),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_79),
.B(n_89),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_0),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_107),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_43),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_52),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_44),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_9),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_42),
.Y(n_97)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_42),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_54),
.B1(n_52),
.B2(n_47),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_109),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_70),
.A3(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_111),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_70),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_0),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_5),
.B(n_6),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_126),
.B(n_11),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_122),
.B(n_123),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_120)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_121),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_25),
.B1(n_38),
.B2(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_11),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_21),
.B1(n_35),
.B2(n_34),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_114),
.C(n_108),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_134),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_17),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_118),
.B1(n_125),
.B2(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_143),
.B1(n_129),
.B2(n_130),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_110),
.B(n_109),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_128),
.B(n_132),
.C(n_127),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_147),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_144),
.C(n_134),
.Y(n_149)
);

AOI31xp33_ASAP7_75t_L g151 ( 
.A1(n_149),
.A2(n_138),
.A3(n_139),
.B(n_148),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_145),
.B1(n_139),
.B2(n_150),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_133),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_12),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_22),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_27),
.B(n_28),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_29),
.Y(n_157)
);


endmodule