module real_jpeg_26716_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_322, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_322;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx11_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_0),
.B(n_198),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_3),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_44),
.B1(n_46),
.B2(n_110),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_3),
.A2(n_22),
.B1(n_26),
.B2(n_110),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_110),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_59),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_5),
.A2(n_22),
.B1(n_26),
.B2(n_59),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_5),
.A2(n_44),
.B1(n_46),
.B2(n_59),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_6),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_6),
.A2(n_34),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_57),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_75),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_34),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_22),
.B(n_40),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_25),
.B(n_28),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_38),
.Y(n_192)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_10),
.A2(n_44),
.B1(n_46),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_10),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_53),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_22),
.B1(n_26),
.B2(n_53),
.Y(n_104)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_85),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_83),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_77),
.Y(n_14)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_68),
.C(n_70),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_16),
.A2(n_17),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.C(n_54),
.Y(n_17)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_18),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_18),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_18),
.A2(n_112),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_18),
.B(n_35),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_31),
.B(n_32),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_19),
.A2(n_103),
.B(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_20),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_20),
.B(n_104),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_20),
.B(n_168),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_22),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_22),
.A2(n_24),
.B(n_34),
.C(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_27),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_27),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_27),
.B(n_33),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_30),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_31),
.B(n_34),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_31),
.A2(n_169),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_34),
.A2(n_39),
.B(n_44),
.C(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_34),
.B(n_98),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_47),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_36),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_42),
.B(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_37),
.A2(n_48),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_39),
.B(n_44),
.C(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_38),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_38),
.B(n_52),
.Y(n_145)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_43),
.B(n_49),
.Y(n_164)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_44),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_46),
.B(n_62),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_116),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_49),
.A2(n_261),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_54),
.A2(n_55),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_63),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_60),
.B(n_61),
.C(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_61),
.Y(n_67)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_60),
.A2(n_66),
.B(n_81),
.Y(n_285)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_64),
.B(n_108),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_66),
.B(n_81),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_68),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_68),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_68),
.A2(n_70),
.B1(n_245),
.B2(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_70),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_71),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_74),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_79),
.B(n_121),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_313),
.B(n_319),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_289),
.A3(n_308),
.B1(n_311),
.B2(n_312),
.C(n_322),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_269),
.B(n_288),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_249),
.B(n_268),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_151),
.B(n_231),
.C(n_248),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_137),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_91),
.B(n_137),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_117),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_106),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_93),
.B(n_106),
.C(n_117),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_94),
.B(n_102),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_99),
.B(n_100),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_95),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_96),
.A2(n_97),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_96),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_101),
.Y(n_100)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_97),
.B(n_150),
.Y(n_196)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_100),
.B(n_197),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_103),
.B(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_105),
.B(n_167),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.C(n_113),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_111),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_112),
.B(n_293),
.C(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_119),
.B(n_124),
.C(n_127),
.Y(n_246)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_134),
.B(n_196),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_135),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_138),
.A2(n_139),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_148),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_145),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_203),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_230),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_223),
.B(n_229),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_181),
.B(n_222),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_170),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_155),
.B(n_170),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.C(n_165),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_156),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_160),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_159),
.A2(n_160),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_159),
.B(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_159),
.A2(n_160),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_160),
.A2(n_280),
.B(n_285),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_164),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_169),
.B(n_178),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_177),
.C(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_217),
.B(n_221),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_199),
.B(n_216),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_184),
.B(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_187),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B(n_215),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_201),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_210),
.B(n_214),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_208),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_246),
.B2(n_247),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_240),
.C(n_247),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_238),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_251),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_267),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_263),
.B2(n_264),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_264),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_257),
.C(n_260),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_271),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_286),
.B2(n_287),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_279),
.C(n_287),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_277),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_291),
.C(n_300),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_278),
.B(n_291),
.CI(n_300),
.CON(n_310),
.SN(n_310)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_301),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_301),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_293),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_303),
.C(n_307),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_310),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);


endmodule