module fake_jpeg_410_n_219 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_219);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_38),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_52),
.Y(n_67)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_29),
.B1(n_14),
.B2(n_31),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_78),
.B1(n_95),
.B2(n_16),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_77),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_21),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_36),
.A2(n_14),
.B1(n_29),
.B2(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_89),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g109 ( 
.A(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_40),
.A2(n_25),
.B1(n_17),
.B2(n_23),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_85),
.B1(n_90),
.B2(n_6),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_25),
.B1(n_28),
.B2(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_34),
.B(n_20),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_20),
.B1(n_31),
.B2(n_18),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_53),
.B1(n_16),
.B2(n_7),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_5),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_5),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_16),
.B1(n_7),
.B2(n_9),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_112),
.B1(n_119),
.B2(n_123),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_63),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_121),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_110),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_112)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_12),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_122),
.Y(n_137)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_68),
.B1(n_88),
.B2(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_63),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_98),
.B1(n_71),
.B2(n_91),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_74),
.C(n_94),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_145),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_138),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_78),
.B(n_95),
.C(n_66),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_98),
.B1(n_71),
.B2(n_91),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_144),
.B1(n_113),
.B2(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_65),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_146),
.Y(n_157)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_143),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_72),
.B1(n_65),
.B2(n_82),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_82),
.C(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_103),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_120),
.B1(n_117),
.B2(n_76),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_161),
.B1(n_162),
.B2(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_76),
.B1(n_111),
.B2(n_113),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_166),
.C(n_154),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_124),
.C(n_129),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_132),
.B(n_136),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g182 ( 
.A1(n_167),
.A2(n_174),
.B(n_148),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_136),
.B(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_153),
.B(n_149),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_142),
.B(n_138),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_126),
.B1(n_133),
.B2(n_150),
.Y(n_180)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_159),
.B1(n_162),
.B2(n_126),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_180),
.B1(n_185),
.B2(n_188),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_168),
.B(n_170),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_129),
.C(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_130),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_148),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_181),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_165),
.C(n_164),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.C(n_135),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_175),
.C(n_176),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_182),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_201),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_202),
.B(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_178),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_181),
.B1(n_176),
.B2(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_161),
.B1(n_173),
.B2(n_156),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_155),
.Y(n_203)
);

AOI31xp67_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_196),
.A3(n_195),
.B(n_193),
.Y(n_206)
);

AOI31xp67_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_130),
.A3(n_109),
.B(n_113),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_203),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_207),
.A2(n_197),
.B1(n_155),
.B2(n_111),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_208),
.C(n_143),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_99),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_214),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_217),
.Y(n_219)
);


endmodule