module fake_jpeg_1406_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_36),
.B1(n_29),
.B2(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_35),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_45),
.B1(n_32),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_58),
.B1(n_38),
.B2(n_3),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_52),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_54),
.B1(n_50),
.B2(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_1),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_2),
.B(n_4),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_9),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_2),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_5),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_84),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_83),
.B1(n_69),
.B2(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_6),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_83)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_88),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_72),
.B1(n_15),
.B2(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_93),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_13),
.B1(n_20),
.B2(n_21),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_99)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_95),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_81),
.C(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_100),
.B(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_92),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_87),
.C(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_91),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_98),
.C(n_88),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_109),
.Y(n_110)
);


endmodule