module fake_jpeg_15193_n_352 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_352);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2x1_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_29),
.B1(n_31),
.B2(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_45),
.Y(n_72)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_37),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_40),
.B1(n_25),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_40),
.B1(n_53),
.B2(n_36),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_37),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_36),
.B(n_26),
.C(n_38),
.Y(n_118)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_87),
.Y(n_108)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_40),
.B1(n_20),
.B2(n_26),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_118),
.B(n_38),
.Y(n_120)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_119),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_101),
.B1(n_107),
.B2(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_19),
.A3(n_27),
.B1(n_22),
.B2(n_34),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_117),
.B(n_38),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_61),
.Y(n_122)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_62),
.A2(n_60),
.B1(n_84),
.B2(n_79),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_113),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_29),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_54),
.B1(n_47),
.B2(n_52),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_46),
.B1(n_52),
.B2(n_50),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_76),
.A2(n_26),
.B1(n_36),
.B2(n_34),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_86),
.B(n_112),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_69),
.C(n_85),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_113),
.B(n_77),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_110),
.C(n_58),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_131),
.Y(n_161)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_69),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_134),
.C(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_27),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_101),
.B1(n_119),
.B2(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_140),
.B1(n_148),
.B2(n_19),
.Y(n_168)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_72),
.B1(n_78),
.B2(n_81),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_105),
.C(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_66),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_63),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_112),
.A3(n_117),
.B1(n_45),
.B2(n_44),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_27),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_108),
.Y(n_150)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_141),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_88),
.B1(n_78),
.B2(n_81),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_156),
.B1(n_164),
.B2(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_117),
.B1(n_97),
.B2(n_106),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_158),
.B(n_166),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_61),
.B1(n_109),
.B2(n_98),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_124),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_58),
.B1(n_96),
.B2(n_46),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_0),
.B(n_1),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_45),
.B1(n_50),
.B2(n_47),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_125),
.B1(n_120),
.B2(n_127),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_39),
.B(n_28),
.C(n_32),
.D(n_37),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_147),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_121),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_184),
.C(n_186),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_183),
.B1(n_190),
.B2(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_160),
.B(n_123),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_187),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_142),
.C(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_132),
.C(n_122),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_128),
.B(n_146),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_155),
.B(n_164),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_193),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_138),
.B1(n_150),
.B2(n_98),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_139),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_192),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_126),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_134),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_145),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_133),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_145),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_202),
.B1(n_179),
.B2(n_175),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_159),
.B1(n_156),
.B2(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_206),
.B1(n_217),
.B2(n_149),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_166),
.B1(n_138),
.B2(n_170),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_165),
.B1(n_152),
.B2(n_149),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_56),
.B1(n_19),
.B2(n_23),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_165),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_208),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_172),
.B1(n_150),
.B2(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_39),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_219),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_108),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_176),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_191),
.B1(n_185),
.B2(n_187),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_143),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_133),
.Y(n_216)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_189),
.B1(n_177),
.B2(n_175),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_108),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_212),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_240),
.B1(n_245),
.B2(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_232),
.C(n_241),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_59),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_203),
.B1(n_211),
.B2(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_143),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_236),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_39),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_239),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_136),
.B1(n_23),
.B2(n_56),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_59),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_196),
.B(n_215),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_246),
.A2(n_261),
.B(n_24),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_227),
.A2(n_217),
.B1(n_201),
.B2(n_210),
.Y(n_255)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_260),
.B1(n_263),
.B2(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_205),
.C(n_208),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.C(n_265),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_205),
.C(n_219),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_213),
.B1(n_200),
.B2(n_2),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_241),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_200),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_56),
.C(n_37),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_228),
.B1(n_237),
.B2(n_230),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_269),
.B(n_270),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_226),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_261),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_278),
.C(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_275),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_240),
.CI(n_231),
.CON(n_275),
.SN(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_233),
.C(n_28),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_282),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_24),
.C(n_35),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_262),
.B1(n_263),
.B2(n_251),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_11),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_284),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_24),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_265),
.C(n_246),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_35),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_293),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_251),
.C(n_254),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_272),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_257),
.C(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_298),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_248),
.C(n_253),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_10),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_302),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_10),
.B1(n_18),
.B2(n_4),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_9),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_275),
.B(n_9),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_305),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_277),
.B1(n_283),
.B2(n_284),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_277),
.B(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_285),
.B(n_281),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_307),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_280),
.B(n_12),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_14),
.B(n_17),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_311),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_35),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_35),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_290),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_12),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_315),
.C(n_296),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_321),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_293),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_322),
.A2(n_323),
.B(n_326),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_316),
.B(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_324),
.B(n_325),
.Y(n_333)
);

OA21x2_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_287),
.B(n_294),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_287),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_328),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_305),
.A2(n_304),
.B1(n_12),
.B2(n_4),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_1),
.C(n_3),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_5),
.B(n_6),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_337),
.B(n_323),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_5),
.Y(n_332)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_332),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_6),
.Y(n_335)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_335),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_8),
.B(n_15),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_17),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_338),
.A2(n_329),
.B(n_15),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_333),
.A2(n_321),
.B(n_14),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_340),
.A2(n_331),
.B(n_334),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_343),
.A2(n_337),
.B(n_330),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_345),
.Y(n_348)
);

HB1xp67_ASAP7_75t_SL g347 ( 
.A(n_346),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_348),
.A2(n_342),
.B(n_341),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_347),
.B(n_339),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_16),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_16),
.B(n_342),
.Y(n_352)
);


endmodule