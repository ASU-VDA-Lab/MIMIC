module fake_jpeg_10952_n_196 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_196);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_13),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_9),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_88),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_59),
.B1(n_72),
.B2(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_100),
.B1(n_73),
.B2(n_64),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_83),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_59),
.B1(n_72),
.B2(n_67),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_76),
.B1(n_65),
.B2(n_81),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_68),
.C(n_74),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_79),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_108),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_124),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_111),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_77),
.B(n_61),
.C(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_82),
.B(n_78),
.C(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_118),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_95),
.B1(n_101),
.B2(n_98),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_151)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_21),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_124),
.B1(n_128),
.B2(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_75),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_82),
.B(n_75),
.C(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_4),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_73),
.B1(n_64),
.B2(n_58),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_146),
.B1(n_147),
.B2(n_151),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_22),
.Y(n_168)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_142),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_49),
.B(n_25),
.C(n_28),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_35),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_140),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_10),
.B(n_11),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_154),
.B(n_166),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_11),
.B(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_14),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_161),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_170),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_34),
.C(n_16),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_164),
.C(n_31),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_168),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_47),
.C(n_17),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_14),
.B(n_19),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_146),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_167),
.C(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_178),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_151),
.B1(n_142),
.B2(n_132),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_153),
.B1(n_136),
.B2(n_154),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_165),
.B(n_139),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_171),
.B1(n_179),
.B2(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_185),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_174),
.B(n_167),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_187),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_188),
.C(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_181),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_192),
.A2(n_176),
.B1(n_164),
.B2(n_162),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_177),
.B(n_168),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_45),
.B(n_33),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_32),
.Y(n_196)
);


endmodule