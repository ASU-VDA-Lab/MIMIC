module fake_aes_4421_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x2_ASAP7_75t_L g11 ( .A(n_7), .B(n_6), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
INVx6_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_12), .B(n_13), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_18), .B(n_16), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_11), .B(n_13), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_18), .B1(n_21), .B2(n_14), .Y(n_27) );
AOI211xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_14), .B(n_12), .C(n_3), .Y(n_28) );
XNOR2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_1), .Y(n_29) );
NOR3x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_1), .C(n_2), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_2), .Y(n_31) );
NOR3xp33_ASAP7_75t_L g32 ( .A(n_30), .B(n_3), .C(n_8), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AOI22xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_32), .B1(n_9), .B2(n_10), .Y(n_34) );
endmodule