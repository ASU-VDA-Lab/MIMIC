module fake_jpeg_3430_n_142 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_14),
.B(n_29),
.Y(n_56)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_2),
.B(n_3),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_24),
.B(n_26),
.C(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_37),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_30),
.B(n_24),
.C(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_29),
.B1(n_18),
.B2(n_22),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_34),
.B1(n_41),
.B2(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_27),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_37),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_43),
.B(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_62),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_35),
.B1(n_34),
.B2(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_68),
.B1(n_23),
.B2(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_17),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_43),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_40),
.B(n_36),
.C(n_24),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_75),
.B(n_36),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_89),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_41),
.B1(n_48),
.B2(n_14),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_63),
.B1(n_60),
.B2(n_72),
.Y(n_96)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_23),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_58),
.C(n_70),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_77),
.B(n_81),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_66),
.B(n_75),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_103),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_89),
.B1(n_80),
.B2(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_102),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_64),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_88),
.C(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_78),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_114),
.B(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_93),
.B(n_99),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_103),
.C(n_98),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_115),
.C(n_111),
.Y(n_120)
);

AOI21x1_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_95),
.B(n_94),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_121),
.B1(n_118),
.B2(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_78),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_96),
.B(n_107),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_114),
.B1(n_94),
.B2(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_96),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_2),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_87),
.B(n_74),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_96),
.A3(n_87),
.B1(n_23),
.B2(n_6),
.C1(n_10),
.C2(n_11),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_13),
.B(n_23),
.Y(n_137)
);

OAI31xp33_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_127),
.A3(n_129),
.B(n_125),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_139)
);

AOI21x1_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_133),
.B(n_3),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_3),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_139),
.C(n_4),
.Y(n_142)
);


endmodule