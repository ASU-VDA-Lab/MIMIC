module fake_jpeg_7810_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_19),
.B(n_22),
.C(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_19),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_23),
.B1(n_28),
.B2(n_20),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_45),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_48),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_19),
.B1(n_17),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_58),
.B1(n_68),
.B2(n_39),
.Y(n_90)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_52),
.Y(n_94)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_23),
.Y(n_84)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_17),
.B1(n_28),
.B2(n_31),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_69),
.B1(n_20),
.B2(n_21),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_17),
.B1(n_28),
.B2(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_78),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_40),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_85),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_92),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_91),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_35),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_35),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_38),
.C(n_43),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_63),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_112),
.Y(n_139)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_111),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_43),
.B(n_45),
.C(n_66),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_87),
.B(n_81),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_117),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_39),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_120),
.Y(n_130)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_126),
.B1(n_82),
.B2(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_52),
.B1(n_51),
.B2(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_97),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_64),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_62),
.B1(n_45),
.B2(n_46),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_72),
.A2(n_27),
.B1(n_34),
.B2(n_25),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_53),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_86),
.Y(n_133)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_148),
.B1(n_105),
.B2(n_153),
.Y(n_158)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_84),
.B(n_77),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_143),
.B(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_132),
.B(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_140),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_85),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_73),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_87),
.B(n_81),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_108),
.B(n_111),
.Y(n_161)
);

AO22x1_ASAP7_75t_SL g148 ( 
.A1(n_107),
.A2(n_96),
.B1(n_92),
.B2(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_76),
.B1(n_126),
.B2(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_160),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_159),
.B1(n_166),
.B2(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_109),
.B1(n_98),
.B2(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_162),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_102),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_164),
.C(n_174),
.Y(n_184)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_148),
.B(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_98),
.B1(n_114),
.B2(n_121),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_80),
.B1(n_83),
.B2(n_82),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_21),
.B(n_80),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_175),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_73),
.C(n_53),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_134),
.B(n_130),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_93),
.B1(n_76),
.B2(n_101),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_0),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_1),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_141),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_88),
.C(n_103),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_151),
.C(n_132),
.Y(n_190)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_201),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_183),
.A2(n_200),
.B1(n_99),
.B2(n_27),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_148),
.B1(n_170),
.B2(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_191),
.B1(n_192),
.B2(n_204),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_206),
.C(n_162),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_131),
.B1(n_135),
.B2(n_145),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_131),
.B1(n_145),
.B2(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_198),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_147),
.B(n_155),
.C(n_32),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_205),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_139),
.B1(n_149),
.B2(n_129),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_175),
.C(n_156),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_217),
.C(n_222),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_178),
.B1(n_161),
.B2(n_174),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_216),
.A2(n_225),
.B1(n_231),
.B2(n_202),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_156),
.C(n_157),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_168),
.B1(n_157),
.B2(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_190),
.C(n_204),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_139),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_226),
.C(n_199),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_227),
.B1(n_24),
.B2(n_26),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_189),
.B1(n_195),
.B2(n_182),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_147),
.C(n_144),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_144),
.C(n_33),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_150),
.B1(n_142),
.B2(n_128),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_232),
.B(n_11),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_234),
.B(n_25),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_99),
.B1(n_32),
.B2(n_30),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_205),
.B(n_191),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_256),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_258),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_196),
.C(n_193),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_243),
.C(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_202),
.C(n_33),
.Y(n_243)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_34),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_34),
.C(n_29),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_216),
.B(n_29),
.CI(n_26),
.CON(n_247),
.SN(n_247)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_221),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_34),
.C(n_29),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_249),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_231),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_213),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_1),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_26),
.B1(n_25),
.B2(n_3),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_1),
.C(n_2),
.Y(n_258)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_211),
.A3(n_230),
.B1(n_210),
.B2(n_219),
.C1(n_228),
.C2(n_234),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_263),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_236),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_214),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_269),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_SL g269 ( 
.A1(n_241),
.A2(n_227),
.A3(n_224),
.B1(n_212),
.B2(n_214),
.C1(n_10),
.C2(n_15),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_251),
.B(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_276),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_16),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_257),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_268),
.B(n_262),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_280),
.B(n_291),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_237),
.B(n_238),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_255),
.B1(n_238),
.B2(n_247),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_283),
.B1(n_288),
.B2(n_289),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_247),
.B1(n_254),
.B2(n_248),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_290),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_243),
.C(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_289),
.C(n_274),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_258),
.C(n_253),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_14),
.B(n_13),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_298),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_260),
.B(n_276),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_281),
.B(n_282),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_259),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_273),
.B1(n_272),
.B2(n_13),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_13),
.B1(n_10),
.B2(n_6),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_2),
.C(n_3),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_2),
.C(n_3),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_6),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_4),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_4),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_307),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_287),
.B(n_5),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_309),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_294),
.A2(n_304),
.B(n_303),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_301),
.B1(n_297),
.B2(n_302),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_7),
.B1(n_8),
.B2(n_314),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_6),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_6),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_317),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_7),
.C(n_8),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_321),
.B(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_327),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_310),
.B1(n_7),
.B2(n_8),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_325),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_316),
.B1(n_328),
.B2(n_319),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_7),
.B(n_323),
.C(n_322),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);


endmodule