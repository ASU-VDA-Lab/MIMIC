module fake_jpeg_12093_n_616 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_616);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_616;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx8_ASAP7_75t_SL g50 ( 
.A(n_18),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_62),
.B(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_24),
.B(n_9),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_64),
.B(n_73),
.Y(n_165)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_9),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_33),
.B(n_10),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_18),
.B1(n_8),
.B2(n_12),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_74),
.A2(n_58),
.B1(n_39),
.B2(n_40),
.Y(n_148)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_25),
.B(n_8),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_79),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_30),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_86),
.Y(n_205)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_89),
.B(n_112),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_38),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_93),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_101),
.Y(n_207)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_50),
.Y(n_112)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

BUFx4f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_31),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_122),
.B(n_53),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_43),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_130),
.B(n_144),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_64),
.B(n_43),
.C(n_57),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_57),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_146),
.B(n_13),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_148),
.A2(n_174),
.B1(n_86),
.B2(n_106),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_73),
.A2(n_58),
.B1(n_52),
.B2(n_47),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_154),
.A2(n_157),
.B1(n_163),
.B2(n_175),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_89),
.A2(n_56),
.B1(n_55),
.B2(n_31),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_68),
.B(n_56),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_161),
.B(n_168),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_87),
.A2(n_53),
.B1(n_49),
.B2(n_41),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_55),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_27),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_171),
.B(n_180),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_72),
.A2(n_27),
.B1(n_35),
.B2(n_53),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_85),
.A2(n_35),
.B1(n_39),
.B2(n_52),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_47),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_40),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_184),
.B(n_191),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_63),
.A2(n_32),
.B1(n_28),
.B2(n_44),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_81),
.B1(n_70),
.B2(n_90),
.Y(n_227)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_116),
.A2(n_32),
.B1(n_28),
.B2(n_46),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_46),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_109),
.B(n_53),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_114),
.B(n_53),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_193),
.B(n_202),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_116),
.A2(n_46),
.B1(n_54),
.B2(n_44),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_84),
.B1(n_80),
.B2(n_126),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_127),
.B(n_14),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_209),
.B(n_0),
.Y(n_268)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_139),
.Y(n_211)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_212),
.Y(n_335)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_164),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_214),
.B(n_221),
.Y(n_342)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_215),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_216),
.B(n_230),
.Y(n_284)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_129),
.Y(n_220)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_46),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_152),
.Y(n_224)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_224),
.Y(n_312)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_273),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_235),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_0),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_236),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_136),
.B(n_46),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_231),
.Y(n_316)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_232),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

BUFx8_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_154),
.B(n_0),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_239),
.Y(n_321)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_242),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_243),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_183),
.A2(n_88),
.B1(n_99),
.B2(n_94),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_244),
.A2(n_280),
.B1(n_205),
.B2(n_185),
.Y(n_298)
);

INVx4_ASAP7_75t_SL g245 ( 
.A(n_207),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_245),
.Y(n_317)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_246),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_195),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_248),
.Y(n_340)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_250),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_140),
.A2(n_128),
.B1(n_91),
.B2(n_103),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_251),
.A2(n_254),
.B1(n_259),
.B2(n_264),
.Y(n_289)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_252),
.Y(n_325)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_143),
.A2(n_93),
.B1(n_54),
.B2(n_44),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_146),
.B(n_0),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_262),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_258),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_199),
.A2(n_54),
.B1(n_48),
.B2(n_120),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_188),
.B(n_69),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_261),
.A2(n_278),
.B(n_159),
.Y(n_300)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_179),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_137),
.Y(n_263)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_263),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_181),
.A2(n_48),
.B1(n_12),
.B2(n_18),
.Y(n_264)
);

INVx4_ASAP7_75t_SL g265 ( 
.A(n_147),
.Y(n_265)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_269),
.Y(n_288)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_271),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_163),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_167),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_274),
.B1(n_276),
.B2(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_181),
.A2(n_48),
.B1(n_12),
.B2(n_4),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_275),
.B(n_283),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_142),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_277),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_131),
.A2(n_123),
.B1(n_48),
.B2(n_4),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_132),
.A2(n_7),
.B1(n_16),
.B2(n_4),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_200),
.A2(n_150),
.B1(n_172),
.B2(n_149),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_200),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_281),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_282),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_141),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_298),
.A2(n_240),
.B1(n_243),
.B2(n_248),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_300),
.B(n_6),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_229),
.B(n_156),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_306),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_225),
.B(n_206),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_217),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_271),
.A2(n_169),
.B1(n_153),
.B2(n_189),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_309),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_211),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_310),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_212),
.B(n_182),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_232),
.C(n_281),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_230),
.A2(n_197),
.B1(n_155),
.B2(n_177),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g331 ( 
.A(n_236),
.B(n_147),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_331),
.B(n_231),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_262),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_334),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_256),
.B(n_206),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_235),
.Y(n_347)
);

OAI22x1_ASAP7_75t_SL g341 ( 
.A1(n_261),
.A2(n_147),
.B1(n_197),
.B2(n_150),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_231),
.B1(n_266),
.B2(n_228),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_343),
.B(n_366),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_346),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_349),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_255),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_299),
.B(n_249),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_354),
.Y(n_408)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_218),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_212),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_356),
.B(n_365),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_238),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_362),
.C(n_379),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_292),
.A2(n_198),
.B1(n_138),
.B2(n_278),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_359),
.B1(n_361),
.B2(n_371),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_316),
.A2(n_198),
.B1(n_138),
.B2(n_149),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_335),
.A2(n_172),
.B1(n_178),
.B2(n_160),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_285),
.B(n_221),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_368),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_364),
.A2(n_366),
.B1(n_372),
.B2(n_374),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_263),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_341),
.A2(n_243),
.B1(n_237),
.B2(n_221),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_284),
.A2(n_214),
.B(n_213),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_383),
.B(n_317),
.Y(n_405)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_373),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_335),
.A2(n_160),
.B1(n_178),
.B2(n_205),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_267),
.B1(n_226),
.B2(n_224),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_285),
.A2(n_241),
.B1(n_242),
.B2(n_219),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_315),
.A2(n_260),
.B1(n_258),
.B2(n_269),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_375),
.A2(n_387),
.B1(n_317),
.B2(n_291),
.Y(n_396)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_300),
.A2(n_245),
.B(n_233),
.C(n_265),
.Y(n_377)
);

AO22x1_ASAP7_75t_L g399 ( 
.A1(n_377),
.A2(n_317),
.B1(n_340),
.B2(n_329),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_381),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_276),
.C(n_277),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_288),
.B(n_272),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_234),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_318),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_322),
.A2(n_233),
.B(n_252),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_287),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_384),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_233),
.C(n_215),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_342),
.C(n_336),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_336),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_388),
.A2(n_399),
.B(n_405),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_396),
.A2(n_400),
.B1(n_424),
.B2(n_364),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_397),
.B(n_413),
.C(n_414),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_382),
.A2(n_289),
.B(n_297),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_398),
.A2(n_411),
.B(n_412),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_354),
.A2(n_315),
.B1(n_303),
.B2(n_325),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_402),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_403),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_381),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_418),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_378),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_386),
.A2(n_324),
.B1(n_303),
.B2(n_325),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_311),
.B(n_291),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_377),
.A2(n_311),
.B(n_305),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_357),
.B(n_332),
.C(n_296),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_362),
.B(n_328),
.C(n_321),
.Y(n_414)
);

AO22x2_ASAP7_75t_L g418 ( 
.A1(n_352),
.A2(n_338),
.B1(n_326),
.B2(n_330),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_346),
.A2(n_295),
.B(n_338),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_419),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_422),
.B(n_383),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_347),
.A2(n_327),
.B1(n_294),
.B2(n_293),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_353),
.A2(n_327),
.B1(n_305),
.B2(n_329),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_426),
.A2(n_371),
.B1(n_361),
.B2(n_375),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_427),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_408),
.A2(n_345),
.B1(n_365),
.B2(n_356),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_428),
.A2(n_432),
.B1(n_442),
.B2(n_444),
.Y(n_476)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_394),
.Y(n_429)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_429),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_431),
.B(n_398),
.Y(n_486)
);

OAI22x1_ASAP7_75t_SL g432 ( 
.A1(n_403),
.A2(n_358),
.B1(n_372),
.B2(n_345),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_433),
.A2(n_435),
.B1(n_437),
.B2(n_443),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_394),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_434),
.B(n_445),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_423),
.A2(n_386),
.B1(n_369),
.B2(n_350),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_436),
.B(n_414),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_391),
.A2(n_351),
.B1(n_384),
.B2(n_380),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_439),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_408),
.A2(n_349),
.B1(n_374),
.B2(n_385),
.Y(n_442)
);

OAI22x1_ASAP7_75t_L g443 ( 
.A1(n_403),
.A2(n_386),
.B1(n_387),
.B2(n_290),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_395),
.A2(n_379),
.B1(n_380),
.B2(n_348),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_395),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_362),
.B1(n_348),
.B2(n_363),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_446),
.A2(n_453),
.B1(n_407),
.B2(n_461),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_391),
.A2(n_355),
.B1(n_368),
.B2(n_370),
.Y(n_447)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_420),
.A2(n_376),
.B1(n_373),
.B2(n_290),
.Y(n_448)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_417),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_451),
.Y(n_475)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_401),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_308),
.C(n_313),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_397),
.C(n_424),
.Y(n_482)
);

AOI22x1_ASAP7_75t_L g457 ( 
.A1(n_399),
.A2(n_330),
.B1(n_308),
.B2(n_313),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_457),
.A2(n_411),
.B(n_400),
.Y(n_483)
);

OAI221xp5_ASAP7_75t_SL g458 ( 
.A1(n_416),
.A2(n_344),
.B1(n_339),
.B2(n_312),
.C(n_314),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_458),
.B(n_399),
.Y(n_492)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_460),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_389),
.B(n_312),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_392),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_462),
.B(n_469),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_438),
.Y(n_465)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_465),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_466),
.B(n_485),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_467),
.A2(n_468),
.B1(n_486),
.B2(n_491),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_446),
.A2(n_389),
.B1(n_393),
.B2(n_412),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_406),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_406),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_472),
.B(n_474),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_413),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_460),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_480),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g480 ( 
.A(n_453),
.B(n_415),
.CI(n_419),
.CON(n_480),
.SN(n_480)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_485),
.C(n_487),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_483),
.A2(n_427),
.B1(n_441),
.B2(n_457),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_409),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_442),
.B(n_415),
.C(n_393),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_450),
.A2(n_452),
.B(n_440),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_489),
.B(n_405),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_450),
.A2(n_452),
.B(n_440),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_428),
.B(n_420),
.C(n_421),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_449),
.C(n_434),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_454),
.A2(n_404),
.B1(n_410),
.B2(n_396),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_492),
.A2(n_439),
.B1(n_451),
.B2(n_459),
.Y(n_503)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_479),
.Y(n_493)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_493),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_429),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_495),
.B(n_497),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_454),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_498),
.B(n_499),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_432),
.C(n_443),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_500),
.B(n_501),
.C(n_519),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_457),
.C(n_435),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_475),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_502),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_503),
.B(n_471),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_514),
.Y(n_525)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_475),
.Y(n_505)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_507),
.A2(n_512),
.B1(n_468),
.B2(n_467),
.Y(n_530)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_484),
.Y(n_508)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_508),
.Y(n_535)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_464),
.Y(n_509)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_509),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_427),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_511),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_476),
.A2(n_441),
.B1(n_433),
.B2(n_404),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_470),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_476),
.A2(n_390),
.B1(n_418),
.B2(n_430),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_480),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_463),
.A2(n_426),
.B1(n_430),
.B2(n_425),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_517),
.A2(n_518),
.B1(n_483),
.B2(n_481),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_491),
.A2(n_425),
.B1(n_418),
.B2(n_402),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_314),
.C(n_418),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_524),
.A2(n_528),
.B1(n_533),
.B2(n_507),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_506),
.A2(n_490),
.B1(n_473),
.B2(n_487),
.Y(n_528)
);

CKINVDCx14_ASAP7_75t_R g529 ( 
.A(n_516),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_539),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_530),
.A2(n_536),
.B1(n_517),
.B2(n_479),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_506),
.A2(n_518),
.B1(n_501),
.B2(n_500),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_538),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_494),
.B(n_478),
.Y(n_537)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_537),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_497),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_493),
.B(n_478),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_486),
.C(n_489),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_540),
.B(n_512),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_418),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_541),
.B(n_543),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_519),
.B(n_418),
.Y(n_543)
);

OAI221xp5_ASAP7_75t_L g544 ( 
.A1(n_535),
.A2(n_504),
.B1(n_495),
.B2(n_496),
.C(n_520),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_544),
.A2(n_546),
.B1(n_560),
.B2(n_561),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_547),
.A2(n_528),
.B1(n_531),
.B2(n_543),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_523),
.B(n_510),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_522),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_513),
.C(n_496),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_550),
.B(n_552),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_529),
.A2(n_486),
.B(n_480),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_551),
.A2(n_557),
.B(n_559),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_513),
.C(n_511),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_539),
.C(n_525),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_402),
.C(n_339),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_556),
.C(n_527),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_526),
.B(n_286),
.C(n_3),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_536),
.A2(n_286),
.B(n_7),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_530),
.A2(n_286),
.B(n_13),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_533),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_524),
.A2(n_2),
.B1(n_16),
.B2(n_531),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_523),
.B(n_16),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_562),
.B(n_534),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_570),
.Y(n_584)
);

FAx1_ASAP7_75t_SL g566 ( 
.A(n_551),
.B(n_540),
.CI(n_541),
.CON(n_566),
.SN(n_566)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_568),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_567),
.Y(n_579)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_548),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_572),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_558),
.B(n_526),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_522),
.C(n_525),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_573),
.B(n_575),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_546),
.A2(n_535),
.B1(n_521),
.B2(n_537),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_574),
.A2(n_560),
.B1(n_561),
.B2(n_554),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_548),
.A2(n_521),
.B(n_527),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_576),
.A2(n_578),
.B(n_557),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_542),
.C(n_2),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_577),
.B(n_576),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_555),
.A2(n_542),
.B(n_545),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_580),
.B(n_563),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_565),
.B(n_556),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_582),
.B(n_591),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_563),
.A2(n_547),
.B(n_559),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_585),
.B(n_566),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_586),
.B(n_587),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_572),
.B(n_573),
.C(n_567),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_566),
.A2(n_549),
.B(n_562),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_588),
.A2(n_581),
.B(n_583),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_570),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_578),
.B(n_577),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_587),
.B(n_571),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_595),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_589),
.C(n_579),
.Y(n_595)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_596),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_598),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_580),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_599),
.B(n_600),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_600),
.A2(n_585),
.B(n_579),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_601),
.A2(n_595),
.B(n_564),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_SL g606 ( 
.A(n_593),
.B(n_597),
.C(n_592),
.Y(n_606)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_606),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_605),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_607),
.B(n_608),
.C(n_610),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_575),
.C(n_604),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_609),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_612),
.A2(n_602),
.B(n_606),
.Y(n_613)
);

BUFx24_ASAP7_75t_SL g614 ( 
.A(n_613),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_611),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_615),
.Y(n_616)
);


endmodule