module fake_aes_5867_n_422 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_422);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_422;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_134;
wire n_233;
wire n_82;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_414;
wire n_350;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g59 ( .A(n_12), .Y(n_59) );
INVx1_ASAP7_75t_L g60 ( .A(n_10), .Y(n_60) );
INVx1_ASAP7_75t_L g61 ( .A(n_53), .Y(n_61) );
INVx1_ASAP7_75t_L g62 ( .A(n_26), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_38), .Y(n_63) );
INVx1_ASAP7_75t_L g64 ( .A(n_17), .Y(n_64) );
INVx1_ASAP7_75t_L g65 ( .A(n_55), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_5), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_46), .Y(n_67) );
INVx1_ASAP7_75t_SL g68 ( .A(n_24), .Y(n_68) );
INVxp33_ASAP7_75t_SL g69 ( .A(n_21), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_42), .Y(n_70) );
INVxp67_ASAP7_75t_SL g71 ( .A(n_20), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_9), .Y(n_72) );
CKINVDCx14_ASAP7_75t_R g73 ( .A(n_5), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_18), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_2), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_1), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_41), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_57), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_43), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_12), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_44), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_18), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_36), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_30), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_13), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_33), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_2), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_17), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_51), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_34), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_0), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_0), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_56), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_13), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_90), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_61), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_61), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_73), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_74), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_62), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_64), .B(n_1), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_63), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_63), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_65), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_64), .B(n_3), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_87), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_65), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_87), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_67), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_82), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_109), .B(n_84), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_97), .B(n_95), .Y(n_118) );
CKINVDCx11_ASAP7_75t_R g119 ( .A(n_112), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_97), .B(n_101), .Y(n_120) );
INVx4_ASAP7_75t_L g121 ( .A(n_110), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_110), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_101), .B(n_82), .Y(n_123) );
NOR2xp33_ASAP7_75t_SL g124 ( .A(n_100), .B(n_95), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_107), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_99), .B(n_69), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_110), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_104), .B(n_78), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_96), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
OR2x2_ASAP7_75t_SL g133 ( .A(n_103), .B(n_66), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_104), .A2(n_66), .B1(n_93), .B2(n_72), .Y(n_134) );
INVx4_ASAP7_75t_SL g135 ( .A(n_111), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_111), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_111), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_106), .A2(n_80), .B1(n_60), .B2(n_76), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_120), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_125), .Y(n_141) );
NOR2xp33_ASAP7_75t_R g142 ( .A(n_131), .B(n_106), .Y(n_142) );
NOR3xp33_ASAP7_75t_SL g143 ( .A(n_117), .B(n_103), .C(n_108), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_127), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_123), .B(n_115), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_118), .B(n_115), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_123), .B(n_116), .Y(n_147) );
INVx1_ASAP7_75t_SL g148 ( .A(n_125), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_124), .B(n_108), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_133), .A2(n_116), .B1(n_98), .B2(n_113), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_130), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_139), .B(n_98), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_119), .Y(n_155) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
BUFx8_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_127), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
INVx1_ASAP7_75t_SL g161 ( .A(n_139), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_121), .B(n_114), .Y(n_163) );
NAND2xp33_ASAP7_75t_R g164 ( .A(n_122), .B(n_114), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
AND2x4_ASAP7_75t_SL g166 ( .A(n_127), .B(n_98), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_134), .B(n_102), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_156), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_152), .B(n_102), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_148), .B(n_68), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_152), .B(n_102), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_140), .B(n_105), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_140), .B(n_105), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_146), .A2(n_105), .B1(n_113), .B2(n_75), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_145), .B(n_113), .Y(n_181) );
BUFx12f_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_161), .A2(n_111), .B1(n_72), .B2(n_75), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_145), .B(n_114), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_147), .A2(n_137), .B(n_132), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_145), .B(n_111), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_157), .B(n_94), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_151), .A2(n_91), .B1(n_93), .B2(n_71), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_158), .B(n_91), .Y(n_196) );
CKINVDCx6p67_ASAP7_75t_R g197 ( .A(n_145), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
INVx8_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_171), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_178), .A2(n_153), .B1(n_143), .B2(n_158), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_172), .B(n_167), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_185), .B(n_162), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_185), .A2(n_167), .B1(n_163), .B2(n_149), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_188), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_197), .B(n_163), .Y(n_208) );
AND2x6_ASAP7_75t_L g209 ( .A(n_188), .B(n_164), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_188), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_179), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_197), .A2(n_163), .B1(n_160), .B2(n_157), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_179), .A2(n_85), .B1(n_77), .B2(n_92), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_197), .A2(n_199), .B1(n_172), .B2(n_196), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_171), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_199), .A2(n_59), .B1(n_88), .B2(n_166), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_172), .B(n_114), .Y(n_217) );
AOI221xp5_ASAP7_75t_L g218 ( .A1(n_184), .A2(n_85), .B1(n_92), .B2(n_77), .C(n_83), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_172), .A2(n_79), .B1(n_81), .B2(n_86), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_199), .A2(n_166), .B1(n_89), .B2(n_156), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_199), .A2(n_166), .B1(n_165), .B2(n_132), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_199), .A2(n_165), .B1(n_137), .B2(n_128), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_199), .A2(n_128), .B1(n_129), .B2(n_138), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_172), .B(n_3), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_210), .Y(n_225) );
OAI221xp5_ASAP7_75t_L g226 ( .A1(n_201), .A2(n_194), .B1(n_196), .B2(n_186), .C(n_183), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_206), .A2(n_180), .B1(n_177), .B2(n_196), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_206), .B(n_177), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_201), .A2(n_189), .B(n_190), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_209), .Y(n_230) );
AND2x6_ASAP7_75t_SL g231 ( .A(n_224), .B(n_182), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_211), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_209), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_211), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_213), .A2(n_189), .B(n_190), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g236 ( .A1(n_210), .A2(n_186), .B1(n_193), .B2(n_182), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_200), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_203), .A2(n_184), .B1(n_181), .B2(n_177), .Y(n_238) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_218), .A2(n_180), .B1(n_184), .B2(n_181), .C(n_194), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_203), .A2(n_181), .B1(n_173), .B2(n_193), .Y(n_240) );
AOI21xp33_ASAP7_75t_SL g241 ( .A1(n_207), .A2(n_193), .B(n_191), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_200), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_208), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_202), .B(n_192), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
OAI221xp5_ASAP7_75t_L g246 ( .A1(n_226), .A2(n_214), .B1(n_204), .B2(n_219), .C(n_213), .Y(n_246) );
OAI33xp33_ASAP7_75t_L g247 ( .A1(n_227), .A2(n_219), .A3(n_232), .B1(n_217), .B2(n_244), .B3(n_234), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_228), .B(n_205), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_232), .Y(n_249) );
OAI211xp5_ASAP7_75t_L g250 ( .A1(n_236), .A2(n_212), .B(n_216), .C(n_183), .Y(n_250) );
OR2x6_ASAP7_75t_L g251 ( .A(n_230), .B(n_193), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_242), .Y(n_252) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_229), .A2(n_215), .B(n_205), .Y(n_253) );
OAI211xp5_ASAP7_75t_L g254 ( .A1(n_226), .A2(n_210), .B(n_208), .C(n_220), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_234), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_227), .A2(n_215), .B1(n_221), .B2(n_195), .Y(n_256) );
OAI332xp33_ASAP7_75t_L g257 ( .A1(n_244), .A2(n_192), .A3(n_195), .B1(n_198), .B2(n_182), .B3(n_9), .C1(n_10), .C2(n_11), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_228), .B(n_198), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_234), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_242), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_239), .A2(n_209), .B1(n_187), .B2(n_176), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_237), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
OAI31xp33_ASAP7_75t_SL g265 ( .A1(n_246), .A2(n_243), .A3(n_239), .B(n_229), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_252), .B(n_230), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_252), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_252), .B(n_230), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g269 ( .A1(n_257), .A2(n_238), .B1(n_240), .B2(n_235), .C(n_243), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_245), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_260), .B(n_262), .Y(n_271) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_256), .A2(n_235), .B(n_241), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_249), .Y(n_273) );
NOR3xp33_ASAP7_75t_SL g274 ( .A(n_246), .B(n_231), .C(n_241), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_260), .B(n_233), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_260), .B(n_233), .Y(n_276) );
AOI33xp33_ASAP7_75t_L g277 ( .A1(n_261), .A2(n_128), .A3(n_129), .B1(n_222), .B2(n_8), .B3(n_11), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_262), .Y(n_278) );
OAI31xp33_ASAP7_75t_L g279 ( .A1(n_254), .A2(n_225), .A3(n_231), .B(n_187), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_262), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_253), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_263), .B(n_233), .Y(n_283) );
NAND2xp67_ASAP7_75t_L g284 ( .A(n_258), .B(n_233), .Y(n_284) );
OAI33xp33_ASAP7_75t_L g285 ( .A1(n_256), .A2(n_4), .A3(n_6), .B1(n_7), .B2(n_8), .B3(n_14), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_255), .B(n_225), .Y(n_286) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_250), .A2(n_225), .B(n_175), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_259), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_259), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_263), .B(n_230), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_265), .B(n_264), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_271), .B(n_253), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_271), .B(n_253), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_271), .B(n_253), .Y(n_295) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_270), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_273), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_290), .B(n_264), .Y(n_299) );
OAI33xp33_ASAP7_75t_L g300 ( .A1(n_280), .A2(n_257), .A3(n_6), .B1(n_7), .B2(n_14), .B3(n_15), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_290), .B(n_248), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_280), .B(n_248), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_265), .B(n_258), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_288), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_269), .B(n_254), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_270), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_284), .B(n_4), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_289), .B(n_245), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_267), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
NOR3xp33_ASAP7_75t_L g312 ( .A(n_285), .B(n_250), .C(n_247), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_267), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_267), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_278), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_283), .B(n_291), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_274), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_279), .B(n_175), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_278), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_281), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_284), .B(n_15), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_281), .B(n_251), .Y(n_323) );
NOR3xp33_ASAP7_75t_SL g324 ( .A(n_285), .B(n_16), .C(n_19), .Y(n_324) );
NOR2xp33_ASAP7_75t_R g325 ( .A(n_283), .B(n_209), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_281), .B(n_251), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_319), .A2(n_287), .B(n_279), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_305), .A2(n_251), .B1(n_291), .B2(n_283), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_292), .B(n_272), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_302), .B(n_291), .Y(n_330) );
OA21x2_ASAP7_75t_L g331 ( .A1(n_303), .A2(n_282), .B(n_266), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_300), .A2(n_272), .B1(n_276), .B2(n_275), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_296), .Y(n_333) );
OAI21xp33_ASAP7_75t_SL g334 ( .A1(n_307), .A2(n_277), .B(n_251), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_318), .A2(n_272), .B(n_282), .C(n_251), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_297), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_324), .A2(n_276), .B1(n_275), .B2(n_268), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_322), .A2(n_268), .B(n_266), .C(n_209), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_310), .B(n_209), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_317), .B(n_22), .Y(n_340) );
XNOR2x1_ASAP7_75t_L g341 ( .A(n_317), .B(n_23), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_317), .A2(n_170), .B1(n_223), .B2(n_187), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_313), .Y(n_343) );
OAI211xp5_ASAP7_75t_L g344 ( .A1(n_312), .A2(n_170), .B(n_175), .C(n_129), .Y(n_344) );
OAI322xp33_ASAP7_75t_L g345 ( .A1(n_298), .A2(n_138), .A3(n_136), .B1(n_174), .B2(n_176), .C1(n_170), .C2(n_175), .Y(n_345) );
AND4x1_ASAP7_75t_L g346 ( .A(n_325), .B(n_209), .C(n_27), .D(n_28), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_308), .A2(n_176), .B1(n_174), .B2(n_175), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_311), .B(n_25), .Y(n_348) );
AOI32xp33_ASAP7_75t_L g349 ( .A1(n_306), .A2(n_174), .A3(n_29), .B1(n_31), .B2(n_32), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_304), .Y(n_350) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_306), .B(n_175), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_301), .B(n_138), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_320), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_326), .A2(n_175), .B1(n_136), .B2(n_37), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_301), .A2(n_136), .B1(n_135), .B2(n_144), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_323), .A2(n_135), .B1(n_168), .B2(n_144), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_293), .A2(n_168), .B1(n_144), .B2(n_159), .C(n_169), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_331), .B(n_294), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_333), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_354), .B(n_294), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_358), .B(n_295), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g366 ( .A(n_329), .B(n_309), .C(n_316), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_334), .B(n_315), .Y(n_367) );
AOI22x1_ASAP7_75t_L g368 ( .A1(n_327), .A2(n_326), .B1(n_315), .B2(n_323), .Y(n_368) );
NOR3xp33_ASAP7_75t_SL g369 ( .A(n_338), .B(n_316), .C(n_309), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_336), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_360), .B(n_332), .Y(n_371) );
NOR4xp25_ASAP7_75t_SL g372 ( .A(n_341), .B(n_321), .C(n_39), .D(n_40), .Y(n_372) );
XNOR2xp5_ASAP7_75t_L g373 ( .A(n_346), .B(n_321), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_353), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_335), .B(n_135), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_330), .B(n_35), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_350), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_328), .B(n_45), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_352), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_348), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_339), .B(n_47), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_340), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_347), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_368), .A2(n_351), .B1(n_342), .B2(n_344), .Y(n_385) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_365), .B(n_345), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_363), .B(n_356), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_367), .A2(n_349), .B(n_355), .C(n_356), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_380), .B(n_359), .Y(n_390) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_378), .B(n_357), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_371), .B(n_357), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_367), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_361), .B(n_52), .Y(n_394) );
XNOR2x1_ASAP7_75t_L g395 ( .A(n_362), .B(n_58), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_375), .B(n_135), .C(n_159), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_386), .A2(n_375), .B(n_368), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_390), .B(n_384), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_389), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_389), .Y(n_400) );
NAND3x1_ASAP7_75t_L g401 ( .A(n_391), .B(n_381), .C(n_376), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_395), .A2(n_373), .B(n_366), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_393), .A2(n_383), .B1(n_392), .B2(n_394), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_385), .A2(n_379), .B1(n_373), .B2(n_382), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_385), .B(n_369), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_387), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g407 ( .A1(n_388), .A2(n_382), .B(n_374), .C(n_370), .Y(n_407) );
AOI211xp5_ASAP7_75t_SL g408 ( .A1(n_396), .A2(n_372), .B(n_364), .C(n_377), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_390), .A2(n_367), .B1(n_380), .B2(n_386), .Y(n_409) );
AOI21xp33_ASAP7_75t_SL g410 ( .A1(n_395), .A2(n_389), .B(n_367), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_399), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_404), .A2(n_405), .B1(n_409), .B2(n_407), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_400), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_410), .A2(n_403), .B(n_397), .C(n_402), .Y(n_414) );
INVx4_ASAP7_75t_L g415 ( .A(n_411), .Y(n_415) );
XNOR2xp5_ASAP7_75t_L g416 ( .A(n_412), .B(n_404), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_413), .B(n_406), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_415), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_417), .Y(n_419) );
XOR2xp5_ASAP7_75t_L g420 ( .A(n_418), .B(n_416), .Y(n_420) );
AO221x1_ASAP7_75t_L g421 ( .A1(n_420), .A2(n_419), .B1(n_414), .B2(n_401), .C(n_408), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_421), .A2(n_419), .B(n_398), .Y(n_422) );
endmodule