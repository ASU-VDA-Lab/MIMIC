module fake_netlist_5_1_n_774 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_774);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_774;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_40),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_72),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_129),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_38),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_6),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_21),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_35),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_15),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_105),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_88),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_141),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_49),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_85),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_94),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_15),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_63),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_60),
.B(n_73),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_61),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_50),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_6),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_20),
.B(n_131),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_67),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_136),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_27),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_127),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_99),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_143),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_75),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_65),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_23),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_31),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

OR2x6_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_195),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_0),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_17),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_0),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_18),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_181),
.B(n_1),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_161),
.B(n_2),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_161),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_191),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_162),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_19),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_171),
.B(n_5),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_180),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_173),
.B(n_9),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_213),
.Y(n_264)
);

NOR2x1p5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_163),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_167),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_217),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_218),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_235),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_225),
.A2(n_256),
.B1(n_224),
.B2(n_231),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_233),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_168),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_215),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_224),
.A2(n_185),
.B1(n_202),
.B2(n_204),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_231),
.B(n_205),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_225),
.B(n_169),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_212),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_210),
.C(n_206),
.Y(n_307)
);

AO21x2_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_200),
.B(n_197),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_235),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_227),
.B(n_172),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_175),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_290),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_229),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_297),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_272),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_277),
.B(n_229),
.Y(n_323)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_283),
.B(n_247),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_222),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_309),
.B(n_277),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_298),
.A2(n_227),
.B1(n_229),
.B2(n_252),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_252),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_245),
.C(n_246),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_298),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_223),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_293),
.A2(n_252),
.B(n_241),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_264),
.B(n_223),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_224),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_271),
.A2(n_228),
.B(n_259),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_271),
.B(n_224),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_259),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_259),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_303),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_305),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_226),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_295),
.B(n_226),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_265),
.A2(n_257),
.B1(n_238),
.B2(n_239),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_270),
.B(n_234),
.C(n_236),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_294),
.B(n_250),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_275),
.A2(n_183),
.B1(n_184),
.B2(n_186),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_251),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_276),
.B(n_234),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_281),
.B(n_188),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_306),
.B(n_251),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_300),
.B(n_251),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_286),
.B(n_193),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_300),
.B(n_251),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_311),
.B(n_304),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_311),
.B(n_251),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_268),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_304),
.B(n_254),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_284),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_288),
.B(n_254),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_284),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_254),
.Y(n_372)
);

NOR2x1p5_ASAP7_75t_L g373 ( 
.A(n_266),
.B(n_236),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_310),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_268),
.B(n_194),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_269),
.B(n_254),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_285),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_269),
.B(n_254),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_SL g379 ( 
.A(n_301),
.B(n_241),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g380 ( 
.A(n_285),
.B(n_255),
.C(n_221),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_287),
.B(n_221),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_269),
.B(n_255),
.Y(n_382)
);

NOR3xp33_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_344),
.C(n_329),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_320),
.A2(n_301),
.B(n_292),
.Y(n_384)
);

AOI21x1_ASAP7_75t_L g385 ( 
.A1(n_340),
.A2(n_292),
.B(n_291),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_317),
.B(n_287),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_291),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_331),
.A2(n_267),
.B(n_278),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_255),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g390 ( 
.A1(n_341),
.A2(n_266),
.B(n_267),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_301),
.B(n_269),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_339),
.C(n_353),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_334),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

CKINVDCx10_ASAP7_75t_R g395 ( 
.A(n_322),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_L g396 ( 
.A1(n_323),
.A2(n_278),
.B(n_273),
.C(n_220),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_335),
.A2(n_301),
.B(n_274),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_R g398 ( 
.A(n_324),
.B(n_22),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_338),
.A2(n_301),
.B(n_274),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_353),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_328),
.B(n_255),
.Y(n_402)
);

O2A1O1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_321),
.A2(n_273),
.B(n_220),
.C(n_255),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_358),
.A2(n_220),
.B(n_274),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_316),
.A2(n_274),
.B(n_241),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_326),
.A2(n_241),
.B1(n_11),
.B2(n_12),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_24),
.Y(n_407)
);

BUFx4f_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

O2A1O1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_357),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_327),
.A2(n_89),
.B1(n_158),
.B2(n_157),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_342),
.B(n_25),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_346),
.B(n_10),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_365),
.A2(n_87),
.B(n_156),
.Y(n_413)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_347),
.A2(n_13),
.B(n_14),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_325),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_363),
.B(n_14),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_343),
.A2(n_91),
.B1(n_26),
.B2(n_28),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_L g419 ( 
.A1(n_355),
.A2(n_16),
.B(n_29),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_367),
.A2(n_95),
.B(n_30),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_32),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_373),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_356),
.A2(n_97),
.B1(n_33),
.B2(n_34),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_324),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_375),
.B(n_16),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_354),
.A2(n_36),
.B(n_37),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_377),
.B(n_39),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_345),
.B(n_41),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_369),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_348),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_318),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_345),
.B(n_54),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_319),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_345),
.B(n_55),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_350),
.B(n_56),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_380),
.A2(n_57),
.B(n_59),
.Y(n_439)
);

AOI21xp33_ASAP7_75t_L g440 ( 
.A1(n_374),
.A2(n_62),
.B(n_64),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_380),
.A2(n_66),
.B(n_68),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_349),
.B(n_361),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_359),
.A2(n_69),
.B(n_70),
.Y(n_443)
);

A2O1A1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_370),
.A2(n_74),
.B(n_77),
.C(n_78),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_325),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_364),
.A2(n_79),
.B(n_80),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_345),
.B(n_82),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_345),
.B(n_83),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_368),
.B(n_86),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_372),
.A2(n_93),
.B(n_96),
.Y(n_451)
);

INVx6_ASAP7_75t_SL g452 ( 
.A(n_395),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_393),
.B(n_382),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_392),
.A2(n_378),
.B1(n_362),
.B2(n_101),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_394),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_396),
.A2(n_379),
.B(n_362),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_383),
.B(n_362),
.Y(n_459)
);

AO22x2_ASAP7_75t_L g460 ( 
.A1(n_427),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_412),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_415),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_387),
.A2(n_103),
.B(n_106),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_107),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g466 ( 
.A1(n_385),
.A2(n_108),
.B(n_109),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_389),
.B(n_111),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_425),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_400),
.A2(n_112),
.B(n_113),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_388),
.A2(n_114),
.B(n_115),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_401),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_122),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_384),
.A2(n_125),
.B(n_126),
.Y(n_473)
);

AOI221xp5_ASAP7_75t_L g474 ( 
.A1(n_414),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_137),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_446),
.A2(n_138),
.B(n_139),
.Y(n_476)
);

CKINVDCx9p33_ASAP7_75t_R g477 ( 
.A(n_408),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_410),
.A2(n_140),
.B1(n_142),
.B2(n_144),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_391),
.A2(n_146),
.B(n_149),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_436),
.B(n_152),
.Y(n_480)
);

A2O1A1Ixp33_ASAP7_75t_L g481 ( 
.A1(n_419),
.A2(n_153),
.B(n_155),
.C(n_160),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_430),
.A2(n_435),
.B(n_448),
.Y(n_482)
);

AOI21x1_ASAP7_75t_SL g483 ( 
.A1(n_438),
.A2(n_411),
.B(n_422),
.Y(n_483)
);

AOI21x1_ASAP7_75t_SL g484 ( 
.A1(n_407),
.A2(n_447),
.B(n_437),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_450),
.A2(n_390),
.B(n_397),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_434),
.Y(n_486)
);

AO21x2_ASAP7_75t_L g487 ( 
.A1(n_404),
.A2(n_451),
.B(n_439),
.Y(n_487)
);

BUFx12f_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

AOI211x1_ASAP7_75t_L g489 ( 
.A1(n_416),
.A2(n_441),
.B(n_423),
.C(n_429),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_408),
.B(n_398),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_405),
.A2(n_428),
.B(n_413),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_402),
.B(n_442),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_421),
.A2(n_443),
.B(n_403),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_431),
.A2(n_424),
.B(n_418),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_432),
.B(n_433),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_415),
.A2(n_417),
.B(n_445),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_409),
.A2(n_406),
.B(n_442),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_445),
.Y(n_498)
);

OAI21xp33_ASAP7_75t_L g499 ( 
.A1(n_444),
.A2(n_440),
.B(n_417),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_392),
.B(n_334),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_395),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_393),
.B(n_330),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_387),
.A2(n_338),
.B(n_404),
.Y(n_505)
);

AOI21xp33_ASAP7_75t_L g506 ( 
.A1(n_504),
.A2(n_461),
.B(n_456),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_485),
.B(n_493),
.Y(n_507)
);

AOI21x1_ASAP7_75t_L g508 ( 
.A1(n_467),
.A2(n_505),
.B(n_472),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_484),
.A2(n_483),
.B(n_469),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_482),
.A2(n_466),
.B(n_479),
.Y(n_510)
);

AOI21xp33_ASAP7_75t_L g511 ( 
.A1(n_456),
.A2(n_501),
.B(n_503),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_474),
.A2(n_476),
.B1(n_495),
.B2(n_460),
.Y(n_512)
);

OAI21x1_ASAP7_75t_SL g513 ( 
.A1(n_476),
.A2(n_464),
.B(n_470),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_464),
.B(n_481),
.C(n_497),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_473),
.A2(n_494),
.B(n_457),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_462),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_465),
.B(n_489),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_459),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_468),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_499),
.A2(n_487),
.B(n_463),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_458),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_488),
.Y(n_526)
);

OAI21x1_ASAP7_75t_SL g527 ( 
.A1(n_475),
.A2(n_471),
.B(n_496),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_487),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_463),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_499),
.A2(n_463),
.B(n_480),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_454),
.A2(n_457),
.B(n_478),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_490),
.A2(n_458),
.B1(n_471),
.B2(n_477),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_452),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

CKINVDCx11_ASAP7_75t_R g535 ( 
.A(n_452),
.Y(n_535)
);

NOR2x1_ASAP7_75t_R g536 ( 
.A(n_502),
.B(n_322),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_333),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_468),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_491),
.A2(n_485),
.B(n_493),
.Y(n_539)
);

AOI221xp5_ASAP7_75t_L g540 ( 
.A1(n_461),
.A2(n_332),
.B1(n_394),
.B2(n_414),
.C(n_296),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_456),
.B(n_309),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_491),
.A2(n_485),
.B(n_493),
.Y(n_543)
);

NOR2x1_ASAP7_75t_SL g544 ( 
.A(n_463),
.B(n_458),
.Y(n_544)
);

AO31x2_ASAP7_75t_L g545 ( 
.A1(n_505),
.A2(n_390),
.A3(n_396),
.B(n_481),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_501),
.B(n_333),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_462),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

AND2x4_ASAP7_75t_SL g549 ( 
.A(n_458),
.B(n_503),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_547),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_548),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_514),
.A2(n_517),
.B(n_509),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_523),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_518),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_535),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_525),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_538),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_515),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_519),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_516),
.Y(n_561)
);

INVx8_ASAP7_75t_L g562 ( 
.A(n_537),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_522),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_525),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_517),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_529),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_546),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_522),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_514),
.A2(n_509),
.B(n_507),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_537),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_544),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_506),
.B(n_512),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_535),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_538),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_540),
.B(n_511),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_549),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_545),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_541),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_545),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_524),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

BUFx4f_ASAP7_75t_SL g582 ( 
.A(n_526),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_520),
.B(n_531),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_549),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_539),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_580),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_580),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_579),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_579),
.Y(n_592)
);

AND2x4_ASAP7_75t_SL g593 ( 
.A(n_553),
.B(n_527),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_570),
.B(n_520),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_586),
.B(n_543),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_554),
.B(n_532),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_575),
.A2(n_513),
.B1(n_530),
.B2(n_534),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_539),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_557),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_567),
.B(n_536),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_553),
.B(n_543),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_510),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_568),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_550),
.B(n_510),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_553),
.B(n_556),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_563),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_568),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_561),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_577),
.Y(n_611)
);

NOR2x1p5_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_508),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_562),
.B(n_533),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_560),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_584),
.B(n_533),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_562),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_572),
.A2(n_558),
.B1(n_584),
.B2(n_585),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_585),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_568),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_568),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_558),
.B(n_559),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_588),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_564),
.B(n_558),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_576),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_552),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_552),
.B(n_571),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_620),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_602),
.B(n_587),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_620),
.Y(n_632)
);

OR2x6_ASAP7_75t_SL g633 ( 
.A(n_616),
.B(n_573),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_603),
.B(n_552),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_616),
.A2(n_581),
.B1(n_578),
.B2(n_576),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_591),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_597),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_602),
.B(n_565),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_SL g640 ( 
.A1(n_598),
.A2(n_565),
.B(n_583),
.C(n_569),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_589),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_603),
.B(n_569),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_601),
.B(n_574),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_592),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_628),
.B(n_583),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_589),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_614),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_590),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_614),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_576),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_600),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_599),
.B(n_574),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_602),
.B(n_573),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_623),
.B(n_582),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_602),
.B(n_555),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_596),
.B(n_555),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_594),
.B(n_596),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_607),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_626),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_626),
.B(n_610),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_610),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_594),
.B(n_605),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_605),
.B(n_619),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_629),
.B(n_595),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_617),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_635),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_651),
.B(n_617),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_662),
.B(n_595),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_639),
.B(n_629),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_658),
.B(n_660),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_634),
.B(n_595),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_643),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_641),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_637),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_657),
.B(n_611),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_659),
.B(n_606),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_634),
.B(n_612),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_657),
.B(n_611),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_644),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_652),
.B(n_665),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_641),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_664),
.B(n_611),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_638),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_664),
.B(n_612),
.Y(n_684)
);

AND3x2_ASAP7_75t_L g685 ( 
.A(n_655),
.B(n_613),
.C(n_615),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_630),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_639),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_646),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_632),
.Y(n_689)
);

OAI21xp33_ASAP7_75t_L g690 ( 
.A1(n_656),
.A2(n_593),
.B(n_606),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_645),
.B(n_624),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_646),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_648),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_645),
.B(n_625),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_682),
.B(n_642),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_682),
.B(n_642),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_670),
.B(n_667),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_687),
.B(n_639),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_673),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_666),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_674),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_687),
.B(n_653),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_684),
.B(n_655),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_687),
.B(n_653),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_680),
.B(n_663),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_683),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_673),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_679),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_684),
.B(n_655),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_686),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_671),
.B(n_668),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_689),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_681),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_695),
.B(n_669),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_SL g715 ( 
.A(n_702),
.B(n_685),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_699),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_698),
.A2(n_690),
.B1(n_653),
.B2(n_631),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_697),
.A2(n_633),
.B1(n_672),
.B2(n_677),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_705),
.B(n_677),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_700),
.B(n_636),
.C(n_676),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_695),
.B(n_669),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_702),
.B(n_654),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_701),
.B(n_693),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_707),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_715),
.A2(n_633),
.B1(n_704),
.B2(n_711),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_SL g726 ( 
.A1(n_718),
.A2(n_703),
.B1(n_709),
.B2(n_698),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_723),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_SL g728 ( 
.A1(n_717),
.A2(n_704),
.B(n_698),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_716),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_719),
.B(n_706),
.Y(n_730)
);

OAI211xp5_ASAP7_75t_L g731 ( 
.A1(n_726),
.A2(n_720),
.B(n_706),
.C(n_718),
.Y(n_731)
);

AOI322xp5_ASAP7_75t_L g732 ( 
.A1(n_725),
.A2(n_722),
.A3(n_696),
.B1(n_721),
.B2(n_714),
.C1(n_724),
.C2(n_712),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_728),
.A2(n_710),
.B(n_708),
.Y(n_733)
);

OAI221xp5_ASAP7_75t_L g734 ( 
.A1(n_730),
.A2(n_707),
.B1(n_713),
.B2(n_699),
.C(n_671),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_SL g735 ( 
.A(n_727),
.B(n_652),
.C(n_713),
.Y(n_735)
);

AOI21xp33_ASAP7_75t_L g736 ( 
.A1(n_729),
.A2(n_631),
.B(n_692),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_736),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_SL g738 ( 
.A1(n_731),
.A2(n_733),
.B(n_735),
.Y(n_738)
);

NOR2x1_ASAP7_75t_SL g739 ( 
.A(n_732),
.B(n_639),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_734),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_731),
.A2(n_631),
.B(n_640),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_738),
.B(n_604),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_740),
.B(n_696),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_741),
.B(n_604),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_742),
.B(n_737),
.C(n_739),
.Y(n_745)
);

BUFx8_ASAP7_75t_SL g746 ( 
.A(n_744),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_743),
.B(n_737),
.C(n_627),
.Y(n_747)
);

NAND3x1_ASAP7_75t_L g748 ( 
.A(n_746),
.B(n_649),
.C(n_647),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_747),
.B(n_669),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_745),
.B(n_650),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_747),
.B(n_650),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_747),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_752),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_748),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_750),
.A2(n_749),
.B1(n_751),
.B2(n_627),
.Y(n_755)
);

NOR2x1_ASAP7_75t_L g756 ( 
.A(n_750),
.B(n_621),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_752),
.B(n_675),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_753),
.A2(n_618),
.B1(n_609),
.B2(n_621),
.Y(n_758)
);

AOI222xp33_ASAP7_75t_L g759 ( 
.A1(n_754),
.A2(n_640),
.B1(n_593),
.B2(n_661),
.C1(n_663),
.C2(n_606),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_756),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_757),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_755),
.A2(n_688),
.B(n_681),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_760),
.Y(n_763)
);

AOI21xp33_ASAP7_75t_SL g764 ( 
.A1(n_758),
.A2(n_622),
.B(n_615),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_762),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_763),
.B(n_759),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_SL g768 ( 
.A1(n_765),
.A2(n_604),
.B1(n_621),
.B2(n_608),
.Y(n_768)
);

AOI211x1_ASAP7_75t_L g769 ( 
.A1(n_766),
.A2(n_694),
.B(n_691),
.C(n_678),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_764),
.A2(n_622),
.B1(n_597),
.B2(n_608),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_767),
.A2(n_608),
.B(n_597),
.Y(n_771)
);

OA21x2_ASAP7_75t_L g772 ( 
.A1(n_771),
.A2(n_770),
.B(n_768),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_772),
.B(n_769),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_773),
.A2(n_593),
.B(n_618),
.Y(n_774)
);


endmodule