module fake_jpeg_18192_n_165 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_33),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_R g43 ( 
.A(n_39),
.B(n_27),
.Y(n_43)
);

OR2x2_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_48),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_51),
.B1(n_18),
.B2(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_27),
.B(n_28),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_59),
.C(n_32),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_23),
.B1(n_28),
.B2(n_19),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_61),
.B1(n_17),
.B2(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_15),
.Y(n_64)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_21),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_29),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_70),
.B1(n_4),
.B2(n_8),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_33),
.B1(n_37),
.B2(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_63),
.A2(n_77),
.B1(n_81),
.B2(n_10),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_15),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_74),
.B(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_71),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_20),
.B1(n_37),
.B2(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_54),
.B(n_47),
.C(n_50),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_29),
.B1(n_38),
.B2(n_5),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_80),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_36),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_59),
.B(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_29),
.B1(n_32),
.B2(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_13),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_85),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_33),
.C(n_32),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_59),
.C(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_14),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_96),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_47),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_84),
.C(n_62),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_46),
.C(n_47),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_57),
.C(n_8),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_63),
.B1(n_68),
.B2(n_79),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_4),
.B(n_9),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_105),
.B(n_95),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_9),
.B(n_10),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_86),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_112),
.B(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_119),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_78),
.B(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_95),
.B(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_108),
.B1(n_99),
.B2(n_98),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_103),
.C(n_90),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_131),
.C(n_110),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_123),
.B1(n_124),
.B2(n_117),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_103),
.C(n_100),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_103),
.B(n_105),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_140),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_115),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_144),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_124),
.B1(n_119),
.B2(n_117),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_128),
.C(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_142),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_148),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_141),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_127),
.B(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_133),
.Y(n_152)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_110),
.A3(n_101),
.B1(n_134),
.B2(n_130),
.C(n_114),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_130),
.A3(n_115),
.B1(n_137),
.B2(n_96),
.C1(n_143),
.C2(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_156),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_147),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_102),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.C(n_154),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

AOI31xp67_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_152),
.A3(n_149),
.B(n_102),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_159),
.C(n_160),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_79),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);


endmodule