module real_jpeg_14836_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_3),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_3),
.A2(n_61),
.B(n_64),
.C(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_103),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_30),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_SL g232 ( 
.A1(n_3),
.A2(n_30),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_3),
.B(n_47),
.C(n_52),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_3),
.A2(n_33),
.B1(n_37),
.B2(n_158),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_3),
.A2(n_87),
.B1(n_88),
.B2(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_3),
.B(n_42),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_33),
.B1(n_37),
.B2(n_165),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_165),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_6),
.A2(n_33),
.B1(n_37),
.B2(n_68),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_68),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_27),
.B1(n_64),
.B2(n_65),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_7),
.A2(n_27),
.B1(n_51),
.B2(n_52),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_9),
.A2(n_33),
.B1(n_37),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_57),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_11),
.A2(n_41),
.B1(n_64),
.B2(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_11),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_11),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_13),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_13),
.A2(n_33),
.B1(n_37),
.B2(n_161),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_161),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_14),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_33),
.B1(n_37),
.B2(n_147),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_147),
.Y(n_249)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_19),
.B(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.C(n_85),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_20),
.B(n_75),
.CI(n_85),
.CON(n_149),
.SN(n_149)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_59),
.B2(n_74),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_43),
.B2(n_58),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_23),
.B(n_58),
.C(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_26),
.A2(n_42),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_28),
.A2(n_30),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_SL g219 ( 
.A(n_28),
.B(n_35),
.C(n_37),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_30),
.A2(n_62),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_31),
.A2(n_32),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_31),
.A2(n_32),
.B1(n_164),
.B2(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_31),
.A2(n_113),
.B(n_166),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_31),
.A2(n_32),
.B1(n_186),
.B2(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_31),
.A2(n_39),
.B(n_115),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_32),
.A2(n_83),
.B(n_116),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx5_ASAP7_75t_SL g37 ( 
.A(n_33),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_33),
.A2(n_36),
.B(n_217),
.C(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_33),
.B(n_241),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_40),
.B(n_84),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_42),
.B(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_43),
.A2(n_58),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_50),
.B(n_55),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_44),
.A2(n_55),
.B(n_97),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_44),
.A2(n_77),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_45),
.A2(n_78),
.B1(n_95),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_45),
.A2(n_78),
.B1(n_213),
.B2(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_45),
.A2(n_78),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_45),
.A2(n_78),
.B1(n_234),
.B2(n_244),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_50),
.A2(n_79),
.B(n_143),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_50),
.B(n_158),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_51),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_88),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_78),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_74),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_69),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_63),
.B1(n_71),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_60),
.A2(n_71),
.B1(n_160),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_60),
.A2(n_71),
.B1(n_146),
.B2(n_191),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_72)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_70),
.A2(n_103),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_71),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_76),
.B(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B(n_98),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_98),
.B1(n_99),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_86),
.A2(n_93),
.B1(n_94),
.B2(n_128),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_90),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_87),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_87),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_87),
.A2(n_88),
.B1(n_247),
.B2(n_255),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_87),
.A2(n_137),
.B(n_249),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_88),
.B(n_139),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_88),
.B(n_158),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_91),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_89),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_89),
.A2(n_138),
.B(n_175),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_89),
.A2(n_174),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_91),
.A2(n_174),
.B(n_200),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_103),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_150),
.B(n_312),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_149),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_125),
.B(n_149),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_130),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_126),
.B(n_129),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_130),
.A2(n_131),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_144),
.C(n_145),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_132),
.A2(n_133),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_141),
.Y(n_284)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_144),
.B(n_145),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_149),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_306),
.B(n_311),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_294),
.B(n_305),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_202),
.B(n_280),
.C(n_293),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_187),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_154),
.B(n_187),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_170),
.C(n_180),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_167),
.C(n_169),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_171),
.B1(n_180),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_177),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_185),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_188),
.B(n_195),
.C(n_201),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_190),
.B(n_192),
.C(n_193),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_196),
.B(n_197),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_278),
.B(n_279),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_222),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_205),
.B(n_208),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.C(n_214),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_214),
.B1(n_215),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_220),
.B1(n_221),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_235),
.B(n_277),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_227),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_233),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_271),
.B(n_276),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_261),
.B(n_270),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_250),
.B(n_260),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_245),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_242),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_256),
.B(n_259),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_266),
.C(n_269),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_292),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_292),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_288),
.C(n_291),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_304),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_302),
.B2(n_303),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_303),
.C(n_304),
.Y(n_310)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);


endmodule