module fake_netlist_6_4897_n_1168 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_58, n_116, n_280, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1168);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_58;
input n_116;
input n_280;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1168;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_760;
wire n_680;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1079;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_726;
wire n_671;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_1164;
wire n_310;
wire n_509;
wire n_575;
wire n_368;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_840;
wire n_392;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_1153;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_685;
wire n_597;
wire n_832;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_814;
wire n_389;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_826;
wire n_383;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_544;
wire n_372;
wire n_468;
wire n_1078;
wire n_923;
wire n_504;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1163;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_843;
wire n_772;
wire n_656;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_838;
wire n_380;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_559;
wire n_334;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_719;
wire n_565;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_527;
wire n_620;
wire n_683;
wire n_811;
wire n_630;
wire n_312;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_394;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_689;
wire n_345;
wire n_354;
wire n_799;
wire n_505;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_550;
wire n_487;
wire n_1125;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_1167;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_420;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_410;
wire n_398;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_59),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_122),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_94),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_78),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_274),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_129),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_197),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_88),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_3),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_191),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_107),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_185),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_135),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_235),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_193),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_97),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_48),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_112),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_85),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_246),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_242),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_64),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_84),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_267),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_170),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_101),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_213),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_249),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_9),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_90),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_272),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_27),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_123),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_109),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_82),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_121),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_167),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_92),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_67),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_130),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_276),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_245),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_47),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_34),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_163),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_98),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_127),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_181),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_243),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_68),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_244),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_211),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_166),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_3),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_224),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_160),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_142),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_136),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_232),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_83),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_113),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_137),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_132),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_271),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_119),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_273),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_5),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_268),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_171),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_217),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_23),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_204),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_46),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_50),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_143),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_174),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_169),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_116),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_161),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_222),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_206),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_149),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_157),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_240),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_187),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_16),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_93),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_80),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_205),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_200),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_199),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_151),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_96),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_100),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_120),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_165),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_270),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_38),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_214),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_41),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_216),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_190),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_125),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_52),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_57),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_262),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_89),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_49),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_139),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_275),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_43),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_263),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_172),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_45),
.Y(n_403)
);

BUFx10_ASAP7_75t_L g404 ( 
.A(n_202),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_51),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_104),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_105),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_55),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_77),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_65),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_2),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_30),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_178),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_141),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_17),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_54),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_73),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_108),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_39),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_150),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_76),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_145),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_261),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_35),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_210),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_277),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_266),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_6),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_148),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_256),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_24),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_6),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_8),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_66),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_26),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_159),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_252),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_221),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_195),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_32),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_279),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_115),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_180),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_248),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_265),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_175),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_37),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_15),
.Y(n_448)
);

BUFx2_ASAP7_75t_SL g449 ( 
.A(n_146),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_201),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_114),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_15),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_238),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_212),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_218),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_56),
.Y(n_456)
);

BUFx5_ASAP7_75t_L g457 ( 
.A(n_12),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_138),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_278),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_457),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_296),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_457),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_457),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_305),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_290),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_324),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_343),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_285),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_287),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_288),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_289),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_294),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_282),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_291),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_292),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_297),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_332),
.B(n_0),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_295),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_319),
.B(n_0),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_284),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_428),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_301),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_286),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_303),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_419),
.B(n_1),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_298),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_333),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_300),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_448),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_307),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_418),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_308),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_299),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_309),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_311),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_376),
.B(n_1),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_317),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_304),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_306),
.Y(n_503)
);

INVxp33_ASAP7_75t_SL g504 ( 
.A(n_302),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_325),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_310),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_312),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_293),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_326),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_370),
.B(n_2),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_327),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_342),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_328),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_331),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_443),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_315),
.B(n_4),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_338),
.Y(n_518)
);

INVxp33_ASAP7_75t_SL g519 ( 
.A(n_356),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_339),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_344),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_360),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_348),
.B(n_4),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_346),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_350),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_369),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_314),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_316),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_353),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_318),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_283),
.B(n_5),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_321),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_372),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_362),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_313),
.B(n_7),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_415),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_363),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_381),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_393),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_395),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_322),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_335),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_378),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_293),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_323),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_397),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_379),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_451),
.B(n_320),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_403),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_407),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_382),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_412),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_384),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_414),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_422),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_329),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_391),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_425),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_434),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_545),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_468),
.B(n_367),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_509),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_491),
.B(n_385),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_471),
.B(n_387),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_509),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_461),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_466),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_475),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_478),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_466),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_479),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_549),
.A2(n_438),
.B(n_437),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_462),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_463),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_488),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_543),
.B(n_409),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_469),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_474),
.B(n_427),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_543),
.B(n_440),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_476),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_480),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_472),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_490),
.B(n_447),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_494),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_523),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_496),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_492),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_501),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_524),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_510),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_522),
.B(n_335),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_504),
.B(n_373),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_502),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_512),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_503),
.B(n_456),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_507),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_562),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_514),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_485),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_515),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_561),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_493),
.A2(n_452),
.B1(n_432),
.B2(n_431),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_528),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_518),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_520),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_525),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_526),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_530),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_535),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_538),
.B(n_293),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_539),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_537),
.B(n_459),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_540),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_541),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_547),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_529),
.B(n_458),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_551),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_560),
.B(n_405),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_553),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_516),
.B(n_361),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_555),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_556),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_559),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_465),
.B(n_361),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_483),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_481),
.B(n_433),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_519),
.B(n_453),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_517),
.B(n_337),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_495),
.B(n_400),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_464),
.B(n_400),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_477),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_506),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_511),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_610),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_631),
.A2(n_489),
.B1(n_500),
.B2(n_532),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_638),
.B(n_531),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_570),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_533),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_563),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_624),
.A2(n_489),
.B1(n_500),
.B2(n_532),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_602),
.B(n_542),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_585),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_590),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_564),
.B(n_546),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_574),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_590),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_585),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_585),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_571),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_567),
.B(n_557),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_598),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_571),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_624),
.A2(n_536),
.B1(n_467),
.B2(n_470),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_571),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_598),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_581),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_572),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_644),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_572),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_572),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_573),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_638),
.B(n_646),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_608),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_638),
.B(n_330),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_598),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_637),
.B(n_467),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_609),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_611),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_633),
.B(n_337),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_601),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_576),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_646),
.B(n_337),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_582),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_575),
.Y(n_689)
);

INVxp67_ASAP7_75t_SL g690 ( 
.A(n_576),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_577),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_578),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_576),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_645),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_579),
.Y(n_695)
);

BUFx4_ASAP7_75t_L g696 ( 
.A(n_591),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_588),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_586),
.B(n_536),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_640),
.B(n_558),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_599),
.B(n_470),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_646),
.A2(n_449),
.B1(n_349),
.B2(n_377),
.Y(n_701)
);

INVx6_ASAP7_75t_L g702 ( 
.A(n_584),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_611),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_593),
.B(n_334),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_611),
.Y(n_705)
);

NAND2x1p5_ASAP7_75t_L g706 ( 
.A(n_614),
.B(n_349),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_593),
.Y(n_707)
);

NOR2x1p5_ASAP7_75t_L g708 ( 
.A(n_615),
.B(n_336),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_595),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_595),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_612),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_632),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_607),
.B(n_484),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_605),
.B(n_554),
.Y(n_714)
);

INVx6_ASAP7_75t_L g715 ( 
.A(n_584),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_587),
.Y(n_716)
);

NAND2x1p5_ASAP7_75t_L g717 ( 
.A(n_589),
.B(n_349),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_600),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_600),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_593),
.B(n_340),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_617),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_629),
.B(n_487),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_596),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_616),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_632),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_566),
.A2(n_377),
.B1(n_390),
.B2(n_446),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_628),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_632),
.Y(n_728)
);

NOR2x1p5_ASAP7_75t_L g729 ( 
.A(n_650),
.B(n_587),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_698),
.A2(n_639),
.B1(n_566),
.B2(n_421),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_652),
.A2(n_424),
.B1(n_406),
.B2(n_603),
.Y(n_731)
);

AO22x2_ASAP7_75t_L g732 ( 
.A1(n_681),
.A2(n_642),
.B1(n_643),
.B2(n_641),
.Y(n_732)
);

AO22x2_ASAP7_75t_L g733 ( 
.A1(n_700),
.A2(n_647),
.B1(n_655),
.B2(n_713),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_677),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_709),
.Y(n_735)
);

XOR2xp5_ASAP7_75t_L g736 ( 
.A(n_723),
.B(n_497),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_709),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_694),
.B(n_673),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_699),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_660),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_707),
.B(n_606),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_714),
.Y(n_742)
);

OAI221xp5_ASAP7_75t_L g743 ( 
.A1(n_649),
.A2(n_620),
.B1(n_617),
.B2(n_618),
.C(n_619),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_685),
.A2(n_641),
.B1(n_513),
.B2(n_521),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_653),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_659),
.B(n_499),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_654),
.A2(n_619),
.B1(n_620),
.B2(n_618),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_710),
.A2(n_592),
.B1(n_594),
.B2(n_583),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_657),
.B(n_621),
.Y(n_749)
);

AND2x2_ASAP7_75t_SL g750 ( 
.A(n_722),
.B(n_527),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_678),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_665),
.B(n_580),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_710),
.Y(n_753)
);

AO22x2_ASAP7_75t_L g754 ( 
.A1(n_718),
.A2(n_534),
.B1(n_544),
.B2(n_548),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_679),
.B(n_552),
.Y(n_755)
);

AO22x2_ASAP7_75t_L g756 ( 
.A1(n_718),
.A2(n_613),
.B1(n_8),
.B2(n_10),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_682),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_719),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_676),
.A2(n_580),
.B1(n_635),
.B2(n_634),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_719),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_721),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_721),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_711),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_648),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_668),
.A2(n_651),
.B1(n_648),
.B2(n_689),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_651),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_691),
.A2(n_623),
.B1(n_625),
.B2(n_626),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_692),
.Y(n_768)
);

AO22x2_ASAP7_75t_L g769 ( 
.A1(n_695),
.A2(n_627),
.B1(n_10),
.B2(n_11),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_728),
.B(n_597),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_658),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_661),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_724),
.Y(n_773)
);

OAI221xp5_ASAP7_75t_L g774 ( 
.A1(n_726),
.A2(n_636),
.B1(n_630),
.B2(n_604),
.C(n_597),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_727),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_702),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_669),
.B(n_604),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_672),
.B(n_565),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_671),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_697),
.B(n_565),
.Y(n_780)
);

AND2x6_ASAP7_75t_L g781 ( 
.A(n_671),
.B(n_377),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_688),
.Y(n_782)
);

AO22x2_ASAP7_75t_L g783 ( 
.A1(n_696),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_688),
.Y(n_784)
);

OAI221xp5_ASAP7_75t_L g785 ( 
.A1(n_701),
.A2(n_408),
.B1(n_345),
.B2(n_347),
.C(n_351),
.Y(n_785)
);

AO22x2_ASAP7_75t_L g786 ( 
.A1(n_704),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_786)
);

AO22x2_ASAP7_75t_L g787 ( 
.A1(n_720),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_702),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_715),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_662),
.B(n_568),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_684),
.B(n_341),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_715),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_656),
.B(n_568),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_717),
.B(n_352),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_666),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_728),
.B(n_354),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_666),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_656),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_664),
.B(n_390),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_663),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_670),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_708),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_664),
.B(n_355),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_742),
.B(n_716),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_739),
.B(n_716),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_730),
.B(n_728),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_738),
.B(n_667),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_SL g808 ( 
.A(n_802),
.B(n_667),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_746),
.B(n_706),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_SL g810 ( 
.A(n_729),
.B(n_667),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_734),
.B(n_780),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_SL g812 ( 
.A(n_788),
.B(n_674),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_755),
.B(n_674),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_731),
.B(n_674),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_750),
.B(n_675),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_768),
.B(n_675),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_735),
.B(n_737),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_753),
.B(n_675),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_SL g819 ( 
.A(n_789),
.B(n_686),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_758),
.B(n_686),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_760),
.B(n_761),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_762),
.B(n_686),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_792),
.B(n_690),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_764),
.B(n_693),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_766),
.B(n_693),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_771),
.B(n_693),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_772),
.B(n_712),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_784),
.B(n_712),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_741),
.B(n_725),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_SL g830 ( 
.A(n_776),
.B(n_725),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_752),
.B(n_684),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_779),
.B(n_670),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_782),
.B(n_680),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_794),
.B(n_680),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_765),
.B(n_683),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_759),
.B(n_683),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_765),
.B(n_749),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_778),
.B(n_703),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_751),
.B(n_703),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_796),
.B(n_705),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_757),
.B(n_705),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_SL g842 ( 
.A(n_770),
.B(n_357),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_747),
.B(n_684),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_747),
.B(n_684),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_740),
.B(n_663),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_SL g846 ( 
.A(n_795),
.B(n_358),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_763),
.B(n_359),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_SL g848 ( 
.A(n_797),
.B(n_364),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_773),
.B(n_365),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_745),
.B(n_687),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_SL g851 ( 
.A(n_801),
.B(n_366),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_733),
.B(n_687),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_798),
.B(n_390),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_SL g854 ( 
.A1(n_844),
.A2(n_785),
.B(n_793),
.C(n_790),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_836),
.A2(n_800),
.B(n_775),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_831),
.A2(n_803),
.B(n_791),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_817),
.A2(n_777),
.B(n_799),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_806),
.A2(n_743),
.B(n_774),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_821),
.A2(n_733),
.B1(n_732),
.B2(n_748),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_850),
.A2(n_845),
.B(n_833),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_807),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_835),
.B(n_809),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_814),
.A2(n_732),
.B(n_748),
.C(n_368),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_839),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_837),
.B(n_823),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_823),
.B(n_767),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_811),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_832),
.A2(n_767),
.B(n_687),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_843),
.A2(n_687),
.B(n_781),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_852),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_829),
.B(n_446),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_815),
.B(n_446),
.Y(n_872)
);

INVx6_ASAP7_75t_L g873 ( 
.A(n_808),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_828),
.A2(n_781),
.B(n_29),
.Y(n_874)
);

AOI211x1_ASAP7_75t_L g875 ( 
.A1(n_818),
.A2(n_769),
.B(n_786),
.C(n_787),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_841),
.Y(n_876)
);

AO21x1_ASAP7_75t_L g877 ( 
.A1(n_840),
.A2(n_769),
.B(n_756),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_810),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_805),
.B(n_736),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_804),
.B(n_371),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_838),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_820),
.A2(n_781),
.B(n_31),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_834),
.A2(n_813),
.B(n_827),
.Y(n_883)
);

NAND3xp33_ASAP7_75t_L g884 ( 
.A(n_849),
.B(n_848),
.C(n_846),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_851),
.Y(n_885)
);

O2A1O1Ixp5_ASAP7_75t_SL g886 ( 
.A1(n_853),
.A2(n_744),
.B(n_754),
.C(n_783),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_822),
.A2(n_380),
.B(n_374),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_877),
.A2(n_825),
.B1(n_824),
.B2(n_826),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_866),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_859),
.A2(n_816),
.B1(n_404),
.B2(n_830),
.Y(n_890)
);

OA21x2_ASAP7_75t_L g891 ( 
.A1(n_863),
.A2(n_853),
.B(n_847),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_862),
.B(n_842),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_855),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_865),
.A2(n_417),
.B1(n_386),
.B2(n_455),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_860),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_SL g896 ( 
.A(n_873),
.B(n_383),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_864),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_870),
.B(n_404),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_861),
.B(n_819),
.Y(n_899)
);

OAI21x1_ASAP7_75t_SL g900 ( 
.A1(n_883),
.A2(n_812),
.B(n_33),
.Y(n_900)
);

AO21x2_ASAP7_75t_L g901 ( 
.A1(n_856),
.A2(n_622),
.B(n_389),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_864),
.Y(n_902)
);

AND2x2_ASAP7_75t_SL g903 ( 
.A(n_878),
.B(n_18),
.Y(n_903)
);

BUFx8_ASAP7_75t_L g904 ( 
.A(n_867),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_854),
.A2(n_392),
.B(n_388),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_884),
.A2(n_396),
.B(n_394),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_875),
.B(n_28),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_858),
.A2(n_426),
.B1(n_454),
.B2(n_450),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_878),
.Y(n_909)
);

AOI21x1_ASAP7_75t_L g910 ( 
.A1(n_868),
.A2(n_622),
.B(n_445),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_858),
.A2(n_420),
.B1(n_444),
.B2(n_442),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_874),
.A2(n_182),
.B(n_281),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_876),
.A2(n_416),
.B(n_441),
.Y(n_913)
);

OA21x2_ASAP7_75t_L g914 ( 
.A1(n_882),
.A2(n_413),
.B(n_439),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_880),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_876),
.Y(n_916)
);

AOI221xp5_ASAP7_75t_L g917 ( 
.A1(n_875),
.A2(n_881),
.B1(n_885),
.B2(n_879),
.C(n_887),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_897),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_897),
.B(n_872),
.Y(n_919)
);

INVxp33_ASAP7_75t_L g920 ( 
.A(n_898),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_916),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_916),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_904),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_902),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_895),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_909),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_889),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_915),
.B(n_871),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_909),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_909),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_909),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_899),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_SL g933 ( 
.A1(n_907),
.A2(n_892),
.B(n_891),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_907),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_903),
.B(n_886),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_895),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_907),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_907),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_904),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_903),
.B(n_873),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_917),
.B(n_869),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_893),
.A2(n_857),
.B(n_177),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_893),
.Y(n_943)
);

AO22x1_ASAP7_75t_L g944 ( 
.A1(n_904),
.A2(n_410),
.B1(n_430),
.B2(n_429),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_908),
.A2(n_622),
.B(n_423),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_908),
.A2(n_402),
.B1(n_401),
.B2(n_399),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_911),
.B(n_36),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_912),
.A2(n_164),
.B(n_280),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_912),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_900),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_891),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_906),
.Y(n_952)
);

BUFx10_ASAP7_75t_L g953 ( 
.A(n_940),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_932),
.Y(n_954)
);

NAND2xp33_ASAP7_75t_R g955 ( 
.A(n_940),
.B(n_923),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_924),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_927),
.B(n_911),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_929),
.B(n_888),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_935),
.B(n_890),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_SL g960 ( 
.A(n_947),
.B(n_896),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_918),
.B(n_921),
.Y(n_961)
);

BUFx4f_ASAP7_75t_L g962 ( 
.A(n_930),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_928),
.B(n_910),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_935),
.B(n_890),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_931),
.B(n_888),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_930),
.B(n_398),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_922),
.B(n_891),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_930),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_926),
.B(n_913),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_920),
.B(n_894),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_939),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_930),
.Y(n_972)
);

XOR2xp5_ASAP7_75t_L g973 ( 
.A(n_920),
.B(n_905),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_943),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_R g975 ( 
.A(n_952),
.B(n_914),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_SL g976 ( 
.A(n_947),
.B(n_901),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_919),
.B(n_901),
.Y(n_977)
);

XOR2xp5_ASAP7_75t_L g978 ( 
.A(n_944),
.B(n_946),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_926),
.B(n_40),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_943),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_934),
.B(n_914),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_925),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_919),
.B(n_914),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_941),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_R g985 ( 
.A(n_926),
.B(n_42),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_937),
.B(n_53),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_938),
.B(n_58),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_950),
.B(n_60),
.Y(n_988)
);

AND2x2_ASAP7_75t_SL g989 ( 
.A(n_946),
.B(n_951),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_933),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_956),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_954),
.B(n_933),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_977),
.B(n_925),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_983),
.B(n_936),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_961),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_974),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_980),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_967),
.B(n_936),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_982),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_981),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_958),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_958),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_965),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_965),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_959),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_968),
.B(n_949),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_968),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_972),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_964),
.B(n_949),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_989),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_970),
.B(n_949),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_962),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_976),
.B(n_942),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_957),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_978),
.A2(n_945),
.B1(n_948),
.B2(n_942),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_953),
.B(n_948),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_953),
.B(n_18),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_973),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_969),
.B(n_19),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_969),
.B(n_19),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_997),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_1008),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_1011),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_991),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_995),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_1000),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_1001),
.B(n_1011),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_1000),
.B(n_960),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1005),
.B(n_971),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_997),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_1008),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_996),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1005),
.B(n_986),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1009),
.B(n_987),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_1010),
.A2(n_1015),
.B(n_986),
.C(n_990),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1009),
.Y(n_1036)
);

AOI322xp5_ASAP7_75t_L g1037 ( 
.A1(n_1010),
.A2(n_955),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_24),
.C2(n_25),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_999),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1002),
.B(n_968),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1004),
.B(n_966),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_992),
.B(n_975),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1030),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_L g1043 ( 
.A(n_1031),
.B(n_1014),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1026),
.B(n_994),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1036),
.B(n_1018),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1021),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1021),
.Y(n_1047)
);

AO21x1_ASAP7_75t_L g1048 ( 
.A1(n_1041),
.A2(n_1020),
.B(n_1019),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1036),
.B(n_1001),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_1031),
.B(n_1006),
.Y(n_1050)
);

OR2x6_ASAP7_75t_SL g1051 ( 
.A(n_1033),
.B(n_1003),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1038),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1040),
.B(n_1017),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_1027),
.B(n_993),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1027),
.B(n_993),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1026),
.B(n_994),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1023),
.B(n_993),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_1023),
.B(n_998),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1025),
.B(n_998),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1034),
.B(n_1016),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1042),
.Y(n_1061)
);

OAI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1053),
.A2(n_1035),
.B1(n_1037),
.B2(n_1028),
.C(n_1017),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_1043),
.B(n_1022),
.Y(n_1063)
);

OAI221xp5_ASAP7_75t_L g1064 ( 
.A1(n_1050),
.A2(n_1035),
.B1(n_1019),
.B2(n_1020),
.C(n_1024),
.Y(n_1064)
);

AO221x2_ASAP7_75t_L g1065 ( 
.A1(n_1048),
.A2(n_1032),
.B1(n_1029),
.B2(n_1022),
.C(n_988),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1060),
.B(n_1039),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1045),
.B(n_1022),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_1059),
.Y(n_1068)
);

AO221x2_ASAP7_75t_L g1069 ( 
.A1(n_1052),
.A2(n_1022),
.B1(n_21),
.B2(n_22),
.C(n_25),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1054),
.A2(n_1016),
.B1(n_1012),
.B2(n_1007),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_1059),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_1051),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_1054),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1044),
.B(n_1013),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1044),
.B(n_1013),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1047),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1056),
.B(n_1006),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1056),
.B(n_1006),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1065),
.A2(n_1050),
.B1(n_1057),
.B2(n_1055),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1071),
.B(n_1058),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1061),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_1065),
.A2(n_963),
.B1(n_985),
.B2(n_979),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_L g1083 ( 
.A(n_1062),
.B(n_1012),
.C(n_1007),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1076),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_1068),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1069),
.A2(n_1049),
.B1(n_1046),
.B2(n_622),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_1063),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1073),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_1072),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1067),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1074),
.B(n_20),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_1077),
.Y(n_1092)
);

AOI21xp33_ASAP7_75t_L g1093 ( 
.A1(n_1064),
.A2(n_20),
.B(n_61),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1066),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1078),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1070),
.B(n_62),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1075),
.B(n_63),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1069),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1072),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1072),
.B(n_69),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1081),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1083),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_1080),
.B(n_74),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1083),
.A2(n_75),
.B1(n_79),
.B2(n_81),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1087),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1084),
.Y(n_1106)
);

OAI332xp33_ASAP7_75t_L g1107 ( 
.A1(n_1089),
.A2(n_86),
.A3(n_87),
.B1(n_91),
.B2(n_95),
.B3(n_99),
.C1(n_102),
.C2(n_103),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1099),
.B(n_106),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1091),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1098),
.A2(n_110),
.B(n_111),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1098),
.A2(n_117),
.B(n_118),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1095),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1082),
.A2(n_1086),
.B1(n_1079),
.B2(n_1085),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1092),
.B(n_124),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1109),
.B(n_1100),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1110),
.A2(n_1093),
.B1(n_1090),
.B2(n_1088),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1106),
.B(n_1094),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1113),
.B(n_1093),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1101),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1112),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1105),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1111),
.A2(n_1097),
.B1(n_1096),
.B2(n_131),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1103),
.B(n_126),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_1114),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1108),
.B(n_128),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1102),
.B(n_133),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1104),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1107),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_L g1129 ( 
.A(n_1107),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1121),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1115),
.B(n_134),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_1124),
.Y(n_1132)
);

XOR2xp5_ASAP7_75t_L g1133 ( 
.A(n_1122),
.B(n_140),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1119),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1123),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1117),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1117),
.Y(n_1137)
);

INVxp67_ASAP7_75t_SL g1138 ( 
.A(n_1118),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1138),
.B(n_1128),
.C(n_1127),
.Y(n_1139)
);

NAND4xp75_ASAP7_75t_L g1140 ( 
.A(n_1136),
.B(n_1129),
.C(n_1120),
.D(n_1126),
.Y(n_1140)
);

OAI211xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1138),
.A2(n_1116),
.B(n_1125),
.C(n_152),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_1130),
.B(n_144),
.C(n_147),
.Y(n_1142)
);

OA211x2_ASAP7_75t_L g1143 ( 
.A1(n_1131),
.A2(n_153),
.B(n_154),
.C(n_155),
.Y(n_1143)
);

NOR3xp33_ASAP7_75t_L g1144 ( 
.A(n_1132),
.B(n_1135),
.C(n_1137),
.Y(n_1144)
);

O2A1O1Ixp5_ASAP7_75t_L g1145 ( 
.A1(n_1134),
.A2(n_156),
.B(n_158),
.C(n_162),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1139),
.A2(n_1133),
.B1(n_173),
.B2(n_176),
.C(n_179),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_1140),
.B(n_168),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_SL g1148 ( 
.A(n_1141),
.B(n_183),
.C(n_184),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1144),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.C(n_192),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1142),
.A2(n_1145),
.B(n_1143),
.Y(n_1150)
);

NAND4xp75_ASAP7_75t_L g1151 ( 
.A(n_1147),
.B(n_194),
.C(n_198),
.D(n_203),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1148),
.Y(n_1152)
);

NOR4xp25_ASAP7_75t_L g1153 ( 
.A(n_1146),
.B(n_207),
.C(n_208),
.D(n_209),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1153),
.B(n_1150),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_SL g1155 ( 
.A(n_1152),
.B(n_1149),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1154),
.Y(n_1156)
);

AOI222xp33_ASAP7_75t_L g1157 ( 
.A1(n_1155),
.A2(n_1151),
.B1(n_219),
.B2(n_220),
.C1(n_223),
.C2(n_225),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1156),
.A2(n_215),
.B1(n_226),
.B2(n_227),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1157),
.B(n_228),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1159),
.Y(n_1160)
);

AOI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1158),
.A2(n_229),
.B(n_230),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_1161),
.B1(n_233),
.B2(n_236),
.Y(n_1162)
);

AOI31xp33_ASAP7_75t_L g1163 ( 
.A1(n_1160),
.A2(n_231),
.A3(n_239),
.B(n_241),
.Y(n_1163)
);

XOR2xp5_ASAP7_75t_L g1164 ( 
.A(n_1162),
.B(n_247),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1164),
.A2(n_1163),
.B(n_251),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_1165),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1166),
.A2(n_250),
.B1(n_254),
.B2(n_255),
.C(n_257),
.Y(n_1167)
);

AOI211xp5_ASAP7_75t_L g1168 ( 
.A1(n_1167),
.A2(n_258),
.B(n_259),
.C(n_260),
.Y(n_1168)
);


endmodule