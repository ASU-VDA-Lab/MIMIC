module real_aes_11043_n_266 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_266);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_266;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1457;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_0), .A2(n_37), .B1(n_441), .B2(n_442), .C(n_633), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_0), .A2(n_259), .B1(n_460), .B2(n_464), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g1173 ( .A(n_1), .Y(n_1173) );
XNOR2xp5_ASAP7_75t_L g293 ( .A(n_2), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g1276 ( .A(n_3), .Y(n_1276) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_4), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_5), .A2(n_70), .B1(n_556), .B2(n_888), .Y(n_1063) );
INVx1_ASAP7_75t_L g1089 ( .A(n_5), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_6), .A2(n_254), .B1(n_480), .B2(n_1141), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_6), .A2(n_254), .B1(n_937), .B2(n_1148), .Y(n_1147) );
XNOR2xp5_ASAP7_75t_L g695 ( .A(n_7), .B(n_696), .Y(n_695) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_8), .Y(n_1189) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_9), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_9), .B(n_200), .Y(n_382) );
AND2x2_ASAP7_75t_L g390 ( .A(n_9), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g445 ( .A(n_9), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g1113 ( .A(n_10), .Y(n_1113) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_11), .A2(n_180), .B1(n_359), .B2(n_365), .Y(n_358) );
INVx1_ASAP7_75t_L g447 ( .A(n_11), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_12), .A2(n_92), .B1(n_467), .B2(n_469), .Y(n_719) );
INVx1_ASAP7_75t_L g738 ( .A(n_12), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g1188 ( .A(n_13), .Y(n_1188) );
INVx1_ASAP7_75t_L g599 ( .A(n_14), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_14), .A2(n_75), .B1(n_388), .B2(n_396), .Y(n_608) );
INVx1_ASAP7_75t_L g1311 ( .A(n_15), .Y(n_1311) );
INVx1_ASAP7_75t_L g708 ( .A(n_16), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_17), .A2(n_226), .B1(n_440), .B2(n_441), .C(n_442), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_17), .A2(n_85), .B1(n_467), .B2(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g851 ( .A(n_18), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_18), .A2(n_197), .B1(n_890), .B2(n_891), .Y(n_889) );
XNOR2xp5_ASAP7_75t_L g893 ( .A(n_19), .B(n_894), .Y(n_893) );
AO221x2_ASAP7_75t_L g1246 ( .A1(n_19), .A2(n_54), .B1(n_1230), .B2(n_1239), .C(n_1247), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_20), .A2(n_208), .B1(n_484), .B2(n_487), .C(n_490), .Y(n_483) );
INVx1_ASAP7_75t_L g516 ( .A(n_20), .Y(n_516) );
INVx1_ASAP7_75t_L g1264 ( .A(n_21), .Y(n_1264) );
INVx2_ASAP7_75t_L g309 ( .A(n_22), .Y(n_309) );
OR2x2_ASAP7_75t_L g463 ( .A(n_22), .B(n_307), .Y(n_463) );
INVx1_ASAP7_75t_L g1248 ( .A(n_23), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_24), .A2(n_218), .B1(n_890), .B2(n_891), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_24), .A2(n_218), .B1(n_396), .B2(n_670), .Y(n_1094) );
INVx1_ASAP7_75t_L g311 ( .A(n_25), .Y(n_311) );
BUFx2_ASAP7_75t_L g318 ( .A(n_25), .Y(n_318) );
BUFx2_ASAP7_75t_L g356 ( .A(n_25), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g981 ( .A1(n_26), .A2(n_192), .B1(n_508), .B2(n_921), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_26), .A2(n_192), .B1(n_563), .B2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g907 ( .A(n_27), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_27), .A2(n_191), .B1(n_919), .B2(n_921), .Y(n_918) );
INVx1_ASAP7_75t_L g1309 ( .A(n_28), .Y(n_1309) );
INVx1_ASAP7_75t_L g349 ( .A(n_29), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_29), .A2(n_72), .B1(n_388), .B2(n_396), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_30), .A2(n_108), .B1(n_819), .B2(n_911), .Y(n_1165) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_30), .A2(n_108), .B1(n_441), .B2(n_505), .C(n_633), .Y(n_1183) );
OAI22xp33_ASAP7_75t_L g974 ( .A1(n_31), .A2(n_60), .B1(n_281), .B2(n_860), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_31), .A2(n_164), .B1(n_990), .B2(n_991), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_32), .A2(n_55), .B1(n_503), .B2(n_504), .C(n_505), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_32), .A2(n_55), .B1(n_552), .B2(n_556), .Y(n_551) );
INVx1_ASAP7_75t_L g1028 ( .A(n_33), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_33), .A2(n_58), .B1(n_467), .B2(n_469), .Y(n_1053) );
CKINVDCx16_ASAP7_75t_R g1261 ( .A(n_34), .Y(n_1261) );
INVx1_ASAP7_75t_L g438 ( .A(n_35), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_35), .A2(n_226), .B1(n_460), .B2(n_464), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_36), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_37), .A2(n_57), .B1(n_467), .B2(n_469), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_38), .A2(n_227), .B1(n_911), .B2(n_913), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_38), .A2(n_227), .B1(n_923), .B2(n_930), .Y(n_929) );
XNOR2xp5_ASAP7_75t_L g1054 ( .A(n_39), .B(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1305 ( .A(n_39), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_40), .Y(n_1174) );
AOI22xp33_ASAP7_75t_SL g1170 ( .A1(n_41), .A2(n_44), .B1(n_523), .B2(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1179 ( .A(n_41), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_42), .A2(n_260), .B1(n_508), .B2(n_509), .Y(n_868) );
AOI22xp33_ASAP7_75t_SL g880 ( .A1(n_42), .A2(n_260), .B1(n_881), .B2(n_882), .Y(n_880) );
INVx1_ASAP7_75t_L g593 ( .A(n_43), .Y(n_593) );
OAI211xp5_ASAP7_75t_SL g622 ( .A1(n_43), .A2(n_428), .B(n_623), .C(n_634), .Y(n_622) );
INVx1_ASAP7_75t_L g1178 ( .A(n_44), .Y(n_1178) );
INVx1_ASAP7_75t_L g1487 ( .A(n_45), .Y(n_1487) );
OAI22xp33_ASAP7_75t_L g1497 ( .A1(n_45), .A2(n_78), .B1(n_467), .B2(n_469), .Y(n_1497) );
INVx1_ASAP7_75t_L g806 ( .A(n_46), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_46), .A2(n_142), .B1(n_870), .B2(n_873), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_47), .A2(n_228), .B1(n_822), .B2(n_901), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g941 ( .A1(n_47), .A2(n_228), .B1(n_846), .B2(n_942), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_48), .A2(n_73), .B1(n_489), .B2(n_505), .C(n_633), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_48), .A2(n_73), .B1(n_778), .B2(n_779), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_49), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_50), .A2(n_263), .B1(n_489), .B2(n_490), .C(n_633), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_50), .A2(n_53), .B1(n_467), .B2(n_469), .Y(n_641) );
INVx1_ASAP7_75t_L g371 ( .A(n_51), .Y(n_371) );
INVx1_ASAP7_75t_L g1465 ( .A(n_52), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_52), .A2(n_65), .B1(n_388), .B2(n_396), .Y(n_1470) );
INVx1_ASAP7_75t_L g627 ( .A(n_53), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_56), .A2(n_253), .B1(n_321), .B2(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_56), .A2(n_253), .B1(n_670), .B2(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g685 ( .A(n_57), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g1031 ( .A1(n_58), .A2(n_68), .B1(n_923), .B2(n_1032), .C(n_1033), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_59), .A2(n_141), .B1(n_890), .B2(n_891), .Y(n_1012) );
INVx1_ASAP7_75t_L g1045 ( .A(n_59), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_60), .A2(n_225), .B1(n_964), .B2(n_966), .Y(n_963) );
INVx1_ASAP7_75t_L g818 ( .A(n_61), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_61), .A2(n_125), .B1(n_504), .B2(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g631 ( .A(n_62), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_62), .A2(n_263), .B1(n_464), .B2(n_528), .Y(n_640) );
INVx1_ASAP7_75t_L g1209 ( .A(n_63), .Y(n_1209) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_64), .Y(n_475) );
INVx1_ASAP7_75t_L g1464 ( .A(n_65), .Y(n_1464) );
AO221x1_ASAP7_75t_L g1186 ( .A1(n_66), .A2(n_93), .B1(n_440), .B2(n_442), .C(n_838), .Y(n_1186) );
INVx1_ASAP7_75t_L g1197 ( .A(n_66), .Y(n_1197) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_67), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_68), .A2(n_198), .B1(n_460), .B2(n_464), .Y(n_1052) );
INVx1_ASAP7_75t_L g1120 ( .A(n_69), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_69), .A2(n_135), .B1(n_937), .B2(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1087 ( .A(n_70), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_71), .A2(n_239), .B1(n_518), .B2(n_988), .Y(n_1064) );
OAI211xp5_ASAP7_75t_SL g1076 ( .A1(n_71), .A2(n_428), .B(n_1077), .C(n_1083), .Y(n_1076) );
INVx1_ASAP7_75t_L g353 ( .A(n_72), .Y(n_353) );
INVx1_ASAP7_75t_L g1122 ( .A(n_74), .Y(n_1122) );
AOI22xp33_ASAP7_75t_SL g1150 ( .A1(n_74), .A2(n_203), .B1(n_913), .B2(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g596 ( .A(n_75), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_76), .A2(n_128), .B1(n_453), .B2(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g541 ( .A(n_76), .Y(n_541) );
INVx1_ASAP7_75t_L g1277 ( .A(n_77), .Y(n_1277) );
INVx1_ASAP7_75t_L g1484 ( .A(n_78), .Y(n_1484) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_79), .A2(n_129), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g982 ( .A1(n_79), .A2(n_129), .B1(n_480), .B2(n_921), .Y(n_982) );
INVx1_ASAP7_75t_L g1116 ( .A(n_80), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_80), .A2(n_131), .B1(n_614), .B2(n_919), .Y(n_1138) );
XNOR2x2_ASAP7_75t_L g797 ( .A(n_81), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g958 ( .A(n_82), .Y(n_958) );
OAI222xp33_ASAP7_75t_L g970 ( .A1(n_82), .A2(n_164), .B1(n_181), .B2(n_971), .C1(n_972), .C2(n_973), .Y(n_970) );
INVx1_ASAP7_75t_L g1069 ( .A(n_83), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1082 ( .A1(n_83), .A2(n_174), .B1(n_484), .B2(n_838), .C(n_1033), .Y(n_1082) );
CKINVDCx16_ASAP7_75t_R g1228 ( .A(n_84), .Y(n_1228) );
INVx1_ASAP7_75t_L g436 ( .A(n_85), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_86), .A2(n_106), .B1(n_490), .B2(n_756), .C(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g785 ( .A(n_86), .Y(n_785) );
OAI222xp33_ASAP7_75t_L g1105 ( .A1(n_87), .A2(n_176), .B1(n_222), .B2(n_901), .C1(n_1106), .C2(n_1109), .Y(n_1105) );
INVx1_ASAP7_75t_L g1123 ( .A(n_87), .Y(n_1123) );
AO22x2_ASAP7_75t_L g1100 ( .A1(n_88), .A2(n_1101), .B1(n_1102), .B2(n_1156), .Y(n_1100) );
INVxp67_ASAP7_75t_SL g1101 ( .A(n_88), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_89), .A2(n_113), .B1(n_1136), .B2(n_1144), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_89), .A2(n_113), .B1(n_911), .B2(n_913), .Y(n_1146) );
INVx1_ASAP7_75t_L g307 ( .A(n_90), .Y(n_307) );
INVx1_ASAP7_75t_L g316 ( .A(n_90), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_91), .A2(n_153), .B1(n_913), .B2(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g948 ( .A(n_91), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g740 ( .A1(n_92), .A2(n_211), .B1(n_441), .B2(n_442), .C(n_486), .Y(n_740) );
INVx1_ASAP7_75t_L g1199 ( .A(n_93), .Y(n_1199) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_94), .Y(n_1192) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_95), .A2(n_97), .B1(n_365), .B2(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1035 ( .A(n_95), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_96), .A2(n_136), .B1(n_915), .B2(n_916), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_96), .A2(n_136), .B1(n_480), .B2(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1036 ( .A(n_97), .Y(n_1036) );
INVx1_ASAP7_75t_L g499 ( .A(n_98), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_98), .A2(n_99), .B1(n_561), .B2(n_563), .Y(n_560) );
INVx1_ASAP7_75t_L g500 ( .A(n_99), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_100), .A2(n_232), .B1(n_480), .B2(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g526 ( .A(n_100), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g1244 ( .A1(n_101), .A2(n_139), .B1(n_1233), .B2(n_1236), .Y(n_1244) );
INVx1_ASAP7_75t_L g710 ( .A(n_102), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_102), .A2(n_405), .B1(n_725), .B2(n_729), .C(n_734), .Y(n_724) );
AOI22x1_ASAP7_75t_L g1158 ( .A1(n_103), .A2(n_1159), .B1(n_1160), .B2(n_1200), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g1200 ( .A(n_103), .Y(n_1200) );
OAI22xp33_ASAP7_75t_L g1466 ( .A1(n_104), .A2(n_169), .B1(n_602), .B2(n_604), .Y(n_1466) );
INVx1_ASAP7_75t_L g1494 ( .A(n_104), .Y(n_1494) );
INVx1_ASAP7_75t_L g1112 ( .A(n_105), .Y(n_1112) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_105), .A2(n_222), .B1(n_930), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g787 ( .A(n_106), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_107), .Y(n_1060) );
INVx1_ASAP7_75t_L g1263 ( .A(n_109), .Y(n_1263) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_110), .Y(n_1059) );
INVx1_ASAP7_75t_L g762 ( .A(n_111), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_111), .A2(n_238), .B1(n_326), .B2(n_562), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_112), .A2(n_171), .B1(n_882), .B2(n_986), .Y(n_1062) );
INVx1_ASAP7_75t_L g1091 ( .A(n_112), .Y(n_1091) );
INVx1_ASAP7_75t_L g492 ( .A(n_114), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_114), .A2(n_248), .B1(n_552), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_115), .A2(n_219), .B1(n_753), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_115), .A2(n_219), .B1(n_562), .B2(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g897 ( .A(n_116), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_116), .A2(n_185), .B1(n_489), .B2(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g1015 ( .A(n_117), .Y(n_1015) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_117), .A2(n_405), .B1(n_734), .B2(n_1038), .C(n_1042), .Y(n_1037) );
AO221x2_ASAP7_75t_L g1274 ( .A1(n_118), .A2(n_179), .B1(n_1224), .B2(n_1230), .C(n_1275), .Y(n_1274) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_119), .Y(n_588) );
INVx1_ASAP7_75t_L g1459 ( .A(n_120), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_121), .A2(n_177), .B1(n_913), .B2(n_1167), .Y(n_1166) );
OAI221xp5_ASAP7_75t_L g1185 ( .A1(n_121), .A2(n_428), .B1(n_1186), .B2(n_1187), .C(n_1191), .Y(n_1185) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_122), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_123), .A2(n_213), .B1(n_936), .B2(n_937), .Y(n_1164) );
AOI22xp33_ASAP7_75t_SL g1181 ( .A1(n_123), .A2(n_213), .B1(n_414), .B2(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g592 ( .A(n_124), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_124), .A2(n_405), .B1(n_424), .B2(n_610), .C(n_618), .Y(n_609) );
INVx1_ASAP7_75t_L g801 ( .A(n_125), .Y(n_801) );
INVx1_ASAP7_75t_L g272 ( .A(n_126), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_127), .Y(n_904) );
INVx1_ASAP7_75t_L g542 ( .A(n_128), .Y(n_542) );
INVx1_ASAP7_75t_L g711 ( .A(n_130), .Y(n_711) );
OAI211xp5_ASAP7_75t_SL g735 ( .A1(n_130), .A2(n_428), .B(n_736), .C(n_741), .Y(n_735) );
INVx1_ASAP7_75t_L g1115 ( .A(n_131), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g1245 ( .A1(n_132), .A2(n_167), .B1(n_1230), .B2(n_1239), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_133), .A2(n_223), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g788 ( .A(n_133), .Y(n_788) );
INVx1_ASAP7_75t_L g839 ( .A(n_134), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_134), .A2(n_202), .B1(n_556), .B2(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g1119 ( .A(n_135), .Y(n_1119) );
INVx1_ASAP7_75t_L g1249 ( .A(n_137), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_138), .A2(n_216), .B1(n_453), .B2(n_494), .Y(n_760) );
INVx1_ASAP7_75t_L g791 ( .A(n_138), .Y(n_791) );
INVx1_ASAP7_75t_L g1468 ( .A(n_140), .Y(n_1468) );
INVx1_ASAP7_75t_L g1049 ( .A(n_141), .Y(n_1049) );
INVx1_ASAP7_75t_L g815 ( .A(n_142), .Y(n_815) );
INVx1_ASAP7_75t_L g792 ( .A(n_143), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_144), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_145), .A2(n_234), .B1(n_936), .B2(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g944 ( .A(n_145), .Y(n_944) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_146), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_147), .A2(n_221), .B1(n_602), .B2(n_604), .Y(n_716) );
INVx1_ASAP7_75t_L g743 ( .A(n_147), .Y(n_743) );
INVx1_ASAP7_75t_L g976 ( .A(n_148), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_148), .A2(n_151), .B1(n_890), .B2(n_891), .Y(n_993) );
INVx1_ASAP7_75t_L g714 ( .A(n_149), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_149), .A2(n_250), .B1(n_388), .B2(n_396), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_150), .A2(n_175), .B1(n_487), .B2(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_150), .A2(n_175), .B1(n_556), .B2(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g977 ( .A(n_151), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_152), .A2(n_157), .B1(n_1233), .B2(n_1236), .Y(n_1252) );
INVx1_ASAP7_75t_L g940 ( .A(n_153), .Y(n_940) );
AOI22x1_ASAP7_75t_SL g950 ( .A1(n_154), .A2(n_951), .B1(n_994), .B2(n_995), .Y(n_950) );
INVx1_ASAP7_75t_L g994 ( .A(n_154), .Y(n_994) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_155), .Y(n_324) );
INVx1_ASAP7_75t_L g1074 ( .A(n_156), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_158), .A2(n_207), .B1(n_1224), .B2(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g955 ( .A(n_159), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_159), .A2(n_225), .B1(n_836), .B2(n_867), .Y(n_983) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_160), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_160), .B(n_272), .Y(n_1212) );
AND3x2_ASAP7_75t_L g1227 ( .A(n_160), .B(n_272), .C(n_1215), .Y(n_1227) );
XNOR2xp5_ASAP7_75t_L g570 ( .A(n_161), .B(n_571), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_162), .Y(n_606) );
INVx1_ASAP7_75t_L g661 ( .A(n_163), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_163), .A2(n_405), .B1(n_424), .B2(n_673), .C(n_679), .Y(n_672) );
INVx1_ASAP7_75t_L g1462 ( .A(n_165), .Y(n_1462) );
OAI221xp5_ASAP7_75t_L g1479 ( .A1(n_165), .A2(n_428), .B1(n_1480), .B2(n_1486), .C(n_1492), .Y(n_1479) );
INVx2_ASAP7_75t_L g285 ( .A(n_166), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g1457 ( .A(n_168), .Y(n_1457) );
INVx1_ASAP7_75t_L g1493 ( .A(n_169), .Y(n_1493) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_170), .Y(n_329) );
INVx1_ASAP7_75t_L g1092 ( .A(n_171), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_172), .A2(n_196), .B1(n_508), .B2(n_509), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_172), .A2(n_196), .B1(n_548), .B2(n_550), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_173), .A2(n_211), .B1(n_464), .B2(n_528), .Y(n_718) );
INVx1_ASAP7_75t_L g739 ( .A(n_173), .Y(n_739) );
INVx1_ASAP7_75t_L g1071 ( .A(n_174), .Y(n_1071) );
INVx1_ASAP7_75t_L g1125 ( .A(n_176), .Y(n_1125) );
INVx1_ASAP7_75t_L g1184 ( .A(n_177), .Y(n_1184) );
AOI22xp5_ASAP7_75t_L g1238 ( .A1(n_178), .A2(n_184), .B1(n_1230), .B2(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g451 ( .A(n_180), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_181), .Y(n_957) );
INVx1_ASAP7_75t_L g820 ( .A(n_182), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_182), .A2(n_217), .B1(n_844), .B2(n_846), .Y(n_843) );
INVx1_ASAP7_75t_L g1215 ( .A(n_183), .Y(n_1215) );
XNOR2xp5_ASAP7_75t_L g1448 ( .A(n_184), .B(n_1449), .Y(n_1448) );
AOI22xp5_ASAP7_75t_L g1503 ( .A1(n_184), .A2(n_1504), .B1(n_1508), .B2(n_1512), .Y(n_1503) );
INVx1_ASAP7_75t_L g903 ( .A(n_185), .Y(n_903) );
CKINVDCx16_ASAP7_75t_R g1260 ( .A(n_186), .Y(n_1260) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_187), .A2(n_190), .B1(n_602), .B2(n_604), .Y(n_667) );
INVx1_ASAP7_75t_L g690 ( .A(n_187), .Y(n_690) );
INVx1_ASAP7_75t_L g1307 ( .A(n_188), .Y(n_1307) );
INVx1_ASAP7_75t_L g342 ( .A(n_189), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_189), .A2(n_405), .B1(n_408), .B2(n_415), .C(n_424), .Y(n_404) );
INVx1_ASAP7_75t_L g689 ( .A(n_190), .Y(n_689) );
INVx1_ASAP7_75t_L g906 ( .A(n_191), .Y(n_906) );
XNOR2xp5_ASAP7_75t_L g1000 ( .A(n_193), .B(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1021 ( .A(n_194), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_195), .A2(n_240), .B1(n_633), .B2(n_836), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_195), .A2(n_240), .B1(n_888), .B2(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g855 ( .A(n_197), .Y(n_855) );
INVx1_ASAP7_75t_L g1030 ( .A(n_198), .Y(n_1030) );
INVx1_ASAP7_75t_L g650 ( .A(n_199), .Y(n_650) );
INVx1_ASAP7_75t_L g287 ( .A(n_200), .Y(n_287) );
INVx2_ASAP7_75t_L g391 ( .A(n_200), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_201), .A2(n_230), .B1(n_881), .B2(n_1019), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_201), .A2(n_230), .B1(n_670), .B2(n_671), .Y(n_1050) );
INVx1_ASAP7_75t_L g858 ( .A(n_202), .Y(n_858) );
INVx1_ASAP7_75t_L g1130 ( .A(n_203), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_204), .Y(n_1010) );
INVx1_ASAP7_75t_L g1461 ( .A(n_205), .Y(n_1461) );
OAI221xp5_ASAP7_75t_L g1471 ( .A1(n_205), .A2(n_405), .B1(n_424), .B2(n_1472), .C(n_1476), .Y(n_1471) );
AOI22xp5_ASAP7_75t_L g1232 ( .A1(n_206), .A2(n_237), .B1(n_1233), .B2(n_1236), .Y(n_1232) );
INVx1_ASAP7_75t_L g529 ( .A(n_208), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_209), .A2(n_258), .B1(n_351), .B2(n_549), .Y(n_657) );
INVx1_ASAP7_75t_L g675 ( .A(n_209), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_210), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_212), .B(n_749), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_214), .Y(n_336) );
INVx1_ASAP7_75t_L g701 ( .A(n_215), .Y(n_701) );
INVx1_ASAP7_75t_L g790 ( .A(n_216), .Y(n_790) );
INVx1_ASAP7_75t_L g826 ( .A(n_217), .Y(n_826) );
INVx1_ASAP7_75t_L g1017 ( .A(n_220), .Y(n_1017) );
OAI211xp5_ASAP7_75t_SL g1023 ( .A1(n_220), .A2(n_428), .B(n_1024), .C(n_1034), .Y(n_1023) );
INVx1_ASAP7_75t_L g742 ( .A(n_221), .Y(n_742) );
INVx1_ASAP7_75t_L g784 ( .A(n_223), .Y(n_784) );
INVx1_ASAP7_75t_L g721 ( .A(n_224), .Y(n_721) );
INVx1_ASAP7_75t_L g654 ( .A(n_229), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_229), .A2(n_486), .B(n_505), .Y(n_681) );
INVx1_ASAP7_75t_L g1217 ( .A(n_231), .Y(n_1217) );
INVx1_ASAP7_75t_L g521 ( .A(n_232), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g1455 ( .A(n_233), .Y(n_1455) );
INVx1_ASAP7_75t_L g946 ( .A(n_234), .Y(n_946) );
INVx1_ASAP7_75t_L g703 ( .A(n_235), .Y(n_703) );
INVx1_ASAP7_75t_L g1216 ( .A(n_236), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_236), .B(n_1214), .Y(n_1221) );
INVx1_ASAP7_75t_L g763 ( .A(n_238), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_239), .A2(n_405), .B1(n_734), .B2(n_1085), .C(n_1090), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g601 ( .A1(n_241), .A2(n_243), .B1(n_602), .B2(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g636 ( .A(n_241), .Y(n_636) );
INVx1_ASAP7_75t_L g664 ( .A(n_242), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_242), .A2(n_428), .B(n_683), .C(n_688), .Y(n_682) );
INVx1_ASAP7_75t_L g637 ( .A(n_243), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_244), .Y(n_1011) );
INVx2_ASAP7_75t_L g284 ( .A(n_245), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_246), .B(n_532), .Y(n_531) );
XNOR2xp5_ASAP7_75t_L g647 ( .A(n_247), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g510 ( .A(n_248), .Y(n_510) );
INVx1_ASAP7_75t_L g1483 ( .A(n_249), .Y(n_1483) );
OAI22xp33_ASAP7_75t_L g1496 ( .A1(n_249), .A2(n_255), .B1(n_464), .B2(n_528), .Y(n_1496) );
INVx1_ASAP7_75t_L g715 ( .A(n_250), .Y(n_715) );
INVx1_ASAP7_75t_L g759 ( .A(n_251), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_251), .A2(n_262), .B1(n_518), .B2(n_537), .Y(n_781) );
INVx1_ASAP7_75t_L g1453 ( .A(n_252), .Y(n_1453) );
INVx1_ASAP7_75t_L g1488 ( .A(n_255), .Y(n_1488) );
BUFx3_ASAP7_75t_L g301 ( .A(n_256), .Y(n_301) );
INVx1_ASAP7_75t_L g328 ( .A(n_256), .Y(n_328) );
BUFx3_ASAP7_75t_L g302 ( .A(n_257), .Y(n_302) );
INVx1_ASAP7_75t_L g323 ( .A(n_257), .Y(n_323) );
INVx1_ASAP7_75t_L g678 ( .A(n_258), .Y(n_678) );
INVx1_ASAP7_75t_L g686 ( .A(n_259), .Y(n_686) );
XOR2xp5_ASAP7_75t_L g1505 ( .A(n_261), .B(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g765 ( .A(n_262), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_264), .Y(n_1068) );
INVx1_ASAP7_75t_L g345 ( .A(n_265), .Y(n_345) );
OAI211xp5_ASAP7_75t_L g427 ( .A1(n_265), .A2(n_428), .B(n_433), .C(n_446), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_288), .B(n_1201), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_275), .Y(n_269) );
AND2x4_ASAP7_75t_L g1502 ( .A(n_270), .B(n_276), .Y(n_1502) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_SL g1511 ( .A(n_271), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_271), .B(n_273), .Y(n_1517) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_273), .B(n_1511), .Y(n_1510) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x6_ASAP7_75t_L g861 ( .A(n_278), .B(n_356), .Y(n_861) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g423 ( .A(n_279), .B(n_287), .Y(n_423) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g505 ( .A(n_280), .B(n_506), .Y(n_505) );
INVx8_ASAP7_75t_L g857 ( .A(n_281), .Y(n_857) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
INVx1_ASAP7_75t_L g421 ( .A(n_282), .Y(n_421) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_282), .Y(n_619) );
BUFx2_ASAP7_75t_L g733 ( .A(n_282), .Y(n_733) );
OR2x6_ASAP7_75t_L g860 ( .A(n_282), .B(n_850), .Y(n_860) );
INVx2_ASAP7_75t_SL g1478 ( .A(n_282), .Y(n_1478) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g385 ( .A(n_284), .B(n_285), .Y(n_385) );
INVx2_ASAP7_75t_L g393 ( .A(n_284), .Y(n_393) );
AND2x4_ASAP7_75t_L g402 ( .A(n_284), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g419 ( .A(n_284), .Y(n_419) );
INVx1_ASAP7_75t_L g432 ( .A(n_284), .Y(n_432) );
INVx1_ASAP7_75t_L g395 ( .A(n_285), .Y(n_395) );
INVx2_ASAP7_75t_L g403 ( .A(n_285), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_285), .B(n_393), .Y(n_412) );
INVx1_ASAP7_75t_L g418 ( .A(n_285), .Y(n_418) );
INVx1_ASAP7_75t_L g450 ( .A(n_285), .Y(n_450) );
AND2x4_ASAP7_75t_L g845 ( .A(n_286), .B(n_450), .Y(n_845) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g846 ( .A(n_287), .B(n_847), .Y(n_846) );
OR2x2_ASAP7_75t_L g973 ( .A(n_287), .B(n_847), .Y(n_973) );
XOR2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_642), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_567), .B2(n_568), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
XNOR2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_472), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND4x1_ASAP7_75t_L g294 ( .A(n_295), .B(n_370), .C(n_386), .D(n_458), .Y(n_294) );
NOR3xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_312), .C(n_358), .Y(n_295) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_296), .Y(n_573) );
NOR3xp33_ASAP7_75t_SL g651 ( .A(n_296), .B(n_652), .C(n_667), .Y(n_651) );
NOR3xp33_ASAP7_75t_SL g697 ( .A(n_296), .B(n_698), .C(n_716), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_296), .A2(n_543), .B1(n_603), .B2(n_790), .C(n_791), .Y(n_789) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_296), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1172 ( .A1(n_296), .A2(n_543), .B1(n_603), .B2(n_1173), .C(n_1174), .Y(n_1172) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_303), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g780 ( .A(n_299), .Y(n_780) );
AND2x4_ASAP7_75t_L g829 ( .A(n_299), .B(n_830), .Y(n_829) );
BUFx6f_ASAP7_75t_L g899 ( .A(n_299), .Y(n_899) );
BUFx6f_ASAP7_75t_L g992 ( .A(n_299), .Y(n_992) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_300), .Y(n_538) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x4_ASAP7_75t_L g322 ( .A(n_301), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g369 ( .A(n_301), .Y(n_369) );
AND2x4_ASAP7_75t_L g327 ( .A(n_302), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_303), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_SL g364 ( .A(n_304), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_304), .B(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g604 ( .A(n_304), .B(n_366), .Y(n_604) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_305), .B(n_310), .Y(n_304) );
AND2x2_ASAP7_75t_L g374 ( .A(n_305), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g357 ( .A(n_308), .B(n_316), .Y(n_357) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g315 ( .A(n_309), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g804 ( .A(n_309), .Y(n_804) );
INVx1_ASAP7_75t_L g809 ( .A(n_309), .Y(n_809) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_309), .Y(n_814) );
OR2x6_ASAP7_75t_L g878 ( .A(n_310), .B(n_443), .Y(n_878) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g462 ( .A(n_311), .B(n_463), .Y(n_462) );
OAI33xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .A3(n_330), .B1(n_341), .B2(n_346), .B3(n_354), .Y(n_312) );
OAI33xp33_ASAP7_75t_L g574 ( .A1(n_313), .A2(n_575), .A3(n_583), .B1(n_589), .B2(n_594), .B3(n_600), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_313), .A2(n_653), .B1(n_658), .B2(n_660), .Y(n_652) );
OAI33xp33_ASAP7_75t_L g698 ( .A1(n_313), .A2(n_600), .A3(n_699), .B1(n_704), .B2(n_709), .B3(n_712), .Y(n_698) );
INVx1_ASAP7_75t_SL g1163 ( .A(n_313), .Y(n_1163) );
OAI33xp33_ASAP7_75t_L g1451 ( .A1(n_313), .A2(n_600), .A3(n_1452), .B1(n_1456), .B2(n_1460), .B3(n_1463), .Y(n_1451) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
OR2x6_ASAP7_75t_L g546 ( .A(n_314), .B(n_317), .Y(n_546) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g774 ( .A(n_315), .Y(n_774) );
INVx1_ASAP7_75t_L g833 ( .A(n_316), .Y(n_833) );
INVx2_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
BUFx2_ASAP7_75t_L g513 ( .A(n_317), .Y(n_513) );
OR2x2_ASAP7_75t_L g773 ( .A(n_317), .B(n_774), .Y(n_773) );
AND2x4_ASAP7_75t_L g865 ( .A(n_317), .B(n_423), .Y(n_865) );
AND2x4_ASAP7_75t_L g979 ( .A(n_317), .B(n_423), .Y(n_979) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g457 ( .A(n_318), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_324), .B1(n_325), .B2(n_329), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_320), .A2(n_576), .B1(n_577), .B2(n_582), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g1463 ( .A1(n_320), .A2(n_461), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_322), .Y(n_471) );
INVx2_ASAP7_75t_SL g524 ( .A(n_322), .Y(n_524) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_322), .Y(n_549) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_322), .Y(n_562) );
AND2x6_ASAP7_75t_L g807 ( .A(n_322), .B(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_L g1148 ( .A(n_322), .Y(n_1148) );
BUFx2_ASAP7_75t_L g1153 ( .A(n_322), .Y(n_1153) );
INVx1_ASAP7_75t_L g335 ( .A(n_323), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_324), .A2(n_329), .B1(n_409), .B2(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_326), .Y(n_550) );
INVx1_ASAP7_75t_L g702 ( .A(n_326), .Y(n_702) );
INVx1_ASAP7_75t_L g1454 ( .A(n_326), .Y(n_1454) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_327), .Y(n_352) );
INVx1_ASAP7_75t_L g461 ( .A(n_327), .Y(n_461) );
INVx1_ASAP7_75t_L g564 ( .A(n_327), .Y(n_564) );
INVx2_ASAP7_75t_L g581 ( .A(n_327), .Y(n_581) );
INVx1_ASAP7_75t_L g334 ( .A(n_328), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_336), .B1(n_337), .B2(n_340), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_331), .A2(n_342), .B1(n_343), .B2(n_345), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_331), .A2(n_705), .B1(n_706), .B2(n_708), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_331), .A2(n_655), .B1(n_710), .B2(n_711), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g1460 ( .A1(n_331), .A2(n_1458), .B1(n_1461), .B2(n_1462), .Y(n_1460) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g468 ( .A(n_332), .Y(n_468) );
INVx2_ASAP7_75t_L g1014 ( .A(n_332), .Y(n_1014) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g584 ( .A(n_333), .Y(n_584) );
INVx1_ASAP7_75t_L g591 ( .A(n_333), .Y(n_591) );
OR2x2_ASAP7_75t_L g964 ( .A(n_333), .B(n_965), .Y(n_964) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g339 ( .A(n_334), .B(n_335), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_336), .A2(n_340), .B1(n_416), .B2(n_420), .C(n_422), .Y(n_415) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx4f_ASAP7_75t_L g344 ( .A(n_339), .Y(n_344) );
INVx2_ASAP7_75t_L g465 ( .A(n_339), .Y(n_465) );
INVx1_ASAP7_75t_L g587 ( .A(n_339), .Y(n_587) );
INVx1_ASAP7_75t_L g663 ( .A(n_339), .Y(n_663) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_343), .Y(n_1016) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g655 ( .A(n_344), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B1(n_350), .B2(n_353), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_350), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_352), .Y(n_666) );
AND2x6_ASAP7_75t_L g816 ( .A(n_352), .B(n_803), .Y(n_816) );
INVx2_ASAP7_75t_L g883 ( .A(n_352), .Y(n_883) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_352), .Y(n_1171) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI33xp33_ASAP7_75t_L g771 ( .A1(n_355), .A2(n_772), .A3(n_775), .B1(n_777), .B2(n_781), .B3(n_782), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g931 ( .A(n_355), .B(n_932), .C(n_935), .Y(n_931) );
INVx1_ASAP7_75t_L g1155 ( .A(n_355), .Y(n_1155) );
AOI33xp33_ASAP7_75t_L g1162 ( .A1(n_355), .A2(n_1163), .A3(n_1164), .B1(n_1165), .B2(n_1166), .B3(n_1170), .Y(n_1162) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x4_ASAP7_75t_L g373 ( .A(n_356), .B(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g566 ( .A(n_356), .B(n_357), .Y(n_566) );
INVx2_ASAP7_75t_L g540 ( .A(n_359), .Y(n_540) );
INVx2_ASAP7_75t_L g603 ( .A(n_359), .Y(n_603) );
INVx1_ASAP7_75t_L g1006 ( .A(n_359), .Y(n_1006) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g825 ( .A(n_362), .Y(n_825) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g375 ( .A(n_363), .B(n_369), .Y(n_375) );
INVx2_ASAP7_75t_L g543 ( .A(n_365), .Y(n_543) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x6_ASAP7_75t_L g827 ( .A(n_368), .B(n_809), .Y(n_827) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g532 ( .A(n_372), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_372), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_372), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_372), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g749 ( .A(n_372), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_372), .B(n_1021), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_372), .B(n_1074), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_372), .B(n_1468), .Y(n_1467) );
OR2x6_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
AOI222xp33_ASAP7_75t_L g1196 ( .A1(n_373), .A2(n_517), .B1(n_527), .B2(n_1188), .C1(n_1192), .C2(n_1197), .Y(n_1196) );
INVx2_ASAP7_75t_L g519 ( .A(n_375), .Y(n_519) );
INVx6_ASAP7_75t_L g555 ( .A(n_375), .Y(n_555) );
BUFx2_ASAP7_75t_L g778 ( .A(n_375), .Y(n_778) );
AND2x4_ASAP7_75t_L g812 ( .A(n_375), .B(n_813), .Y(n_812) );
NOR2xp67_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx2_ASAP7_75t_L g638 ( .A(n_377), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_383), .Y(n_378) );
AND2x2_ASAP7_75t_L g448 ( .A(n_379), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g635 ( .A(n_379), .B(n_449), .Y(n_635) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x6_ASAP7_75t_L g424 ( .A(n_380), .B(n_425), .Y(n_424) );
OR2x6_ASAP7_75t_L g453 ( .A(n_380), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g497 ( .A(n_380), .Y(n_497) );
OR2x2_ASAP7_75t_L g734 ( .A(n_380), .B(n_425), .Y(n_734) );
INVx1_ASAP7_75t_L g1195 ( .A(n_380), .Y(n_1195) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g923 ( .A(n_383), .Y(n_923) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
INVx2_ASAP7_75t_SL g486 ( .A(n_384), .Y(n_486) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_385), .Y(n_407) );
OAI31xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_404), .A3(n_427), .B(n_455), .Y(n_386) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_389), .A2(n_397), .B1(n_499), .B2(n_500), .Y(n_498) );
INVx3_ASAP7_75t_L g670 ( .A(n_389), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_389), .A2(n_397), .B1(n_762), .B2(n_763), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_389), .A2(n_397), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx2_ASAP7_75t_L g399 ( .A(n_390), .Y(n_399) );
AND2x4_ASAP7_75t_L g406 ( .A(n_390), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g444 ( .A(n_391), .Y(n_444) );
INVx1_ASAP7_75t_L g506 ( .A(n_391), .Y(n_506) );
BUFx2_ASAP7_75t_L g480 ( .A(n_392), .Y(n_480) );
BUFx2_ASAP7_75t_L g508 ( .A(n_392), .Y(n_508) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_392), .Y(n_753) );
AND2x4_ASAP7_75t_L g849 ( .A(n_392), .B(n_850), .Y(n_849) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_392), .Y(n_872) );
INVx1_ASAP7_75t_L g920 ( .A(n_392), .Y(n_920) );
BUFx6f_ASAP7_75t_L g1182 ( .A(n_392), .Y(n_1182) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g454 ( .A(n_393), .Y(n_454) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g671 ( .A(n_397), .Y(n_671) );
AND2x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
AND2x4_ASAP7_75t_L g429 ( .A(n_398), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g928 ( .A(n_400), .Y(n_928) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g768 ( .A(n_401), .Y(n_768) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_402), .Y(n_414) );
INVx3_ASAP7_75t_L g617 ( .A(n_402), .Y(n_617) );
INVx1_ASAP7_75t_L g854 ( .A(n_402), .Y(n_854) );
AND2x4_ASAP7_75t_L g431 ( .A(n_403), .B(n_432), .Y(n_431) );
CKINVDCx6p67_ASAP7_75t_R g405 ( .A(n_406), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_406), .A2(n_502), .B1(n_507), .B2(n_510), .C(n_511), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_406), .A2(n_511), .B1(n_765), .B2(n_766), .C(n_767), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_406), .A2(n_1181), .B1(n_1183), .B2(n_1184), .Y(n_1180) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_407), .Y(n_633) );
BUFx2_ASAP7_75t_L g756 ( .A(n_407), .Y(n_756) );
INVx3_ASAP7_75t_L g1137 ( .A(n_407), .Y(n_1137) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g674 ( .A(n_410), .Y(n_674) );
INVx2_ASAP7_75t_L g684 ( .A(n_410), .Y(n_684) );
INVx2_ASAP7_75t_L g737 ( .A(n_410), .Y(n_737) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g1027 ( .A(n_411), .Y(n_1027) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g435 ( .A(n_412), .Y(n_435) );
BUFx2_ASAP7_75t_L g626 ( .A(n_412), .Y(n_626) );
INVx2_ASAP7_75t_SL g509 ( .A(n_413), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_413), .A2(n_684), .B1(n_685), .B2(n_686), .C(n_687), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_413), .A2(n_737), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_736) );
INVx4_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g437 ( .A(n_414), .Y(n_437) );
INVx2_ASAP7_75t_SL g482 ( .A(n_414), .Y(n_482) );
BUFx3_ASAP7_75t_L g873 ( .A(n_414), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_416), .A2(n_585), .B1(n_588), .B2(n_619), .C(n_620), .Y(n_618) );
BUFx3_ASAP7_75t_L g680 ( .A(n_416), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_416), .B(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1482 ( .A(n_416), .Y(n_1482) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x2_ASAP7_75t_L g426 ( .A(n_418), .B(n_419), .Y(n_426) );
INVx1_ASAP7_75t_L g847 ( .A(n_419), .Y(n_847) );
OAI221xp5_ASAP7_75t_L g1480 ( .A1(n_420), .A2(n_1481), .B1(n_1483), .B2(n_1484), .C(n_1485), .Y(n_1480) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g1088 ( .A(n_421), .Y(n_1088) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_422), .A2(n_1010), .B1(n_1011), .B2(n_1039), .C(n_1041), .Y(n_1038) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_422), .A2(n_1086), .B1(n_1087), .B2(n_1088), .C(n_1089), .Y(n_1085) );
BUFx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g621 ( .A(n_423), .Y(n_621) );
INVx2_ASAP7_75t_L g511 ( .A(n_424), .Y(n_511) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g730 ( .A(n_426), .Y(n_730) );
INVx2_ASAP7_75t_L g972 ( .A(n_426), .Y(n_972) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_426), .Y(n_1040) );
INVx8_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_429), .A2(n_479), .B1(n_483), .B2(n_492), .C(n_493), .Y(n_478) );
AOI221xp5_ASAP7_75t_SL g751 ( .A1(n_429), .A2(n_752), .B1(n_755), .B2(n_759), .C(n_760), .Y(n_751) );
INVx1_ASAP7_75t_L g758 ( .A(n_430), .Y(n_758) );
BUFx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g441 ( .A(n_431), .Y(n_441) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_431), .Y(n_489) );
BUFx6f_ASAP7_75t_L g838 ( .A(n_431), .Y(n_838) );
AND2x4_ASAP7_75t_L g840 ( .A(n_431), .B(n_841), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_437), .B2(n_438), .C(n_439), .Y(n_433) );
INVx1_ASAP7_75t_L g1044 ( .A(n_434), .Y(n_1044) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_435), .Y(n_612) );
INVx2_ASAP7_75t_L g1190 ( .A(n_435), .Y(n_1190) );
BUFx3_ASAP7_75t_L g867 ( .A(n_440), .Y(n_867) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g842 ( .A(n_444), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_451), .B2(n_452), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_448), .A2(n_452), .B1(n_742), .B2(n_743), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_448), .A2(n_452), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_448), .A2(n_452), .B1(n_1059), .B2(n_1060), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_448), .A2(n_452), .B1(n_1493), .B2(n_1494), .Y(n_1492) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_452), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_452), .A2(n_635), .B1(n_689), .B2(n_690), .Y(n_688) );
CKINVDCx11_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
OAI31xp33_ASAP7_75t_L g668 ( .A1(n_455), .A2(n_669), .A3(n_672), .B(n_682), .Y(n_668) );
OAI31xp33_ASAP7_75t_L g1075 ( .A1(n_455), .A2(n_1076), .A3(n_1084), .B(n_1094), .Y(n_1075) );
OAI21xp5_ASAP7_75t_L g1175 ( .A1(n_455), .A2(n_1176), .B(n_1185), .Y(n_1175) );
BUFx8_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g832 ( .A(n_457), .B(n_833), .Y(n_832) );
AND2x4_ASAP7_75t_L g967 ( .A(n_457), .B(n_833), .Y(n_967) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .Y(n_458) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
OR2x6_ASAP7_75t_L g528 ( .A(n_461), .B(n_462), .Y(n_528) );
INVx2_ASAP7_75t_L g776 ( .A(n_461), .Y(n_776) );
OR2x6_ASAP7_75t_L g464 ( .A(n_462), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g467 ( .A(n_462), .B(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g469 ( .A(n_462), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g520 ( .A(n_462), .Y(n_520) );
CKINVDCx6p67_ASAP7_75t_R g530 ( .A(n_464), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_465), .A2(n_590), .B1(n_592), .B2(n_593), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_465), .A2(n_1009), .B1(n_1010), .B2(n_1011), .C(n_1012), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1458 ( .A(n_465), .Y(n_1458) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g890 ( .A(n_471), .Y(n_890) );
BUFx4f_ASAP7_75t_L g915 ( .A(n_471), .Y(n_915) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
XNOR2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_475), .A2(n_1223), .B1(n_1228), .B2(n_1229), .Y(n_1222) );
NOR4xp75_ASAP7_75t_L g476 ( .A(n_477), .B(n_514), .C(n_531), .D(n_533), .Y(n_476) );
AOI31xp33_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_498), .A3(n_501), .B(n_512), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g503 ( .A(n_486), .Y(n_503) );
AOI211xp5_ASAP7_75t_L g939 ( .A1(n_487), .A2(n_840), .B(n_940), .C(n_941), .Y(n_939) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g504 ( .A(n_488), .Y(n_504) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g1485 ( .A(n_490), .Y(n_1485) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g1033 ( .A(n_491), .Y(n_1033) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_495), .A2(n_1127), .B1(n_1173), .B2(n_1174), .Y(n_1194) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g1121 ( .A1(n_504), .A2(n_1122), .B1(n_1123), .B2(n_1124), .C1(n_1125), .C2(n_1126), .Y(n_1121) );
INVx1_ASAP7_75t_L g850 ( .A(n_506), .Y(n_850) );
INVx2_ASAP7_75t_L g744 ( .A(n_512), .Y(n_744) );
CKINVDCx8_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
OAI31xp33_ASAP7_75t_L g1022 ( .A1(n_513), .A2(n_1023), .A3(n_1037), .B(n_1050), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_525), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B1(n_521), .B2(n_522), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_517), .A2(n_522), .B1(n_787), .B2(n_788), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_517), .A2(n_522), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g888 ( .A(n_519), .Y(n_888) );
AND2x2_ASAP7_75t_L g522 ( .A(n_520), .B(n_523), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g1198 ( .A1(n_522), .A2(n_530), .B1(n_1189), .B2(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g936 ( .A(n_524), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B1(n_529), .B2(n_530), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_527), .A2(n_530), .B1(n_784), .B2(n_785), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_527), .A2(n_530), .B1(n_1068), .B2(n_1069), .Y(n_1067) );
CKINVDCx6p67_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
NAND3xp33_ASAP7_75t_SL g533 ( .A(n_534), .B(n_539), .C(n_544), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND3xp33_ASAP7_75t_SL g1057 ( .A(n_536), .B(n_1058), .C(n_1061), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_537), .Y(n_559) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g557 ( .A(n_538), .Y(n_557) );
BUFx4f_ASAP7_75t_L g819 ( .A(n_538), .Y(n_819) );
BUFx3_ASAP7_75t_L g988 ( .A(n_538), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B1(n_542), .B2(n_543), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_543), .A2(n_1006), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
AOI33xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .A3(n_551), .B1(n_558), .B2(n_560), .B3(n_565), .Y(n_544) );
AOI33xp33_ASAP7_75t_L g879 ( .A1(n_545), .A2(n_565), .A3(n_880), .B1(n_884), .B2(n_887), .B3(n_889), .Y(n_879) );
AOI33xp33_ASAP7_75t_L g984 ( .A1(n_545), .A2(n_566), .A3(n_985), .B1(n_987), .B2(n_989), .B3(n_993), .Y(n_984) );
AOI33xp33_ASAP7_75t_L g1061 ( .A1(n_545), .A2(n_565), .A3(n_1062), .B1(n_1063), .B2(n_1064), .B3(n_1065), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_SL g1007 ( .A1(n_546), .A2(n_658), .B1(n_1008), .B2(n_1013), .Y(n_1007) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g595 ( .A(n_549), .Y(n_595) );
INVx1_ASAP7_75t_L g700 ( .A(n_549), .Y(n_700) );
BUFx3_ASAP7_75t_L g881 ( .A(n_549), .Y(n_881) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g805 ( .A(n_555), .Y(n_805) );
INVx2_ASAP7_75t_L g886 ( .A(n_555), .Y(n_886) );
INVx2_ASAP7_75t_L g912 ( .A(n_555), .Y(n_912) );
BUFx6f_ASAP7_75t_L g934 ( .A(n_555), .Y(n_934) );
INVx1_ASAP7_75t_L g1151 ( .A(n_555), .Y(n_1151) );
INVx2_ASAP7_75t_SL g1169 ( .A(n_555), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_556), .B(n_955), .Y(n_954) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_SL g713 ( .A(n_562), .Y(n_713) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g598 ( .A(n_564), .Y(n_598) );
INVx1_ASAP7_75t_L g891 ( .A(n_564), .Y(n_891) );
BUFx4f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx4_ASAP7_75t_L g600 ( .A(n_566), .Y(n_600) );
BUFx4f_ASAP7_75t_L g659 ( .A(n_566), .Y(n_659) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND4x1_ASAP7_75t_L g571 ( .A(n_572), .B(n_605), .C(n_607), .D(n_639), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .C(n_601), .Y(n_572) );
NOR3xp33_ASAP7_75t_SL g1450 ( .A(n_573), .B(n_1451), .C(n_1466), .Y(n_1450) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_576), .A2(n_582), .B1(n_611), .B2(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g916 ( .A(n_579), .Y(n_916) );
INVx1_ASAP7_75t_L g937 ( .A(n_579), .Y(n_937) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B1(n_586), .B2(n_588), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_584), .A2(n_654), .B1(n_655), .B2(n_656), .C(n_657), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_584), .A2(n_661), .B1(n_662), .B2(n_664), .C(n_665), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g1456 ( .A1(n_584), .A2(n_1457), .B1(n_1458), .B2(n_1459), .Y(n_1456) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g1110 ( .A(n_587), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_590), .Y(n_1009) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_599), .Y(n_594) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI31xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .A3(n_622), .B(n_638), .Y(n_607) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g728 ( .A(n_616), .Y(n_728) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_616), .Y(n_754) );
INVx2_ASAP7_75t_L g1491 ( .A(n_616), .Y(n_1491) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_617), .Y(n_630) );
INVx3_ASAP7_75t_L g1048 ( .A(n_617), .Y(n_1048) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_619), .Y(n_1041) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_620), .A2(n_705), .B1(n_708), .B2(n_730), .C(n_731), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g1476 ( .A1(n_620), .A2(n_730), .B1(n_1457), .B2(n_1459), .C(n_1477), .Y(n_1476) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B1(n_628), .B2(n_631), .C(n_632), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g677 ( .A(n_630), .Y(n_677) );
INVx1_ASAP7_75t_L g876 ( .A(n_633), .Y(n_876) );
INVx1_ASAP7_75t_L g769 ( .A(n_638), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_996), .Y(n_642) );
XNOR2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_794), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_746), .B2(n_793), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AO22x2_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_694), .B1(n_695), .B2(n_745), .Y(n_646) );
INVx1_ASAP7_75t_L g745 ( .A(n_647), .Y(n_745) );
AND4x1_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .C(n_668), .D(n_691), .Y(n_648) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_656), .A2(n_680), .B(n_681), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g707 ( .A(n_663), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_678), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_674), .A2(n_701), .B1(n_703), .B2(n_726), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g1472 ( .A1(n_674), .A2(n_1453), .B1(n_1455), .B2(n_1473), .Y(n_1472) );
OAI22xp5_ASAP7_75t_SL g1486 ( .A1(n_674), .A2(n_1487), .B1(n_1488), .B2(n_1489), .Y(n_1486) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND4x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_717), .C(n_720), .D(n_722), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g1452 ( .A1(n_700), .A2(n_1453), .B1(n_1454), .B2(n_1455), .Y(n_1452) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g986 ( .A(n_713), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
OAI31xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .A3(n_735), .B(n_744), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g921 ( .A(n_728), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_728), .A2(n_1188), .B1(n_1189), .B2(n_1190), .Y(n_1187) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_730), .Y(n_1086) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_737), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
OAI31xp33_ASAP7_75t_L g1469 ( .A1(n_744), .A2(n_1470), .A3(n_1471), .B(n_1479), .Y(n_1469) );
INVx2_ASAP7_75t_L g793 ( .A(n_746), .Y(n_793) );
XOR2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_792), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .C(n_770), .Y(n_747) );
AOI31xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_761), .A3(n_764), .B(n_769), .Y(n_750) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g1144 ( .A(n_758), .Y(n_1144) );
INVx1_ASAP7_75t_L g1081 ( .A(n_768), .Y(n_1081) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_783), .C(n_786), .D(n_789), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_772), .B(n_910), .C(n_914), .Y(n_909) );
NAND3xp33_ASAP7_75t_L g1145 ( .A(n_772), .B(n_1146), .C(n_1147), .Y(n_1145) );
INVx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx3_ASAP7_75t_L g913 ( .A(n_780), .Y(n_913) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
XNOR2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_892), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AOI211x1_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_831), .B(n_834), .C(n_862), .Y(n_798) );
NAND4xp25_ASAP7_75t_SL g799 ( .A(n_800), .B(n_810), .C(n_817), .D(n_828), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B1(n_806), .B2(n_807), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_802), .A2(n_812), .B1(n_903), .B2(n_904), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_802), .A2(n_812), .B1(n_1112), .B2(n_1113), .Y(n_1111) );
AND2x4_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
INVx1_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_804), .B(n_1108), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_807), .A2(n_816), .B1(n_906), .B2(n_907), .Y(n_905) );
CKINVDCx6p67_ASAP7_75t_R g961 ( .A(n_807), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_807), .A2(n_816), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
INVx1_ASAP7_75t_L g830 ( .A(n_808), .Y(n_830) );
INVx1_ASAP7_75t_L g965 ( .A(n_808), .Y(n_965) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B1(n_815), .B2(n_816), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_811), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
INVx4_ASAP7_75t_L g966 ( .A(n_812), .Y(n_966) );
AND2x4_ASAP7_75t_L g823 ( .A(n_813), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx4_ASAP7_75t_L g962 ( .A(n_816), .Y(n_962) );
AOI222xp33_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B1(n_820), .B2(n_821), .C1(n_826), .C2(n_827), .Y(n_817) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_823), .A2(n_827), .B1(n_957), .B2(n_958), .Y(n_956) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g1108 ( .A(n_825), .Y(n_1108) );
INVx3_ASAP7_75t_L g901 ( .A(n_827), .Y(n_901) );
INVx5_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AOI211xp5_ASAP7_75t_L g896 ( .A1(n_829), .A2(n_897), .B(n_898), .C(n_900), .Y(n_896) );
CKINVDCx8_ASAP7_75t_R g959 ( .A(n_829), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_829), .B(n_1105), .Y(n_1104) );
AOI221x1_ASAP7_75t_L g1102 ( .A1(n_831), .A2(n_1103), .B1(n_1117), .B2(n_1132), .C(n_1133), .Y(n_1102) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
AO211x2_ASAP7_75t_L g894 ( .A1(n_832), .A2(n_895), .B(n_908), .C(n_938), .Y(n_894) );
AOI31xp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_848), .A3(n_856), .B(n_861), .Y(n_834) );
AOI211xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_839), .B(n_840), .C(n_843), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx2_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_838), .Y(n_930) );
BUFx2_ASAP7_75t_L g1032 ( .A(n_838), .Y(n_1032) );
NOR3xp33_ASAP7_75t_L g969 ( .A(n_840), .B(n_970), .C(n_974), .Y(n_969) );
CKINVDCx11_ASAP7_75t_R g1131 ( .A(n_840), .Y(n_1131) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVxp67_ASAP7_75t_L g1128 ( .A(n_842), .Y(n_1128) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g942 ( .A(n_845), .Y(n_942) );
INVx2_ASAP7_75t_L g971 ( .A(n_845), .Y(n_971) );
INVx1_ASAP7_75t_L g1127 ( .A(n_847), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_851), .B1(n_852), .B2(n_855), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g943 ( .A1(n_849), .A2(n_944), .B1(n_945), .B2(n_946), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_849), .A2(n_945), .B1(n_976), .B2(n_977), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_849), .A2(n_852), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
AND2x4_ASAP7_75t_L g852 ( .A(n_850), .B(n_853), .Y(n_852) );
AND2x4_ASAP7_75t_L g945 ( .A(n_850), .B(n_853), .Y(n_945) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
HB1xp67_ASAP7_75t_L g1475 ( .A(n_854), .Y(n_1475) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_857), .A2(n_904), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_857), .A2(n_949), .B1(n_1113), .B2(n_1130), .Y(n_1129) );
INVx4_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx5_ASAP7_75t_L g949 ( .A(n_860), .Y(n_949) );
AOI31xp33_ASAP7_75t_L g938 ( .A1(n_861), .A2(n_939), .A3(n_943), .B(n_947), .Y(n_938) );
AO21x1_ASAP7_75t_SL g968 ( .A1(n_861), .A2(n_969), .B(n_975), .Y(n_968) );
CKINVDCx16_ASAP7_75t_R g1132 ( .A(n_861), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_879), .Y(n_862) );
AOI33xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_866), .A3(n_868), .B1(n_869), .B2(n_874), .B3(n_877), .Y(n_863) );
BUFx3_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_865), .B(n_926), .C(n_929), .Y(n_925) );
INVx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g1093 ( .A(n_873), .Y(n_1093) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AOI33xp33_ASAP7_75t_L g978 ( .A1(n_877), .A2(n_979), .A3(n_980), .B1(n_981), .B2(n_982), .B3(n_983), .Y(n_978) );
INVx6_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx5_ASAP7_75t_L g924 ( .A(n_878), .Y(n_924) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g1019 ( .A(n_883), .Y(n_1019) );
BUFx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_886), .Y(n_990) );
XNOR2x1_ASAP7_75t_L g892 ( .A(n_893), .B(n_950), .Y(n_892) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_902), .C(n_905), .Y(n_895) );
HB1xp67_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
NAND4xp25_ASAP7_75t_L g908 ( .A(n_909), .B(n_917), .C(n_925), .D(n_931), .Y(n_908) );
BUFx6f_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_922), .C(n_924), .Y(n_917) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g1134 ( .A(n_924), .B(n_1135), .C(n_1138), .Y(n_1134) );
INVx1_ASAP7_75t_L g1029 ( .A(n_927), .Y(n_1029) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g1124 ( .A(n_942), .Y(n_1124) );
AND4x1_ASAP7_75t_L g951 ( .A(n_952), .B(n_968), .C(n_978), .D(n_984), .Y(n_951) );
NAND4xp25_ASAP7_75t_L g995 ( .A(n_952), .B(n_968), .C(n_978), .D(n_984), .Y(n_995) );
OAI31xp33_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_960), .A3(n_963), .B(n_967), .Y(n_952) );
NAND3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_956), .C(n_959), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g1139 ( .A(n_979), .B(n_1140), .C(n_1143), .Y(n_1139) );
BUFx6f_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
AO22x2_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_999), .B1(n_1097), .B2(n_1098), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
AO22x1_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1054), .B1(n_1095), .B2(n_1096), .Y(n_999) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1000), .Y(n_1096) );
AND4x1_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1020), .C(n_1022), .D(n_1051), .Y(n_1001) );
NOR3xp33_ASAP7_75t_SL g1002 ( .A(n_1003), .B(n_1004), .C(n_1007), .Y(n_1002) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
OAI221xp5_ASAP7_75t_L g1013 ( .A1(n_1014), .A2(n_1015), .B1(n_1016), .B2(n_1017), .C(n_1018), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1024 ( .A1(n_1025), .A2(n_1028), .B1(n_1029), .B2(n_1030), .C(n_1031), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1078 ( .A(n_1027), .Y(n_1078) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_1043), .A2(n_1045), .B1(n_1046), .B2(n_1049), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_1047), .Y(n_1046) );
BUFx3_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1048), .Y(n_1142) );
NOR2xp33_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1053), .Y(n_1051) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1054), .Y(n_1095) );
AND3x1_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1073), .C(n_1075), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1066), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1070), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1077 ( .A1(n_1068), .A2(n_1072), .B1(n_1078), .B2(n_1079), .C(n_1082), .Y(n_1077) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
OAI22x1_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1100), .B1(n_1157), .B2(n_1158), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1102), .Y(n_1156) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1111), .C(n_1114), .Y(n_1103) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
NAND4xp25_ASAP7_75t_SL g1117 ( .A(n_1118), .B(n_1121), .C(n_1129), .D(n_1131), .Y(n_1117) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1128), .Y(n_1126) );
NAND4xp25_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1139), .C(n_1145), .D(n_1149), .Y(n_1133) );
A2O1A1Ixp33_ASAP7_75t_L g1191 ( .A1(n_1136), .A2(n_1192), .B(n_1193), .C(n_1195), .Y(n_1191) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
NAND3xp33_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1152), .C(n_1154), .Y(n_1149) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_SL g1157 ( .A(n_1158), .Y(n_1157) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
NAND4xp75_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1175), .C(n_1196), .D(n_1198), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1172), .Y(n_1161) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1180), .Y(n_1176) );
OAI221xp5_ASAP7_75t_SL g1201 ( .A1(n_1202), .A2(n_1442), .B1(n_1444), .B2(n_1498), .C(n_1503), .Y(n_1201) );
AND5x1_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1352), .C(n_1390), .D(n_1402), .E(n_1425), .Y(n_1202) );
A2O1A1Ixp33_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1206), .B(n_1294), .C(n_1328), .Y(n_1203) );
OAI211xp5_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1240), .B(n_1281), .C(n_1283), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1231), .Y(n_1205) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1206), .Y(n_1292) );
INVx3_ASAP7_75t_L g1314 ( .A(n_1206), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1206), .B(n_1273), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1206), .B(n_1327), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1206), .B(n_1338), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1206), .B(n_1231), .Y(n_1384) );
INVx3_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1207), .B(n_1231), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1316 ( .A(n_1207), .B(n_1317), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1222), .Y(n_1207) );
OAI22xp33_ASAP7_75t_L g1208 ( .A1(n_1209), .A2(n_1210), .B1(n_1217), .B2(n_1218), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1262 ( .A1(n_1210), .A2(n_1220), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1275 ( .A1(n_1210), .A2(n_1220), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
BUFx3_ASAP7_75t_L g1310 ( .A(n_1210), .Y(n_1310) );
BUFx6f_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_1211), .A2(n_1220), .B1(n_1248), .B2(n_1249), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1213), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1212), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1212), .Y(n_1235) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1213), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1216), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1515 ( .A(n_1214), .Y(n_1515) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1216), .Y(n_1226) );
HB1xp67_ASAP7_75t_L g1312 ( .A(n_1218), .Y(n_1312) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1221), .Y(n_1237) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1224), .Y(n_1306) );
BUFx3_ASAP7_75t_L g1443 ( .A(n_1224), .Y(n_1443) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1227), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1225), .B(n_1227), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1516 ( .A(n_1225), .Y(n_1516) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
AND2x4_ASAP7_75t_L g1230 ( .A(n_1226), .B(n_1227), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_1229), .A2(n_1259), .B1(n_1260), .B2(n_1261), .Y(n_1258) );
INVx1_ASAP7_75t_SL g1229 ( .A(n_1230), .Y(n_1229) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1230), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1231), .B(n_1273), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1231), .B(n_1273), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1231), .B(n_1274), .Y(n_1317) );
INVx2_ASAP7_75t_L g1327 ( .A(n_1231), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1231), .B(n_1274), .Y(n_1338) );
OAI211xp5_ASAP7_75t_L g1366 ( .A1(n_1231), .A2(n_1367), .B(n_1369), .C(n_1372), .Y(n_1366) );
OAI221xp5_ASAP7_75t_L g1392 ( .A1(n_1231), .A2(n_1281), .B1(n_1393), .B2(n_1395), .C(n_1396), .Y(n_1392) );
OAI211xp5_ASAP7_75t_L g1404 ( .A1(n_1231), .A2(n_1405), .B(n_1407), .C(n_1413), .Y(n_1404) );
AND2x4_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1238), .Y(n_1231) );
AND2x4_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1235), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1236 ( .A(n_1235), .B(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1239), .Y(n_1259) );
AOI211xp5_ASAP7_75t_L g1240 ( .A1(n_1241), .A2(n_1250), .B(n_1265), .C(n_1268), .Y(n_1240) );
AOI21xp33_ASAP7_75t_L g1346 ( .A1(n_1241), .A2(n_1347), .B(n_1349), .Y(n_1346) );
AOI21xp5_ASAP7_75t_L g1400 ( .A1(n_1241), .A2(n_1349), .B(n_1386), .Y(n_1400) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1242), .B(n_1266), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1242), .B(n_1256), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1242), .B(n_1250), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1242), .B(n_1251), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1246), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1243), .B(n_1246), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1243), .B(n_1280), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1243), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1243), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1243), .B(n_1257), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1245), .Y(n_1243) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1246), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1246), .B(n_1322), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1246), .B(n_1256), .Y(n_1337) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1246), .B(n_1256), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1246), .B(n_1250), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1250), .B(n_1321), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1250), .B(n_1359), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1256), .Y(n_1250) );
INVx4_ASAP7_75t_L g1266 ( .A(n_1251), .Y(n_1266) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1251), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1251), .B(n_1282), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_1251), .B(n_1267), .Y(n_1335) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1251), .B(n_1271), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1251), .B(n_1406), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1416 ( .A(n_1251), .B(n_1256), .Y(n_1416) );
AND2x6_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1253), .Y(n_1251) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
OAI22xp5_ASAP7_75t_L g1304 ( .A1(n_1255), .A2(n_1305), .B1(n_1306), .B2(n_1307), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1256), .B(n_1280), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1256), .B(n_1280), .Y(n_1319) );
NOR2xp33_ASAP7_75t_L g1363 ( .A(n_1256), .B(n_1364), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1256), .B(n_1321), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1256), .B(n_1298), .Y(n_1394) );
CKINVDCx6p67_ASAP7_75t_R g1256 ( .A(n_1257), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1257), .B(n_1267), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1257), .B(n_1298), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1345 ( .A(n_1257), .B(n_1322), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1257), .B(n_1321), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1257), .B(n_1359), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1257), .B(n_1279), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1257), .B(n_1322), .Y(n_1424) );
OR2x6_ASAP7_75t_SL g1257 ( .A(n_1258), .B(n_1262), .Y(n_1257) );
NOR2xp33_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1267), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1266), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1266), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1266), .B(n_1374), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1266), .B(n_1424), .Y(n_1430) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1267), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1278), .Y(n_1268) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1269), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1271), .Y(n_1269) );
INVx2_ASAP7_75t_L g1285 ( .A(n_1270), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1270), .B(n_1337), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1270), .B(n_1344), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1270), .B(n_1368), .Y(n_1367) );
OAI21xp33_ASAP7_75t_L g1385 ( .A1(n_1270), .A2(n_1347), .B(n_1386), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1270), .B(n_1399), .Y(n_1398) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_1270), .B(n_1327), .Y(n_1410) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1272), .Y(n_1291) );
O2A1O1Ixp33_ASAP7_75t_L g1341 ( .A1(n_1272), .A2(n_1342), .B(n_1343), .C(n_1346), .Y(n_1341) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1272), .B(n_1423), .Y(n_1422) );
INVx2_ASAP7_75t_SL g1272 ( .A(n_1273), .Y(n_1272) );
INVx2_ASAP7_75t_SL g1273 ( .A(n_1274), .Y(n_1273) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_1274), .Y(n_1357) );
NOR2xp33_ASAP7_75t_L g1380 ( .A(n_1278), .B(n_1381), .Y(n_1380) );
NOR3xp33_ASAP7_75t_L g1388 ( .A(n_1278), .B(n_1314), .C(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
OAI222xp33_ASAP7_75t_L g1315 ( .A1(n_1282), .A2(n_1316), .B1(n_1318), .B2(n_1320), .C1(n_1323), .C2(n_1325), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1401 ( .A(n_1282), .B(n_1316), .Y(n_1401) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_1284), .A2(n_1287), .B1(n_1290), .B2(n_1293), .Y(n_1283) );
NOR2x1_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1285), .B(n_1424), .Y(n_1423) );
NOR2x1_ASAP7_75t_R g1436 ( .A(n_1285), .B(n_1437), .Y(n_1436) );
OR2x2_ASAP7_75t_L g1441 ( .A(n_1285), .B(n_1300), .Y(n_1441) );
AOI221xp5_ASAP7_75t_L g1333 ( .A1(n_1289), .A2(n_1334), .B1(n_1336), .B2(n_1338), .C(n_1339), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1289), .B(n_1340), .Y(n_1339) );
A2O1A1Ixp33_ASAP7_75t_L g1396 ( .A1(n_1289), .A2(n_1303), .B(n_1397), .C(n_1400), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1292), .Y(n_1290) );
O2A1O1Ixp33_ASAP7_75t_SL g1352 ( .A1(n_1292), .A2(n_1353), .B(n_1366), .C(n_1375), .Y(n_1352) );
INVxp67_ASAP7_75t_SL g1294 ( .A(n_1295), .Y(n_1294) );
OAI211xp5_ASAP7_75t_L g1328 ( .A1(n_1295), .A2(n_1329), .B(n_1333), .C(n_1341), .Y(n_1328) );
AOI21xp5_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1313), .B(n_1315), .Y(n_1295) );
OAI21xp5_ASAP7_75t_SL g1296 ( .A1(n_1297), .A2(n_1299), .B(n_1301), .Y(n_1296) );
OAI21xp5_ASAP7_75t_SL g1360 ( .A1(n_1299), .A2(n_1361), .B(n_1365), .Y(n_1360) );
OAI21xp33_ASAP7_75t_SL g1376 ( .A1(n_1299), .A2(n_1377), .B(n_1378), .Y(n_1376) );
INVx2_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
NOR2xp33_ASAP7_75t_L g1411 ( .A(n_1300), .B(n_1412), .Y(n_1411) );
CKINVDCx14_ASAP7_75t_R g1301 ( .A(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1303), .B(n_1314), .Y(n_1313) );
CKINVDCx5p33_ASAP7_75t_R g1331 ( .A(n_1303), .Y(n_1331) );
AOI31xp33_ASAP7_75t_L g1375 ( .A1(n_1303), .A2(n_1376), .A3(n_1379), .B(n_1383), .Y(n_1375) );
OR2x6_ASAP7_75t_SL g1303 ( .A(n_1304), .B(n_1308), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1310), .B1(n_1311), .B2(n_1312), .Y(n_1308) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1313), .Y(n_1403) );
INVx1_ASAP7_75t_SL g1332 ( .A(n_1314), .Y(n_1332) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1316), .Y(n_1391) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1317), .Y(n_1374) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1319), .B(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1320), .Y(n_1340) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1321), .Y(n_1437) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_1324), .A2(n_1343), .B1(n_1384), .B2(n_1385), .C(n_1388), .Y(n_1383) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
AOI21xp5_ASAP7_75t_L g1379 ( .A1(n_1326), .A2(n_1342), .B(n_1380), .Y(n_1379) );
NOR2xp33_ASAP7_75t_L g1395 ( .A(n_1326), .B(n_1357), .Y(n_1395) );
A2O1A1Ixp33_ASAP7_75t_L g1353 ( .A1(n_1327), .A2(n_1354), .B(n_1355), .C(n_1360), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1327), .B(n_1331), .Y(n_1421) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1332), .Y(n_1330) );
OAI21xp33_ASAP7_75t_L g1428 ( .A1(n_1331), .A2(n_1357), .B(n_1429), .Y(n_1428) );
AOI21xp5_ASAP7_75t_L g1435 ( .A1(n_1331), .A2(n_1374), .B(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1336), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1338), .B(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1338), .Y(n_1434) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1343), .Y(n_1433) );
NOR2xp33_ASAP7_75t_L g1409 ( .A(n_1344), .B(n_1368), .Y(n_1409) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1354), .B(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1355), .Y(n_1426) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1358), .Y(n_1355) );
OAI21xp33_ASAP7_75t_L g1413 ( .A1(n_1356), .A2(n_1414), .B(n_1417), .Y(n_1413) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1357), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1359), .B(n_1416), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1359), .B(n_1440), .Y(n_1439) );
AOI211xp5_ASAP7_75t_L g1390 ( .A1(n_1361), .A2(n_1391), .B(n_1392), .C(n_1401), .Y(n_1390) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1367), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1368), .B(n_1371), .Y(n_1370) );
INVxp67_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
AOI22xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1404), .B1(n_1420), .B2(n_1422), .Y(n_1402) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1405), .Y(n_1427) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1406), .Y(n_1412) );
AOI21xp5_ASAP7_75t_L g1407 ( .A1(n_1408), .A2(n_1410), .B(n_1411), .Y(n_1407) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
INVxp67_ASAP7_75t_SL g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
OAI321xp33_ASAP7_75t_L g1425 ( .A1(n_1421), .A2(n_1426), .A3(n_1427), .B1(n_1428), .B2(n_1431), .C(n_1438), .Y(n_1425) );
INVxp33_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
A2O1A1Ixp33_ASAP7_75t_L g1431 ( .A1(n_1432), .A2(n_1433), .B(n_1434), .C(n_1435), .Y(n_1431) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
CKINVDCx5p33_ASAP7_75t_R g1442 ( .A(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
HB1xp67_ASAP7_75t_L g1507 ( .A(n_1449), .Y(n_1507) );
AND4x1_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1467), .C(n_1469), .D(n_1495), .Y(n_1449) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx2_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx2_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
INVx2_ASAP7_75t_SL g1490 ( .A(n_1491), .Y(n_1490) );
NOR2xp33_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1497), .Y(n_1495) );
CKINVDCx14_ASAP7_75t_R g1498 ( .A(n_1499), .Y(n_1498) );
BUFx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
INVxp33_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
CKINVDCx5p33_ASAP7_75t_R g1509 ( .A(n_1510), .Y(n_1509) );
A2O1A1Ixp33_ASAP7_75t_L g1513 ( .A1(n_1511), .A2(n_1514), .B(n_1516), .C(n_1517), .Y(n_1513) );
HB1xp67_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
endmodule