module fake_netlist_6_2775_n_29 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_29);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_29;

wire n_16;
wire n_21;
wire n_10;
wire n_24;
wire n_18;
wire n_15;
wire n_27;
wire n_14;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_19;
wire n_25;

AND2x2_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_3),
.B(n_6),
.Y(n_12)
);

BUFx8_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx5p33_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_2),
.Y(n_19)
);

AO21x2_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_4),
.B(n_8),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_11),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

OAI211xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_19),
.B(n_15),
.C(n_16),
.Y(n_24)
);

BUFx8_ASAP7_75t_SL g25 ( 
.A(n_23),
.Y(n_25)
);

NOR3xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_14),
.C(n_18),
.Y(n_26)
);

NAND4xp25_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_16),
.C(n_13),
.D(n_14),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_7),
.B1(n_20),
.B2(n_15),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_20),
.B1(n_26),
.B2(n_28),
.Y(n_29)
);


endmodule