module fake_jpeg_23686_n_76 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_75;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_19),
.Y(n_29)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_3),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_9),
.B1(n_15),
.B2(n_13),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_20),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_37),
.B1(n_11),
.B2(n_14),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_9),
.B1(n_18),
.B2(n_19),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_34),
.B1(n_15),
.B2(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_19),
.B1(n_20),
.B2(n_16),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_49),
.C(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_20),
.B1(n_8),
.B2(n_14),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_22),
.C(n_11),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_35),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_37),
.C(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_30),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_57),
.B1(n_14),
.B2(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_44),
.Y(n_57)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_49),
.B(n_40),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_50),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_48),
.B(n_47),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_51),
.C(n_50),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_62),
.C(n_60),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_57),
.C(n_5),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_39),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C1(n_7),
.C2(n_1),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_60),
.C(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_67),
.B(n_69),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_6),
.B(n_7),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_72),
.C(n_7),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_0),
.Y(n_76)
);


endmodule