module fake_jpeg_201_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_5),
.B(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_61),
.Y(n_75)
);

NAND2x1_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_2),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_46),
.B1(n_49),
.B2(n_40),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_49),
.B1(n_52),
.B2(n_51),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_83),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_81),
.Y(n_104)
);

OR2x4_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_63),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_37),
.B(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_50),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_44),
.C(n_47),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_63),
.C(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_42),
.B1(n_54),
.B2(n_69),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_41),
.B1(n_35),
.B2(n_34),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_106),
.Y(n_124)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_101),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_24),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_3),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_71),
.B1(n_37),
.B2(n_48),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_16),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_87),
.B(n_71),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_11),
.B(n_12),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_87),
.C(n_41),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_115),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_116),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_123),
.C(n_14),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_26),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_4),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_120),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_129),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_6),
.B(n_8),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_130),
.B(n_131),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_9),
.B(n_10),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_115),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_15),
.B(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_119),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_134),
.C(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_127),
.B1(n_126),
.B2(n_122),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_146),
.B(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_139),
.A3(n_137),
.B1(n_123),
.B2(n_109),
.C1(n_113),
.C2(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_132),
.B1(n_110),
.B2(n_135),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);


endmodule