module fake_jpeg_17863_n_92 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_24),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_0),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_34),
.B1(n_40),
.B2(n_37),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_47),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_17),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_0),
.Y(n_52)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_60),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_35),
.B1(n_32),
.B2(n_3),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_4),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_75),
.B1(n_19),
.B2(n_20),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_18),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_81),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_64),
.C(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_86),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

OAI31xp33_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_67),
.A3(n_77),
.B(n_72),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_72),
.C(n_76),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_27),
.B(n_28),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_29),
.Y(n_92)
);


endmodule