module fake_jpeg_21158_n_203 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_12),
.B1(n_22),
.B2(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_17),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_17),
.B1(n_22),
.B2(n_16),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_13),
.B1(n_21),
.B2(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_28),
.B1(n_29),
.B2(n_24),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_24),
.B(n_16),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_14),
.C(n_26),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_48),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_30),
.B1(n_25),
.B2(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_26),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_33),
.B(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_30),
.B1(n_25),
.B2(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_58),
.B(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_24),
.B1(n_31),
.B2(n_20),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_31),
.B1(n_39),
.B2(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_16),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_65),
.B(n_71),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_74),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_43),
.B(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_31),
.B1(n_37),
.B2(n_39),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_73),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_39),
.B1(n_26),
.B2(n_20),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_20),
.B1(n_21),
.B2(n_13),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_59),
.B1(n_58),
.B2(n_56),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_12),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.C(n_23),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_12),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_86),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_60),
.B1(n_53),
.B2(n_21),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_66),
.B(n_23),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_65),
.B(n_72),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_88),
.B(n_23),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_53),
.B(n_36),
.C(n_60),
.D(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_13),
.B1(n_23),
.B2(n_36),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_96),
.B1(n_69),
.B2(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_36),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_76),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_68),
.C(n_67),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_92),
.C(n_96),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_110),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_76),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_76),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_96),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_80),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_113),
.B(n_4),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_11),
.B1(n_9),
.B2(n_8),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_11),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_116),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_9),
.B1(n_8),
.B2(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_81),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_8),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_85),
.B1(n_81),
.B2(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_122),
.C(n_138),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_91),
.C(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

OAI21x1_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_88),
.B(n_83),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_132),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_131),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_111),
.Y(n_146)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_85),
.A3(n_93),
.B1(n_4),
.B2(n_5),
.C1(n_0),
.C2(n_7),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_112),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_3),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_98),
.B1(n_105),
.B2(n_104),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_110),
.B1(n_109),
.B2(n_105),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_4),
.C(n_5),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_146),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_97),
.B1(n_102),
.B2(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_126),
.B1(n_137),
.B2(n_128),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_98),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_149),
.C(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_4),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_122),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_5),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_138),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_144),
.B1(n_152),
.B2(n_131),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_123),
.B(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_134),
.B1(n_147),
.B2(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_166),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_152),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_165),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_176),
.B1(n_161),
.B2(n_158),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_146),
.CI(n_153),
.CON(n_174),
.SN(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_136),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_183),
.B1(n_173),
.B2(n_174),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_179),
.B(n_181),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_163),
.B(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_159),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_185),
.A3(n_154),
.B1(n_174),
.B2(n_149),
.C(n_181),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_172),
.B1(n_171),
.B2(n_169),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_189),
.A2(n_191),
.B1(n_187),
.B2(n_188),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_6),
.B(n_178),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_5),
.C(n_6),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_6),
.B(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_6),
.B(n_7),
.Y(n_195)
);

NAND2x1_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_200),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_198),
.Y(n_203)
);


endmodule