module real_aes_7175_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_1), .A2(n_143), .B(n_148), .C(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_2), .A2(n_138), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g450 ( .A(n_3), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_4), .B(n_162), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_5), .A2(n_15), .B1(n_711), .B2(n_712), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_5), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_6), .A2(n_138), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g143 ( .A(n_7), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g172 ( .A(n_8), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_9), .B(n_44), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_10), .A2(n_250), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_11), .B(n_153), .Y(n_189) );
INVx1_ASAP7_75t_L g472 ( .A(n_12), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_13), .B(n_152), .Y(n_520) );
INVx1_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_15), .Y(n_711) );
INVx1_ASAP7_75t_L g532 ( .A(n_16), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_17), .A2(n_173), .B(n_198), .C(n_200), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_18), .B(n_162), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_19), .B(n_461), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_20), .A2(n_438), .B1(n_710), .B2(n_713), .C1(n_716), .C2(n_720), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_21), .A2(n_102), .B1(n_113), .B2(n_722), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_22), .B(n_138), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_23), .B(n_258), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_24), .A2(n_152), .B(n_154), .C(n_158), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_25), .B(n_162), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_26), .B(n_153), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_27), .A2(n_156), .B(n_200), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_28), .B(n_153), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_29), .Y(n_218) );
INVx1_ASAP7_75t_L g232 ( .A(n_30), .Y(n_232) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_31), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_32), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_33), .B(n_153), .Y(n_451) );
INVx1_ASAP7_75t_L g255 ( .A(n_34), .Y(n_255) );
INVx1_ASAP7_75t_L g485 ( .A(n_35), .Y(n_485) );
INVx2_ASAP7_75t_L g141 ( .A(n_36), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_37), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_38), .A2(n_152), .B(n_211), .C(n_213), .Y(n_210) );
INVxp67_ASAP7_75t_L g256 ( .A(n_39), .Y(n_256) );
CKINVDCx14_ASAP7_75t_R g209 ( .A(n_40), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_41), .A2(n_148), .B(n_231), .C(n_237), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_42), .A2(n_143), .B(n_148), .C(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_43), .A2(n_90), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_43), .Y(n_122) );
INVx1_ASAP7_75t_L g484 ( .A(n_45), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_46), .A2(n_170), .B(n_171), .C(n_174), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_47), .B(n_153), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_48), .B(n_435), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_49), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_50), .Y(n_252) );
INVx1_ASAP7_75t_L g146 ( .A(n_51), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_52), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_53), .B(n_138), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_54), .A2(n_148), .B1(n_158), .B2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_55), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_56), .Y(n_447) );
CKINVDCx14_ASAP7_75t_R g168 ( .A(n_57), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_58), .A2(n_170), .B(n_213), .C(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_59), .Y(n_513) );
INVx1_ASAP7_75t_L g469 ( .A(n_60), .Y(n_469) );
INVx1_ASAP7_75t_L g144 ( .A(n_61), .Y(n_144) );
INVx1_ASAP7_75t_L g135 ( .A(n_62), .Y(n_135) );
INVx1_ASAP7_75t_SL g212 ( .A(n_63), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_65), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g221 ( .A(n_66), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_SL g460 ( .A1(n_67), .A2(n_213), .B(n_461), .C(n_462), .Y(n_460) );
INVxp67_ASAP7_75t_L g463 ( .A(n_68), .Y(n_463) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_70), .A2(n_138), .B(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_71), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_72), .A2(n_138), .B(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_73), .Y(n_488) );
INVx1_ASAP7_75t_L g507 ( .A(n_74), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_75), .A2(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g196 ( .A(n_76), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_77), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_78), .A2(n_143), .B(n_148), .C(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_79), .A2(n_138), .B(n_145), .Y(n_137) );
INVx1_ASAP7_75t_L g199 ( .A(n_80), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_81), .B(n_233), .Y(n_501) );
INVx2_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
INVx1_ASAP7_75t_L g186 ( .A(n_83), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_84), .B(n_461), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_85), .A2(n_143), .B(n_148), .C(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g108 ( .A(n_86), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g708 ( .A(n_86), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_86), .B(n_110), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_87), .A2(n_148), .B(n_220), .C(n_223), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_88), .B(n_165), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_89), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_90), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_91), .A2(n_143), .B(n_148), .C(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_92), .Y(n_524) );
INVx1_ASAP7_75t_L g459 ( .A(n_93), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_94), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_95), .B(n_233), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_96), .B(n_131), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_97), .B(n_131), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_98), .B(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g155 ( .A(n_99), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_100), .A2(n_138), .B(n_458), .Y(n_457) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g722 ( .A(n_103), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g433 ( .A(n_108), .Y(n_433) );
INVx1_ASAP7_75t_SL g435 ( .A(n_108), .Y(n_435) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_109), .B(n_708), .Y(n_715) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g707 ( .A(n_110), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_436), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g721 ( .A(n_116), .Y(n_721) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_431), .B(n_434), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B1(n_429), .B2(n_430), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_120), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_123), .A2(n_707), .B1(n_717), .B2(n_718), .Y(n_716) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g430 ( .A(n_124), .Y(n_430) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_355), .Y(n_124) );
NOR4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_297), .C(n_327), .D(n_337), .Y(n_125) );
OAI211xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_202), .B(n_260), .C(n_287), .Y(n_126) );
OAI222xp33_ASAP7_75t_L g382 ( .A1(n_127), .A2(n_302), .B1(n_383), .B2(n_384), .C1(n_385), .C2(n_386), .Y(n_382) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_177), .Y(n_127) );
AOI33xp33_ASAP7_75t_L g308 ( .A1(n_128), .A2(n_295), .A3(n_296), .B1(n_309), .B2(n_314), .B3(n_316), .Y(n_308) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_128), .A2(n_366), .B(n_368), .C(n_370), .Y(n_365) );
OR2x2_ASAP7_75t_L g381 ( .A(n_128), .B(n_367), .Y(n_381) );
INVx1_ASAP7_75t_L g414 ( .A(n_128), .Y(n_414) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_164), .Y(n_128) );
INVx2_ASAP7_75t_L g291 ( .A(n_129), .Y(n_291) );
AND2x2_ASAP7_75t_L g307 ( .A(n_129), .B(n_193), .Y(n_307) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_129), .Y(n_342) );
AND2x2_ASAP7_75t_L g371 ( .A(n_129), .B(n_164), .Y(n_371) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_137), .B(n_161), .Y(n_129) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_130), .A2(n_194), .B(n_201), .Y(n_193) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_130), .A2(n_207), .B(n_215), .Y(n_206) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx4_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_131), .A2(n_457), .B(n_464), .Y(n_456) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g248 ( .A(n_132), .Y(n_248) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_133), .B(n_134), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx2_ASAP7_75t_L g250 ( .A(n_138), .Y(n_250) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_139), .B(n_143), .Y(n_183) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g236 ( .A(n_140), .Y(n_236) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
INVx1_ASAP7_75t_L g159 ( .A(n_141), .Y(n_159) );
INVx1_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
INVx3_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
INVx1_ASAP7_75t_L g461 ( .A(n_142), .Y(n_461) );
INVx4_ASAP7_75t_SL g160 ( .A(n_143), .Y(n_160) );
BUFx3_ASAP7_75t_L g237 ( .A(n_143), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_SL g145 ( .A1(n_146), .A2(n_147), .B(n_151), .C(n_160), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_SL g167 ( .A1(n_147), .A2(n_160), .B(n_168), .C(n_169), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_SL g195 ( .A1(n_147), .A2(n_160), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_147), .A2(n_160), .B(n_209), .C(n_210), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_SL g251 ( .A1(n_147), .A2(n_160), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_147), .A2(n_160), .B(n_459), .C(n_460), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_147), .A2(n_160), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_147), .A2(n_160), .B(n_529), .C(n_530), .Y(n_528) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx3_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_149), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_152), .B(n_212), .Y(n_211) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_156), .B(n_199), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g254 ( .A1(n_156), .A2(n_233), .B1(n_255), .B2(n_256), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_156), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_157), .A2(n_188), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g452 ( .A(n_158), .Y(n_452) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g223 ( .A(n_160), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_160), .A2(n_183), .B1(n_482), .B2(n_486), .Y(n_481) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_162), .A2(n_467), .B(n_473), .Y(n_466) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_163), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_163), .A2(n_217), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_163), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_SL g503 ( .A(n_163), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g271 ( .A(n_164), .Y(n_271) );
BUFx3_ASAP7_75t_L g279 ( .A(n_164), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_164), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g290 ( .A(n_164), .B(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_164), .B(n_178), .Y(n_319) );
AND2x2_ASAP7_75t_L g388 ( .A(n_164), .B(n_322), .Y(n_388) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_176), .Y(n_164) );
INVx1_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
INVx2_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_165), .A2(n_183), .B(n_229), .C(n_230), .Y(n_228) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_165), .A2(n_527), .B(n_533), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx5_ASAP7_75t_L g233 ( .A(n_173), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_173), .B(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_173), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g190 ( .A(n_174), .Y(n_190) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g200 ( .A(n_175), .Y(n_200) );
INVx2_ASAP7_75t_SL g282 ( .A(n_177), .Y(n_282) );
OR2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_178), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g324 ( .A(n_178), .Y(n_324) );
AND2x2_ASAP7_75t_L g335 ( .A(n_178), .B(n_291), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_178), .B(n_320), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_178), .B(n_322), .Y(n_367) );
AND2x2_ASAP7_75t_L g426 ( .A(n_178), .B(n_371), .Y(n_426) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g296 ( .A(n_179), .B(n_193), .Y(n_296) );
AND2x2_ASAP7_75t_L g306 ( .A(n_179), .B(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g328 ( .A(n_179), .Y(n_328) );
AND3x2_ASAP7_75t_L g387 ( .A(n_179), .B(n_388), .C(n_389), .Y(n_387) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_191), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_180), .B(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_180), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_180), .B(n_524), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_183), .A2(n_218), .B(n_219), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_183), .A2(n_447), .B(n_448), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_183), .A2(n_507), .B(n_508), .Y(n_506) );
O2A1O1Ixp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_189), .C(n_190), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_187), .A2(n_190), .B(n_221), .C(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_190), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_190), .A2(n_510), .B(n_511), .Y(n_509) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_193), .Y(n_278) );
INVx1_ASAP7_75t_SL g322 ( .A(n_193), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_193), .B(n_271), .C(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_240), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_203), .A2(n_306), .B(n_358), .C(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_205), .B(n_227), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_205), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g374 ( .A(n_205), .Y(n_374) );
AND2x2_ASAP7_75t_L g395 ( .A(n_205), .B(n_242), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_205), .B(n_304), .Y(n_423) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
AND2x2_ASAP7_75t_L g268 ( .A(n_206), .B(n_259), .Y(n_268) );
INVx2_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
AND2x2_ASAP7_75t_L g295 ( .A(n_206), .B(n_242), .Y(n_295) );
AND2x2_ASAP7_75t_L g345 ( .A(n_206), .B(n_227), .Y(n_345) );
INVx1_ASAP7_75t_L g349 ( .A(n_206), .Y(n_349) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_214), .Y(n_521) );
INVx2_ASAP7_75t_SL g259 ( .A(n_216), .Y(n_259) );
BUFx2_ASAP7_75t_L g285 ( .A(n_216), .Y(n_285) );
AND2x2_ASAP7_75t_L g412 ( .A(n_216), .B(n_227), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx1_ASAP7_75t_L g258 ( .A(n_226), .Y(n_258) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_226), .A2(n_516), .B(n_523), .Y(n_515) );
INVx3_ASAP7_75t_SL g242 ( .A(n_227), .Y(n_242) );
AND2x2_ASAP7_75t_L g267 ( .A(n_227), .B(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g274 ( .A(n_227), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g304 ( .A(n_227), .B(n_264), .Y(n_304) );
OR2x2_ASAP7_75t_L g313 ( .A(n_227), .B(n_259), .Y(n_313) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_227), .Y(n_331) );
AND2x2_ASAP7_75t_L g336 ( .A(n_227), .B(n_289), .Y(n_336) );
AND2x2_ASAP7_75t_L g364 ( .A(n_227), .B(n_244), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_227), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g402 ( .A(n_227), .B(n_243), .Y(n_402) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_238), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .C(n_235), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_233), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_236), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g326 ( .A(n_242), .B(n_275), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_242), .B(n_268), .Y(n_354) );
AND2x2_ASAP7_75t_L g372 ( .A(n_242), .B(n_289), .Y(n_372) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_259), .Y(n_243) );
AND2x2_ASAP7_75t_L g273 ( .A(n_244), .B(n_259), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_244), .B(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g311 ( .A(n_244), .Y(n_311) );
OR2x2_ASAP7_75t_L g359 ( .A(n_244), .B(n_279), .Y(n_359) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .B(n_257), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_246), .A2(n_265), .B(n_266), .Y(n_264) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_246), .A2(n_506), .B(n_512), .Y(n_505) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AOI21xp5_ASAP7_75t_SL g497 ( .A1(n_247), .A2(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_248), .A2(n_446), .B(n_453), .Y(n_445) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_248), .A2(n_481), .B(n_487), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_248), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g265 ( .A(n_249), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_257), .Y(n_266) );
AND2x2_ASAP7_75t_L g294 ( .A(n_259), .B(n_264), .Y(n_294) );
INVx1_ASAP7_75t_L g302 ( .A(n_259), .Y(n_302) );
AND2x2_ASAP7_75t_L g397 ( .A(n_259), .B(n_275), .Y(n_397) );
AOI222xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_269), .B1(n_272), .B2(n_276), .C1(n_280), .C2(n_283), .Y(n_260) );
INVx1_ASAP7_75t_L g392 ( .A(n_261), .Y(n_392) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
AND2x2_ASAP7_75t_L g288 ( .A(n_262), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g299 ( .A(n_262), .B(n_268), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_262), .B(n_290), .Y(n_315) );
OAI222xp33_ASAP7_75t_L g337 ( .A1(n_262), .A2(n_338), .B1(n_343), .B2(n_344), .C1(n_352), .C2(n_354), .Y(n_337) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g325 ( .A(n_264), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_264), .B(n_345), .Y(n_385) );
AND2x2_ASAP7_75t_L g396 ( .A(n_264), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g404 ( .A(n_267), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_269), .B(n_320), .Y(n_383) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_271), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g341 ( .A(n_271), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx3_ASAP7_75t_L g286 ( .A(n_274), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g376 ( .A1(n_274), .A2(n_377), .B(n_380), .C(n_382), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_274), .B(n_311), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_274), .B(n_294), .Y(n_416) );
AND2x2_ASAP7_75t_L g289 ( .A(n_275), .B(n_285), .Y(n_289) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g316 ( .A(n_278), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_279), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g368 ( .A(n_279), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g407 ( .A(n_279), .B(n_307), .Y(n_407) );
INVx1_ASAP7_75t_L g419 ( .A(n_279), .Y(n_419) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_282), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g400 ( .A(n_285), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_290), .B(n_292), .C(n_296), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_288), .A2(n_318), .B1(n_333), .B2(n_336), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_289), .B(n_303), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_289), .B(n_311), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_290), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g353 ( .A(n_290), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_290), .B(n_340), .Y(n_360) );
INVx2_ASAP7_75t_L g321 ( .A(n_291), .Y(n_321) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NOR4xp25_ASAP7_75t_L g298 ( .A(n_295), .B(n_299), .C(n_300), .D(n_303), .Y(n_298) );
INVx1_ASAP7_75t_SL g369 ( .A(n_296), .Y(n_369) );
AND2x2_ASAP7_75t_L g413 ( .A(n_296), .B(n_414), .Y(n_413) );
OAI211xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_305), .B(n_308), .C(n_317), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_304), .B(n_374), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_306), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_424) );
INVx1_ASAP7_75t_SL g379 ( .A(n_307), .Y(n_379) );
AND2x2_ASAP7_75t_L g418 ( .A(n_307), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_311), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_315), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_316), .B(n_341), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_323), .B(n_325), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g393 ( .A(n_320), .Y(n_393) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g421 ( .A(n_321), .Y(n_421) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B(n_332), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_328), .Y(n_340) );
OR2x2_ASAP7_75t_L g378 ( .A(n_328), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_331), .A2(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_335), .A2(n_362), .B1(n_365), .B2(n_372), .C(n_373), .Y(n_361) );
INVx1_ASAP7_75t_SL g405 ( .A(n_336), .Y(n_405) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
OR2x2_ASAP7_75t_L g352 ( .A(n_340), .B(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_349), .B2(n_350), .Y(n_344) );
INVx1_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_348), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR4xp25_ASAP7_75t_L g355 ( .A(n_356), .B(n_390), .C(n_403), .D(n_415), .Y(n_355) );
NAND3xp33_ASAP7_75t_SL g356 ( .A(n_357), .B(n_361), .C(n_376), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_359), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_366), .B(n_371), .Y(n_375) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_378), .A2(n_404), .B1(n_405), .B2(n_406), .C(n_408), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_380), .A2(n_395), .B(n_396), .C(n_398), .Y(n_394) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_381), .A2(n_399), .B1(n_401), .B2(n_402), .Y(n_398) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_393), .C(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g409 ( .A(n_402), .Y(n_409) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI21xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_410), .B(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_417), .B1(n_420), .B2(n_422), .C(n_424), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g438 ( .A1(n_430), .A2(n_439), .B1(n_707), .B2(n_709), .Y(n_438) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_434), .A2(n_437), .B(n_721), .Y(n_436) );
INVx1_ASAP7_75t_L g717 ( .A(n_439), .Y(n_717) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_623), .Y(n_439) );
NOR5xp2_ASAP7_75t_L g440 ( .A(n_441), .B(n_546), .C(n_578), .D(n_593), .E(n_610), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_474), .B(n_493), .C(n_534), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_455), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_443), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_443), .B(n_598), .Y(n_661) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_444), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_444), .B(n_490), .Y(n_547) );
AND2x2_ASAP7_75t_L g588 ( .A(n_444), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_444), .B(n_557), .Y(n_592) );
OR2x2_ASAP7_75t_L g629 ( .A(n_444), .B(n_480), .Y(n_629) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g479 ( .A(n_445), .B(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g537 ( .A(n_445), .Y(n_537) );
OR2x2_ASAP7_75t_L g700 ( .A(n_445), .B(n_540), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_455), .A2(n_603), .B1(n_604), .B2(n_607), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_455), .B(n_537), .Y(n_686) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
AND2x2_ASAP7_75t_L g492 ( .A(n_456), .B(n_480), .Y(n_492) );
AND2x2_ASAP7_75t_L g539 ( .A(n_456), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g544 ( .A(n_456), .Y(n_544) );
INVx3_ASAP7_75t_L g557 ( .A(n_456), .Y(n_557) );
OR2x2_ASAP7_75t_L g577 ( .A(n_456), .B(n_540), .Y(n_577) );
AND2x2_ASAP7_75t_L g596 ( .A(n_456), .B(n_466), .Y(n_596) );
BUFx2_ASAP7_75t_L g628 ( .A(n_456), .Y(n_628) );
AND2x4_ASAP7_75t_L g543 ( .A(n_465), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g478 ( .A(n_466), .Y(n_478) );
INVx2_ASAP7_75t_L g491 ( .A(n_466), .Y(n_491) );
OR2x2_ASAP7_75t_L g559 ( .A(n_466), .B(n_540), .Y(n_559) );
AND2x2_ASAP7_75t_L g589 ( .A(n_466), .B(n_480), .Y(n_589) );
AND2x2_ASAP7_75t_L g606 ( .A(n_466), .B(n_537), .Y(n_606) );
AND2x2_ASAP7_75t_L g646 ( .A(n_466), .B(n_557), .Y(n_646) );
AND2x2_ASAP7_75t_SL g682 ( .A(n_466), .B(n_492), .Y(n_682) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp33_ASAP7_75t_SL g475 ( .A(n_476), .B(n_489), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_477), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_478), .A2(n_492), .B(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_478), .B(n_480), .Y(n_676) );
AND2x2_ASAP7_75t_L g612 ( .A(n_479), .B(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g540 ( .A(n_480), .Y(n_540) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_480), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_489), .B(n_537), .Y(n_705) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_490), .A2(n_648), .B1(n_649), .B2(n_654), .Y(n_647) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x2_ASAP7_75t_L g538 ( .A(n_491), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g576 ( .A(n_491), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g613 ( .A(n_491), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_492), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g667 ( .A(n_492), .Y(n_667) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_514), .Y(n_494) );
INVx4_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
AND2x2_ASAP7_75t_L g631 ( .A(n_495), .B(n_598), .Y(n_631) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
INVx3_ASAP7_75t_L g550 ( .A(n_496), .Y(n_550) );
AND2x2_ASAP7_75t_L g564 ( .A(n_496), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g568 ( .A(n_496), .Y(n_568) );
INVx2_ASAP7_75t_L g582 ( .A(n_496), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_496), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g639 ( .A(n_496), .B(n_634), .Y(n_639) );
AND2x2_ASAP7_75t_L g704 ( .A(n_496), .B(n_674), .Y(n_704) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
AND2x2_ASAP7_75t_L g545 ( .A(n_505), .B(n_526), .Y(n_545) );
INVx2_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
INVx1_ASAP7_75t_L g570 ( .A(n_514), .Y(n_570) );
AND2x2_ASAP7_75t_L g616 ( .A(n_514), .B(n_564), .Y(n_616) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_525), .Y(n_514) );
INVx2_ASAP7_75t_L g555 ( .A(n_515), .Y(n_555) );
INVx1_ASAP7_75t_L g563 ( .A(n_515), .Y(n_563) );
AND2x2_ASAP7_75t_L g581 ( .A(n_515), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_515), .B(n_565), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_522), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_521), .Y(n_518) );
AND2x2_ASAP7_75t_L g598 ( .A(n_525), .B(n_555), .Y(n_598) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g551 ( .A(n_526), .Y(n_551) );
AND2x2_ASAP7_75t_L g634 ( .A(n_526), .B(n_565), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_541), .B(n_545), .Y(n_534) );
INVx1_ASAP7_75t_SL g579 ( .A(n_535), .Y(n_579) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_536), .B(n_543), .Y(n_636) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g585 ( .A(n_537), .B(n_540), .Y(n_585) );
AND2x2_ASAP7_75t_L g614 ( .A(n_537), .B(n_558), .Y(n_614) );
OR2x2_ASAP7_75t_L g617 ( .A(n_537), .B(n_577), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_538), .A2(n_630), .B1(n_682), .B2(n_683), .C1(n_685), .C2(n_687), .Y(n_681) );
BUFx2_ASAP7_75t_L g595 ( .A(n_540), .Y(n_595) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g584 ( .A(n_543), .B(n_585), .Y(n_584) );
INVx3_ASAP7_75t_SL g601 ( .A(n_543), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_543), .B(n_595), .Y(n_655) );
AND2x2_ASAP7_75t_L g590 ( .A(n_545), .B(n_550), .Y(n_590) );
INVx1_ASAP7_75t_L g609 ( .A(n_545), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_548), .B1(n_552), .B2(n_556), .C(n_560), .Y(n_546) );
OR2x2_ASAP7_75t_L g618 ( .A(n_548), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g603 ( .A(n_550), .B(n_573), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_550), .B(n_563), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_550), .B(n_598), .Y(n_648) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_550), .Y(n_658) );
NAND2x1_ASAP7_75t_SL g669 ( .A(n_550), .B(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g554 ( .A(n_551), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g574 ( .A(n_551), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_551), .B(n_569), .Y(n_600) );
INVx1_ASAP7_75t_L g666 ( .A(n_551), .Y(n_666) );
INVx1_ASAP7_75t_L g641 ( .A(n_552), .Y(n_641) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g653 ( .A(n_553), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g665 ( .A(n_553), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g670 ( .A(n_554), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_554), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g573 ( .A(n_555), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_555), .B(n_565), .Y(n_586) );
INVx1_ASAP7_75t_L g652 ( .A(n_555), .Y(n_652) );
INVx1_ASAP7_75t_L g673 ( .A(n_556), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI21xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_566), .B(n_575), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
AND2x2_ASAP7_75t_L g706 ( .A(n_562), .B(n_639), .Y(n_706) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g674 ( .A(n_563), .B(n_634), .Y(n_674) );
AOI32xp33_ASAP7_75t_L g587 ( .A1(n_564), .A2(n_570), .A3(n_588), .B1(n_590), .B2(n_591), .Y(n_587) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_564), .A2(n_596), .A3(n_679), .B1(n_690), .B2(n_691), .C1(n_692), .C2(n_694), .Y(n_689) );
INVx2_ASAP7_75t_L g569 ( .A(n_565), .Y(n_569) );
INVx1_ASAP7_75t_L g679 ( .A(n_565), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_570), .B1(n_571), .B2(n_572), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_567), .B(n_573), .Y(n_622) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_568), .B(n_634), .Y(n_684) );
INVx1_ASAP7_75t_L g571 ( .A(n_569), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_569), .B(n_598), .Y(n_688) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_577), .B(n_672), .Y(n_671) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_580), .B1(n_583), .B2(n_586), .C(n_587), .Y(n_578) );
OR2x2_ASAP7_75t_L g599 ( .A(n_580), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g608 ( .A(n_580), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g633 ( .A(n_581), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g637 ( .A(n_591), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B1(n_599), .B2(n_601), .C(n_602), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_595), .A2(n_626), .B1(n_630), .B2(n_631), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_596), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g701 ( .A(n_596), .Y(n_701) );
INVx1_ASAP7_75t_L g695 ( .A(n_598), .Y(n_695) );
INVx1_ASAP7_75t_SL g630 ( .A(n_599), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_601), .B(n_629), .Y(n_691) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_606), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g672 ( .A(n_606), .Y(n_672) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_615), .B1(n_617), .B2(n_618), .C(n_620), .Y(n_610) );
NOR2xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_614), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_612), .A2(n_630), .B1(n_676), .B2(n_677), .Y(n_675) );
CKINVDCx14_ASAP7_75t_R g615 ( .A(n_616), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_617), .A2(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR3xp33_ASAP7_75t_SL g623 ( .A(n_624), .B(n_656), .C(n_680), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_625), .B(n_632), .C(n_640), .D(n_647), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g703 ( .A(n_628), .Y(n_703) );
INVx3_ASAP7_75t_SL g697 ( .A(n_629), .Y(n_697) );
OR2x2_ASAP7_75t_L g702 ( .A(n_629), .B(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B1(n_637), .B2(n_639), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_634), .B(n_652), .Y(n_693) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B(n_644), .Y(n_640) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_659), .B(n_662), .C(n_675), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g690 ( .A(n_661), .Y(n_690) );
AOI222xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_667), .B1(n_668), .B2(n_671), .C1(n_673), .C2(n_674), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND4xp25_ASAP7_75t_SL g699 ( .A(n_672), .B(n_700), .C(n_701), .D(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g680 ( .A(n_681), .B(n_689), .C(n_698), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_698) );
INVx1_ASAP7_75t_L g719 ( .A(n_709), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_710), .Y(n_720) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
endmodule