module real_jpeg_20582_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_0),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_55),
.Y(n_167)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_66),
.B1(n_73),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_3),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_54),
.B1(n_56),
.B2(n_96),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_96),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_96),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_48),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_5),
.A2(n_66),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_54),
.B1(n_56),
.B2(n_74),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_74),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_74),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_6),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_6),
.A2(n_54),
.B(n_71),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_6),
.A2(n_66),
.B1(n_73),
.B2(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_6),
.B(n_76),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_38),
.B(n_42),
.C(n_177),
.D(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_6),
.B(n_38),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_60),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_6),
.A2(n_26),
.B(n_192),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_6),
.A2(n_56),
.B(n_57),
.C(n_126),
.D(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_6),
.B(n_56),
.Y(n_224)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_8),
.B(n_193),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_66),
.B1(n_73),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_11),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_11),
.A2(n_54),
.B1(n_56),
.B2(n_78),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_78),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_78),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_12),
.A2(n_40),
.B1(n_54),
.B2(n_56),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_40),
.Y(n_120)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_104),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_79),
.B2(n_80),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_25),
.B(n_36),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_34),
.B(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_26),
.A2(n_83),
.B1(n_90),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_26),
.A2(n_83),
.B1(n_120),
.B2(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_26),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_26),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_27),
.A2(n_198),
.B(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_30),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_28),
.A2(n_44),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_30),
.B(n_43),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_30),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_32),
.A2(n_167),
.B(n_207),
.Y(n_231)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_39),
.B1(n_58),
.B2(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_38),
.B(n_58),
.Y(n_230)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_43),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_39),
.A2(n_59),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_41),
.A2(n_49),
.B1(n_189),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_41),
.A2(n_222),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_42),
.B(n_141),
.Y(n_140)
);

CKINVDCx9p33_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_49),
.A2(n_92),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_49),
.B(n_142),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_49),
.A2(n_140),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_49),
.B(n_117),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_60),
.B2(n_62),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_58),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_56),
.B1(n_68),
.B2(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_72),
.B(n_75),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_70),
.B1(n_72),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_68),
.B(n_117),
.C(n_118),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_95),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_75),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_83),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_83),
.B(n_117),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_97),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_91),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_100),
.A2(n_123),
.B1(n_124),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_100),
.A2(n_101),
.B(n_148),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.C(n_108),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_107),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_109),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_121),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_111),
.B1(n_121),
.B2(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_169),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_152),
.B(n_168),
.Y(n_131)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_132),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_149),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_149),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.C(n_146),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_153),
.B(n_155),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_158),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_162),
.A2(n_163),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_164),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_254),
.C(n_255),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_248),
.B(n_253),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_234),
.B(n_247),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_216),
.B(n_233),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_194),
.B(n_215),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_183),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_175),
.B(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_179),
.B1(n_180),
.B2(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_199),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_204),
.B(n_214),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_202),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_209),
.B(n_213),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_227),
.B2(n_232),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_226),
.C(n_232),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_224),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_227),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_231),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_243),
.C(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);


endmodule