module fake_jpeg_22111_n_30 (n_3, n_2, n_1, n_0, n_4, n_5, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_25;
wire n_17;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_4),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_8),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_13)
);

AND2x6_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_3),
.B1(n_11),
.B2(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_10),
.B(n_11),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_18),
.B1(n_15),
.B2(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_23),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_26),
.A2(n_23),
.B(n_16),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_9),
.B2(n_14),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_10),
.B(n_17),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_9),
.B(n_21),
.Y(n_30)
);


endmodule