module fake_netlist_1_7009_n_1418 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1418);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1418;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_283;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_281;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_1390;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_90), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_159), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_117), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_256), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_202), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_59), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_128), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_218), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_248), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_187), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_229), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_276), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_154), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_26), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_199), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_238), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_190), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_274), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_189), .Y(n_297) );
NOR2xp67_ASAP7_75t_L g298 ( .A(n_136), .B(n_148), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_28), .Y(n_299) );
CKINVDCx16_ASAP7_75t_R g300 ( .A(n_110), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_129), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_79), .B(n_77), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_102), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_260), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_261), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_233), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_249), .Y(n_307) );
INVxp67_ASAP7_75t_SL g308 ( .A(n_105), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_73), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_21), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_58), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_69), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_156), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_213), .Y(n_314) );
BUFx8_ASAP7_75t_SL g315 ( .A(n_120), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_131), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_255), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_184), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_157), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_188), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_30), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_53), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_50), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_97), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_264), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_210), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
INVxp67_ASAP7_75t_SL g328 ( .A(n_69), .Y(n_328) );
CKINVDCx14_ASAP7_75t_R g329 ( .A(n_139), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_253), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_180), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_231), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_114), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_147), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_34), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_246), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_94), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_51), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_192), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_142), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_228), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_83), .Y(n_343) );
NOR2xp67_ASAP7_75t_L g344 ( .A(n_277), .B(n_38), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_197), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_226), .Y(n_346) );
CKINVDCx16_ASAP7_75t_R g347 ( .A(n_209), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_119), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_194), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_271), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_30), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_75), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_245), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_113), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_193), .Y(n_355) );
NOR2xp67_ASAP7_75t_L g356 ( .A(n_214), .B(n_44), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_141), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_121), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_267), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_171), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_0), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_109), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_122), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_200), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_241), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_191), .B(n_109), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_273), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_14), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_222), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_177), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_272), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_243), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_82), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_100), .Y(n_374) );
INVxp33_ASAP7_75t_L g375 ( .A(n_29), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_102), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_26), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_71), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_103), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_2), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_278), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_205), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_225), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_111), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_269), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_0), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_234), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_145), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_169), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_149), .Y(n_390) );
BUFx10_ASAP7_75t_L g391 ( .A(n_179), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_196), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_144), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_125), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_37), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_18), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_237), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_223), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_275), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_132), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_262), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_1), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_160), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_208), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_62), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_44), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_127), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_2), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_203), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_153), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_183), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_236), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_211), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_265), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_124), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_173), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_235), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_257), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_258), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_133), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_29), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_152), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_140), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_88), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_155), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_116), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_60), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_137), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_250), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_263), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_212), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_221), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_176), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_6), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_195), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_130), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_51), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_68), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_87), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_217), .Y(n_440) );
BUFx6f_ASAP7_75t_SL g441 ( .A(n_9), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_110), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_170), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_268), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_299), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_350), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_350), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_299), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_377), .B(n_1), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_350), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_442), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_283), .B(n_3), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_377), .B(n_4), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_279), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_283), .B(n_7), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_283), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_441), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_350), .Y(n_459) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_280), .A2(n_8), .B(n_9), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_350), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_426), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
AND2x6_ASAP7_75t_L g464 ( .A(n_305), .B(n_112), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_391), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_375), .B(n_8), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_312), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_280), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_281), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_340), .B(n_10), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_312), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_360), .B(n_10), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_305), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_371), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_281), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_315), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_337), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_391), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_315), .Y(n_479) );
CKINVDCx6p67_ASAP7_75t_R g480 ( .A(n_371), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_441), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_337), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_383), .B(n_11), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_360), .B(n_11), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_473), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_472), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_453), .A2(n_300), .B1(n_441), .B2(n_282), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_457), .B(n_405), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_452), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_473), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_456), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_456), .B(n_425), .Y(n_492) );
NOR2x1p5_ASAP7_75t_L g493 ( .A(n_479), .B(n_284), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_456), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_465), .B(n_407), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_476), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_457), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_453), .A2(n_452), .B1(n_466), .B2(n_449), .Y(n_499) );
INVx5_ASAP7_75t_L g500 ( .A(n_464), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_465), .B(n_291), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_453), .B(n_313), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_456), .Y(n_503) );
AND2x6_ASAP7_75t_L g504 ( .A(n_452), .B(n_414), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_472), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_473), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_473), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_456), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_481), .B(n_347), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_458), .B(n_425), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_458), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_481), .B(n_391), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_458), .B(n_330), .Y(n_513) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_446), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_458), .B(n_404), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_473), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_458), .B(n_289), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_458), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_465), .B(n_318), .Y(n_519) );
INVx5_ASAP7_75t_L g520 ( .A(n_464), .Y(n_520) );
INVx4_ASAP7_75t_L g521 ( .A(n_452), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_465), .B(n_378), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_452), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_463), .Y(n_524) );
AO22x2_ASAP7_75t_L g525 ( .A1(n_452), .A2(n_366), .B1(n_302), .B2(n_378), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_465), .B(n_389), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_472), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_465), .B(n_443), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_463), .B(n_289), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
INVx5_ASAP7_75t_L g531 ( .A(n_464), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_463), .B(n_306), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_463), .B(n_306), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_476), .B(n_284), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_521), .B(n_472), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_513), .B(n_478), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_498), .B(n_478), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_487), .A2(n_454), .B1(n_311), .B2(n_395), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_502), .A2(n_483), .B1(n_466), .B2(n_484), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_502), .A2(n_483), .B1(n_466), .B2(n_484), .Y(n_540) );
INVx5_ASAP7_75t_L g541 ( .A(n_504), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_525), .A2(n_483), .B1(n_484), .B2(n_478), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_500), .Y(n_543) );
NAND3xp33_ASAP7_75t_SL g544 ( .A(n_487), .B(n_479), .C(n_451), .Y(n_544) );
INVx4_ASAP7_75t_L g545 ( .A(n_521), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_534), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_525), .A2(n_460), .B1(n_484), .B2(n_464), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_493), .B(n_483), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_525), .A2(n_460), .B1(n_484), .B2(n_464), .Y(n_549) );
INVx8_ASAP7_75t_L g550 ( .A(n_504), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_515), .B(n_480), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_525), .A2(n_460), .B1(n_484), .B2(n_464), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_534), .Y(n_553) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_499), .B(n_460), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_521), .B(n_470), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_488), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_515), .B(n_480), .Y(n_557) );
NOR2xp67_ASAP7_75t_L g558 ( .A(n_496), .B(n_463), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_521), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_525), .A2(n_470), .B1(n_451), .B2(n_282), .Y(n_560) );
BUFx3_ASAP7_75t_L g561 ( .A(n_522), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_495), .B(n_480), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_501), .B(n_480), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_488), .B(n_463), .Y(n_564) );
NOR2x2_ASAP7_75t_L g565 ( .A(n_493), .B(n_454), .Y(n_565) );
BUFx3_ASAP7_75t_L g566 ( .A(n_522), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_504), .A2(n_460), .B1(n_464), .B2(n_462), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_L g568 ( .A1(n_530), .A2(n_455), .B(n_302), .C(n_468), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_486), .A2(n_451), .B1(n_363), .B2(n_364), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_486), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_504), .A2(n_297), .B1(n_364), .B2(n_363), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_504), .A2(n_297), .B1(n_416), .B2(n_372), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_486), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_512), .B(n_445), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_500), .B(n_462), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_489), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_522), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_522), .B(n_474), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_519), .B(n_445), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_491), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_504), .A2(n_460), .B1(n_464), .B2(n_462), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_504), .A2(n_416), .B1(n_372), .B2(n_454), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_489), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_489), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_500), .B(n_285), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_505), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_491), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_526), .B(n_445), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_528), .B(n_448), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_517), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_509), .B(n_292), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_503), .B(n_474), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_503), .B(n_474), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_505), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g595 ( .A1(n_505), .A2(n_311), .B1(n_395), .B2(n_279), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_489), .B(n_290), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_523), .B(n_290), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_494), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_500), .B(n_295), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_523), .B(n_295), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_523), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_527), .A2(n_455), .B1(n_321), .B2(n_361), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_523), .B(n_304), .Y(n_603) );
BUFx4f_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_527), .B(n_325), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_527), .B(n_325), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_530), .B(n_334), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_517), .B(n_321), .Y(n_608) );
NAND2xp33_ASAP7_75t_L g609 ( .A(n_500), .B(n_464), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_492), .B(n_336), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_520), .B(n_336), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_492), .B(n_510), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_497), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_497), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_508), .Y(n_615) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_520), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_510), .B(n_345), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_511), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_529), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_511), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_518), .B(n_345), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_518), .B(n_346), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_524), .Y(n_623) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_520), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_524), .B(n_448), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_529), .B(n_346), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_532), .Y(n_627) );
INVx5_ASAP7_75t_L g628 ( .A(n_520), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_532), .A2(n_324), .B1(n_380), .B2(n_361), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_535), .A2(n_533), .B(n_531), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_627), .B(n_533), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_542), .A2(n_468), .B(n_475), .C(n_469), .Y(n_632) );
INVx6_ASAP7_75t_L g633 ( .A(n_537), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_560), .A2(n_324), .B1(n_438), .B2(n_380), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_590), .B(n_438), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_619), .B(n_439), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_561), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_559), .Y(n_638) );
BUFx3_ASAP7_75t_L g639 ( .A(n_556), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_SL g640 ( .A1(n_547), .A2(n_329), .B(n_490), .C(n_485), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_608), .B(n_439), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_539), .A2(n_308), .B1(n_374), .B2(n_351), .C(n_328), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_545), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_540), .B(n_353), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_584), .Y(n_645) );
BUFx2_ASAP7_75t_L g646 ( .A(n_537), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_546), .Y(n_647) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_564), .A2(n_309), .B(n_310), .C(n_303), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_553), .B(n_406), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_566), .Y(n_650) );
INVx4_ASAP7_75t_L g651 ( .A(n_550), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_577), .Y(n_652) );
NOR2xp33_ASAP7_75t_R g653 ( .A(n_544), .B(n_406), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_548), .B(n_421), .Y(n_654) );
AO21x1_ASAP7_75t_L g655 ( .A1(n_579), .A2(n_469), .B(n_468), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_584), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_580), .Y(n_657) );
INVx4_ASAP7_75t_L g658 ( .A(n_550), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_576), .Y(n_659) );
INVx3_ASAP7_75t_L g660 ( .A(n_545), .Y(n_660) );
BUFx3_ASAP7_75t_L g661 ( .A(n_548), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_583), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g663 ( .A(n_582), .B(n_434), .C(n_421), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_569), .A2(n_434), .B1(n_355), .B2(n_358), .Y(n_664) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_541), .B(n_604), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_541), .B(n_520), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_568), .A2(n_323), .B(n_335), .C(n_322), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_554), .A2(n_464), .B1(n_531), .B2(n_343), .Y(n_668) );
AOI221x1_ASAP7_75t_L g669 ( .A1(n_579), .A2(n_473), .B1(n_475), .B2(n_469), .C(n_468), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_588), .A2(n_469), .B(n_475), .C(n_366), .Y(n_670) );
AO32x2_ASAP7_75t_L g671 ( .A1(n_538), .A2(n_473), .A3(n_475), .B1(n_344), .B2(n_356), .Y(n_671) );
BUFx3_ASAP7_75t_L g672 ( .A(n_595), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_554), .A2(n_467), .B1(n_471), .B2(n_448), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_612), .A2(n_531), .B(n_507), .Y(n_674) );
NAND2x1_ASAP7_75t_SL g675 ( .A(n_571), .B(n_298), .Y(n_675) );
OAI21xp33_ASAP7_75t_SL g676 ( .A1(n_547), .A2(n_471), .B(n_467), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_551), .A2(n_531), .B(n_507), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_629), .B(n_467), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_536), .B(n_353), .Y(n_679) );
OAI21xp33_ASAP7_75t_SL g680 ( .A1(n_549), .A2(n_477), .B(n_471), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_549), .A2(n_482), .B1(n_477), .B2(n_338), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_557), .A2(n_531), .B(n_516), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_591), .B(n_352), .Y(n_683) );
INVx3_ASAP7_75t_L g684 ( .A(n_550), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_558), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_626), .B(n_358), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_567), .A2(n_516), .B(n_506), .Y(n_687) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_601), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_604), .B(n_365), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_552), .A2(n_482), .B1(n_373), .B2(n_376), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_610), .B(n_369), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_572), .A2(n_379), .B1(n_384), .B2(n_368), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_570), .B(n_369), .Y(n_694) );
NAND2xp33_ASAP7_75t_R g695 ( .A(n_617), .B(n_370), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_588), .A2(n_386), .B(n_402), .C(n_396), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_587), .Y(n_697) );
BUFx2_ASAP7_75t_L g698 ( .A(n_570), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_563), .A2(n_516), .B(n_506), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_562), .A2(n_382), .B(n_296), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_589), .B(n_408), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_555), .B(n_424), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_602), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_543), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_574), .B(n_427), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_574), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_573), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_573), .B(n_370), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_621), .B(n_437), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_589), .B(n_362), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_565), .A2(n_390), .B1(n_398), .B2(n_381), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g712 ( .A(n_598), .B(n_362), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_622), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_625), .A2(n_287), .B(n_288), .C(n_286), .Y(n_714) );
BUFx12f_ASAP7_75t_L g715 ( .A(n_543), .Y(n_715) );
BUFx3_ASAP7_75t_L g716 ( .A(n_618), .Y(n_716) );
BUFx3_ASAP7_75t_L g717 ( .A(n_625), .Y(n_717) );
INVxp67_ASAP7_75t_L g718 ( .A(n_596), .Y(n_718) );
O2A1O1Ixp33_ASAP7_75t_L g719 ( .A1(n_578), .A2(n_294), .B(n_301), .C(n_293), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_586), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_605), .B(n_606), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_586), .B(n_381), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_592), .A2(n_314), .B(n_307), .Y(n_723) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_543), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_597), .B(n_600), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_613), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_614), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_567), .B(n_473), .C(n_317), .Y(n_728) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_603), .B(n_607), .Y(n_729) );
AND2x4_ASAP7_75t_L g730 ( .A(n_594), .B(n_316), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_594), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_609), .A2(n_398), .B1(n_399), .B2(n_390), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_581), .A2(n_615), .B1(n_623), .B2(n_620), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_593), .A2(n_326), .B(n_320), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_575), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_581), .B(n_399), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_599), .A2(n_423), .B1(n_433), .B2(n_418), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_575), .B(n_423), .Y(n_738) );
BUFx12f_ASAP7_75t_L g739 ( .A(n_543), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_611), .A2(n_331), .B(n_327), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_585), .A2(n_332), .B(n_339), .C(n_333), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_585), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_616), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_616), .A2(n_341), .B(n_348), .C(n_342), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_616), .B(n_319), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_624), .B(n_385), .Y(n_746) );
O2A1O1Ixp33_ASAP7_75t_L g747 ( .A1(n_628), .A2(n_349), .B(n_357), .C(n_354), .Y(n_747) );
INVxp33_ASAP7_75t_SL g748 ( .A(n_628), .Y(n_748) );
NOR2xp33_ASAP7_75t_R g749 ( .A(n_628), .B(n_12), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_560), .A2(n_359), .B1(n_387), .B2(n_367), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_535), .A2(n_392), .B(n_388), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_561), .Y(n_752) );
NOR2xp33_ASAP7_75t_SL g753 ( .A(n_550), .B(n_393), .Y(n_753) );
BUFx12f_ASAP7_75t_L g754 ( .A(n_556), .Y(n_754) );
BUFx2_ASAP7_75t_L g755 ( .A(n_537), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_627), .B(n_394), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_556), .Y(n_757) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_550), .Y(n_758) );
OR2x6_ASAP7_75t_L g759 ( .A(n_550), .B(n_400), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_627), .B(n_401), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_556), .B(n_403), .Y(n_761) );
CKINVDCx8_ASAP7_75t_R g762 ( .A(n_548), .Y(n_762) );
INVx4_ASAP7_75t_L g763 ( .A(n_550), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_560), .A2(n_412), .B1(n_413), .B2(n_410), .Y(n_764) );
OAI22x1_ASAP7_75t_L g765 ( .A1(n_582), .A2(n_417), .B1(n_419), .B2(n_415), .Y(n_765) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_550), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_561), .Y(n_767) );
AND2x4_ASAP7_75t_L g768 ( .A(n_539), .B(n_422), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_560), .A2(n_429), .B1(n_430), .B2(n_428), .Y(n_769) );
O2A1O1Ixp33_ASAP7_75t_L g770 ( .A1(n_556), .A2(n_432), .B(n_436), .C(n_431), .Y(n_770) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_571), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_556), .B(n_444), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_595), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_535), .A2(n_409), .B(n_397), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_631), .B(n_12), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_663), .A2(n_420), .B1(n_435), .B2(n_411), .Y(n_776) );
BUFx2_ASAP7_75t_L g777 ( .A(n_647), .Y(n_777) );
NAND3xp33_ASAP7_75t_SL g778 ( .A(n_713), .B(n_420), .C(n_411), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_699), .A2(n_440), .B(n_435), .Y(n_779) );
AOI221x1_ASAP7_75t_L g780 ( .A1(n_673), .A2(n_461), .B1(n_459), .B2(n_450), .C(n_446), .Y(n_780) );
AO31x2_ASAP7_75t_L g781 ( .A1(n_655), .A2(n_447), .A3(n_440), .B(n_446), .Y(n_781) );
A2O1A1Ixp33_ASAP7_75t_L g782 ( .A1(n_667), .A2(n_447), .B(n_450), .C(n_446), .Y(n_782) );
O2A1O1Ixp5_ASAP7_75t_L g783 ( .A1(n_670), .A2(n_447), .B(n_450), .C(n_446), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_726), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g785 ( .A1(n_642), .A2(n_446), .B1(n_450), .B2(n_459), .C(n_461), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_654), .B(n_13), .Y(n_786) );
O2A1O1Ixp33_ASAP7_75t_SL g787 ( .A1(n_640), .A2(n_632), .B(n_714), .C(n_733), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_664), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_750), .A2(n_461), .B1(n_459), .B2(n_450), .C(n_446), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_677), .A2(n_514), .B(n_450), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_682), .A2(n_514), .B(n_450), .Y(n_791) );
INVx4_ASAP7_75t_SL g792 ( .A(n_754), .Y(n_792) );
OR2x2_ASAP7_75t_L g793 ( .A(n_649), .B(n_16), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g794 ( .A1(n_725), .A2(n_459), .B(n_461), .C(n_446), .Y(n_794) );
O2A1O1Ixp33_ASAP7_75t_L g795 ( .A1(n_696), .A2(n_18), .B(n_16), .C(n_17), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g796 ( .A1(n_719), .A2(n_461), .B(n_459), .C(n_514), .Y(n_796) );
AO21x1_ASAP7_75t_L g797 ( .A1(n_733), .A2(n_461), .B(n_459), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_687), .A2(n_630), .B(n_674), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_651), .B(n_17), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_773), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_750), .A2(n_461), .B1(n_459), .B2(n_514), .C(n_22), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_727), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_L g803 ( .A1(n_721), .A2(n_514), .B(n_21), .C(n_19), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_657), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_702), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_768), .B(n_19), .Y(n_806) );
BUFx8_ASAP7_75t_L g807 ( .A(n_671), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_756), .B(n_635), .Y(n_808) );
NAND2x1p5_ASAP7_75t_L g809 ( .A(n_698), .B(n_20), .Y(n_809) );
O2A1O1Ixp33_ASAP7_75t_L g810 ( .A1(n_648), .A2(n_23), .B(n_20), .C(n_22), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_771), .A2(n_25), .B1(n_23), .B2(n_24), .Y(n_811) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_753), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_703), .A2(n_24), .B1(n_25), .B2(n_27), .Y(n_813) );
A2O1A1Ixp33_ASAP7_75t_L g814 ( .A1(n_676), .A2(n_27), .B(n_28), .C(n_31), .Y(n_814) );
BUFx2_ASAP7_75t_R g815 ( .A(n_762), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_759), .A2(n_756), .B1(n_691), .B2(n_681), .Y(n_816) );
A2O1A1Ixp33_ASAP7_75t_L g817 ( .A1(n_680), .A2(n_31), .B(n_32), .C(n_33), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_697), .Y(n_818) );
BUFx8_ASAP7_75t_L g819 ( .A(n_671), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_764), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_820) );
A2O1A1Ixp33_ASAP7_75t_L g821 ( .A1(n_709), .A2(n_35), .B(n_36), .C(n_37), .Y(n_821) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_634), .A2(n_35), .B1(n_36), .B2(n_38), .C(n_39), .Y(n_822) );
AOI21xp5_ASAP7_75t_L g823 ( .A1(n_729), .A2(n_118), .B(n_115), .Y(n_823) );
AO31x2_ASAP7_75t_L g824 ( .A1(n_669), .A2(n_39), .A3(n_40), .B(n_41), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_718), .A2(n_736), .B(n_686), .Y(n_825) );
A2O1A1Ixp33_ASAP7_75t_L g826 ( .A1(n_705), .A2(n_41), .B(n_42), .C(n_43), .Y(n_826) );
O2A1O1Ixp33_ASAP7_75t_L g827 ( .A1(n_764), .A2(n_42), .B(n_43), .C(n_45), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_636), .B(n_46), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_768), .B(n_46), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_692), .A2(n_126), .B(n_123), .Y(n_830) );
INVx2_ASAP7_75t_SL g831 ( .A(n_639), .Y(n_831) );
CKINVDCx12_ASAP7_75t_R g832 ( .A(n_759), .Y(n_832) );
AND2x4_ASAP7_75t_L g833 ( .A(n_651), .B(n_658), .Y(n_833) );
CKINVDCx9p33_ASAP7_75t_R g834 ( .A(n_722), .Y(n_834) );
AND2x2_ASAP7_75t_SL g835 ( .A(n_753), .B(n_47), .Y(n_835) );
BUFx8_ASAP7_75t_L g836 ( .A(n_671), .Y(n_836) );
OAI21xp5_ASAP7_75t_L g837 ( .A1(n_728), .A2(n_135), .B(n_134), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_702), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g839 ( .A(n_653), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g840 ( .A(n_683), .B(n_48), .C(n_49), .Y(n_840) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_701), .A2(n_143), .B(n_138), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_711), .A2(n_48), .B1(n_49), .B2(n_50), .C(n_52), .Y(n_842) );
A2O1A1Ixp33_ASAP7_75t_L g843 ( .A1(n_770), .A2(n_52), .B(n_53), .C(n_54), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_769), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_844) );
BUFx12f_ASAP7_75t_L g845 ( .A(n_757), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_715), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_701), .A2(n_150), .B(n_146), .Y(n_847) );
O2A1O1Ixp33_ASAP7_75t_L g848 ( .A1(n_769), .A2(n_55), .B(n_56), .C(n_57), .Y(n_848) );
AND2x4_ASAP7_75t_L g849 ( .A(n_658), .B(n_57), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_638), .Y(n_850) );
INVx4_ASAP7_75t_L g851 ( .A(n_739), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_L g852 ( .A1(n_751), .A2(n_58), .B(n_59), .C(n_60), .Y(n_852) );
AO32x2_ASAP7_75t_L g853 ( .A1(n_673), .A2(n_61), .A3(n_62), .B1(n_63), .B2(n_64), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_661), .B(n_61), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_760), .B(n_63), .Y(n_855) );
O2A1O1Ixp33_ASAP7_75t_L g856 ( .A1(n_693), .A2(n_64), .B(n_65), .C(n_66), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_700), .A2(n_186), .B(n_270), .Y(n_857) );
INVx5_ASAP7_75t_L g858 ( .A(n_759), .Y(n_858) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_704), .Y(n_859) );
OAI21xp5_ASAP7_75t_L g860 ( .A1(n_668), .A2(n_185), .B(n_266), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_693), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_861) );
INVx1_ASAP7_75t_SL g862 ( .A(n_707), .Y(n_862) );
NOR2xp67_ASAP7_75t_L g863 ( .A(n_765), .B(n_67), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_712), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_678), .B(n_68), .Y(n_865) );
AO31x2_ASAP7_75t_L g866 ( .A1(n_774), .A2(n_70), .A3(n_72), .B(n_73), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_720), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_641), .B(n_70), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_695), .Y(n_869) );
BUFx2_ASAP7_75t_L g870 ( .A(n_749), .Y(n_870) );
BUFx6f_ASAP7_75t_L g871 ( .A(n_704), .Y(n_871) );
INVx2_ASAP7_75t_SL g872 ( .A(n_730), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_659), .Y(n_873) );
OAI21x1_ASAP7_75t_L g874 ( .A1(n_712), .A2(n_182), .B(n_259), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_731), .Y(n_875) );
A2O1A1Ixp33_ASAP7_75t_L g876 ( .A1(n_706), .A2(n_72), .B(n_74), .C(n_75), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_717), .B(n_74), .Y(n_877) );
CKINVDCx12_ASAP7_75t_R g878 ( .A(n_738), .Y(n_878) );
AO32x2_ASAP7_75t_L g879 ( .A1(n_675), .A2(n_76), .A3(n_77), .B1(n_78), .B2(n_79), .Y(n_879) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_723), .A2(n_76), .B(n_78), .C(n_80), .Y(n_880) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_644), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_710), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_734), .A2(n_81), .B(n_83), .C(n_84), .Y(n_883) );
O2A1O1Ixp33_ASAP7_75t_L g884 ( .A1(n_761), .A2(n_84), .B(n_85), .C(n_86), .Y(n_884) );
BUFx2_ASAP7_75t_L g885 ( .A(n_633), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_662), .Y(n_886) );
BUFx3_ASAP7_75t_L g887 ( .A(n_716), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_772), .B(n_85), .Y(n_888) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_679), .A2(n_198), .B(n_254), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_742), .Y(n_890) );
O2A1O1Ixp33_ASAP7_75t_L g891 ( .A1(n_744), .A2(n_86), .B(n_87), .C(n_88), .Y(n_891) );
AO31x2_ASAP7_75t_L g892 ( .A1(n_646), .A2(n_755), .A3(n_689), .B(n_740), .Y(n_892) );
BUFx2_ASAP7_75t_L g893 ( .A(n_633), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_746), .A2(n_201), .B(n_252), .Y(n_894) );
O2A1O1Ixp33_ASAP7_75t_L g895 ( .A1(n_747), .A2(n_89), .B(n_90), .C(n_91), .Y(n_895) );
INVx1_ASAP7_75t_SL g896 ( .A(n_694), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_656), .A2(n_204), .B(n_251), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_643), .Y(n_898) );
INVx3_ASAP7_75t_L g899 ( .A(n_763), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_637), .B(n_91), .Y(n_900) );
INVx3_ASAP7_75t_L g901 ( .A(n_763), .Y(n_901) );
BUFx3_ASAP7_75t_L g902 ( .A(n_748), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_650), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_903) );
INVx2_ASAP7_75t_L g904 ( .A(n_643), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_652), .A2(n_92), .B1(n_93), .B2(n_95), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_660), .Y(n_906) );
BUFx2_ASAP7_75t_SL g907 ( .A(n_758), .Y(n_907) );
INVx2_ASAP7_75t_SL g908 ( .A(n_685), .Y(n_908) );
AO31x2_ASAP7_75t_L g909 ( .A1(n_735), .A2(n_95), .A3(n_96), .B(n_97), .Y(n_909) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_737), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_660), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g912 ( .A1(n_708), .A2(n_206), .B(n_247), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_752), .B(n_96), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_645), .Y(n_914) );
O2A1O1Ixp33_ASAP7_75t_L g915 ( .A1(n_741), .A2(n_98), .B(n_99), .C(n_100), .Y(n_915) );
A2O1A1Ixp33_ASAP7_75t_L g916 ( .A1(n_745), .A2(n_98), .B(n_99), .C(n_101), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_767), .Y(n_917) );
O2A1O1Ixp33_ASAP7_75t_L g918 ( .A1(n_690), .A2(n_101), .B(n_103), .C(n_104), .Y(n_918) );
AO31x2_ASAP7_75t_L g919 ( .A1(n_743), .A2(n_704), .A3(n_724), .B(n_732), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_665), .Y(n_920) );
INVx5_ASAP7_75t_L g921 ( .A(n_758), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_666), .A2(n_207), .B(n_244), .Y(n_922) );
BUFx12f_ASAP7_75t_L g923 ( .A(n_766), .Y(n_923) );
CKINVDCx6p67_ASAP7_75t_R g924 ( .A(n_766), .Y(n_924) );
O2A1O1Ixp33_ASAP7_75t_L g925 ( .A1(n_684), .A2(n_104), .B(n_105), .C(n_106), .Y(n_925) );
O2A1O1Ixp33_ASAP7_75t_L g926 ( .A1(n_766), .A2(n_106), .B(n_107), .C(n_108), .Y(n_926) );
AO32x2_ASAP7_75t_L g927 ( .A1(n_724), .A2(n_107), .A3(n_108), .B1(n_111), .B2(n_151), .Y(n_927) );
A2O1A1Ixp33_ASAP7_75t_L g928 ( .A1(n_688), .A2(n_158), .B(n_161), .C(n_162), .Y(n_928) );
OAI21xp5_ASAP7_75t_L g929 ( .A1(n_783), .A2(n_688), .B(n_164), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_804), .Y(n_930) );
AOI21xp33_ASAP7_75t_L g931 ( .A1(n_816), .A2(n_163), .B(n_165), .Y(n_931) );
AO21x1_ASAP7_75t_L g932 ( .A1(n_812), .A2(n_166), .B(n_167), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_862), .B(n_168), .Y(n_933) );
NAND2xp5_ASAP7_75t_SL g934 ( .A(n_858), .B(n_172), .Y(n_934) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_808), .A2(n_174), .B1(n_175), .B2(n_178), .C(n_181), .Y(n_935) );
INVx3_ASAP7_75t_L g936 ( .A(n_833), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_867), .B(n_215), .Y(n_937) );
BUFx6f_ASAP7_75t_L g938 ( .A(n_859), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_818), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_818), .B(n_216), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_777), .B(n_219), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_784), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_882), .B(n_220), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_846), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_875), .B(n_224), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_832), .Y(n_946) );
O2A1O1Ixp33_ASAP7_75t_L g947 ( .A1(n_795), .A2(n_227), .B(n_230), .C(n_232), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_802), .Y(n_948) );
HB1xp67_ASAP7_75t_L g949 ( .A(n_851), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_917), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_917), .Y(n_951) );
INVxp67_ASAP7_75t_L g952 ( .A(n_815), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_793), .B(n_239), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_805), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_838), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_872), .B(n_887), .Y(n_956) );
INVx3_ASAP7_75t_L g957 ( .A(n_833), .Y(n_957) );
OR2x6_ASAP7_75t_L g958 ( .A(n_851), .B(n_799), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_828), .Y(n_959) );
NOR2xp67_ASAP7_75t_L g960 ( .A(n_858), .B(n_845), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_900), .Y(n_961) );
BUFx2_ASAP7_75t_L g962 ( .A(n_923), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_865), .B(n_775), .Y(n_963) );
AO21x2_ASAP7_75t_L g964 ( .A1(n_797), .A2(n_837), .B(n_794), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_809), .Y(n_965) );
OR2x2_ASAP7_75t_L g966 ( .A(n_890), .B(n_806), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_790), .A2(n_791), .B(n_779), .Y(n_967) );
OAI21xp5_ASAP7_75t_L g968 ( .A1(n_782), .A2(n_796), .B(n_803), .Y(n_968) );
OAI21xp33_ASAP7_75t_SL g969 ( .A1(n_835), .A2(n_863), .B(n_874), .Y(n_969) );
AND2x4_ASAP7_75t_L g970 ( .A(n_858), .B(n_864), .Y(n_970) );
NAND2xp5_ASAP7_75t_SL g971 ( .A(n_799), .B(n_849), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_902), .B(n_877), .Y(n_972) );
NAND2xp5_ASAP7_75t_SL g973 ( .A(n_849), .B(n_870), .Y(n_973) );
AOI21xp5_ASAP7_75t_L g974 ( .A1(n_860), .A2(n_830), .B(n_889), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_829), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_861), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_873), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_850), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_886), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_910), .A2(n_786), .B1(n_778), .B2(n_855), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_868), .B(n_888), .Y(n_981) );
AOI221xp5_ASAP7_75t_L g982 ( .A1(n_788), .A2(n_856), .B1(n_822), .B2(n_848), .C(n_827), .Y(n_982) );
INVx2_ASAP7_75t_SL g983 ( .A(n_792), .Y(n_983) );
BUFx3_ASAP7_75t_L g984 ( .A(n_924), .Y(n_984) );
AOI21xp5_ASAP7_75t_L g985 ( .A1(n_894), .A2(n_780), .B(n_823), .Y(n_985) );
BUFx6f_ASAP7_75t_L g986 ( .A(n_859), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_776), .A2(n_854), .B1(n_839), .B2(n_913), .Y(n_987) );
BUFx3_ASAP7_75t_L g988 ( .A(n_831), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_807), .A2(n_819), .B1(n_836), .B2(n_869), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_857), .A2(n_847), .B(n_841), .Y(n_990) );
BUFx4f_ASAP7_75t_SL g991 ( .A(n_792), .Y(n_991) );
A2O1A1Ixp33_ASAP7_75t_L g992 ( .A1(n_810), .A2(n_915), .B(n_895), .C(n_884), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_866), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_866), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_842), .A2(n_807), .B1(n_819), .B2(n_836), .Y(n_995) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_878), .Y(n_996) );
INVx3_ASAP7_75t_L g997 ( .A(n_921), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_921), .Y(n_998) );
NOR2x1_ASAP7_75t_SL g999 ( .A(n_921), .B(n_907), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_881), .A2(n_844), .B1(n_785), .B2(n_821), .C(n_826), .Y(n_1000) );
AOI22xp5_ASAP7_75t_L g1001 ( .A1(n_896), .A2(n_800), .B1(n_820), .B2(n_811), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_914), .B(n_920), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_898), .B(n_906), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_840), .A2(n_893), .B1(n_885), .B2(n_908), .Y(n_1004) );
BUFx6f_ASAP7_75t_L g1005 ( .A(n_859), .Y(n_1005) );
OAI211xp5_ASAP7_75t_L g1006 ( .A1(n_813), .A2(n_903), .B(n_925), .C(n_905), .Y(n_1006) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_891), .A2(n_843), .B1(n_817), .B2(n_814), .C(n_801), .Y(n_1007) );
A2O1A1Ixp33_ASAP7_75t_L g1008 ( .A1(n_918), .A2(n_926), .B(n_916), .C(n_883), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_899), .Y(n_1009) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_899), .B(n_901), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_911), .B(n_853), .Y(n_1011) );
OA21x2_ASAP7_75t_L g1012 ( .A1(n_897), .A2(n_789), .B(n_912), .Y(n_1012) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_904), .B(n_901), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_853), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_853), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_909), .Y(n_1016) );
OR2x6_ASAP7_75t_L g1017 ( .A(n_871), .B(n_876), .Y(n_1017) );
A2O1A1Ixp33_ASAP7_75t_L g1018 ( .A1(n_880), .A2(n_852), .B(n_922), .C(n_928), .Y(n_1018) );
A2O1A1Ixp33_ASAP7_75t_L g1019 ( .A1(n_879), .A2(n_834), .B(n_927), .C(n_824), .Y(n_1019) );
HB1xp67_ASAP7_75t_L g1020 ( .A(n_892), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_927), .A2(n_879), .B1(n_824), .B2(n_892), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_781), .B(n_892), .Y(n_1022) );
INVx2_ASAP7_75t_L g1023 ( .A(n_824), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_879), .A2(n_927), .B1(n_919), .B2(n_909), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_919), .A2(n_595), .B1(n_544), .B2(n_627), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_909), .B(n_919), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_804), .Y(n_1027) );
OAI21xp33_ASAP7_75t_L g1028 ( .A1(n_835), .A2(n_502), .B(n_487), .Y(n_1028) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_804), .Y(n_1030) );
BUFx12f_ASAP7_75t_SL g1031 ( .A(n_851), .Y(n_1031) );
INVx4_ASAP7_75t_SL g1032 ( .A(n_923), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_846), .Y(n_1033) );
AOI21xp5_ASAP7_75t_L g1034 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1034) );
INVx1_ASAP7_75t_SL g1035 ( .A(n_862), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_816), .A2(n_544), .B1(n_538), .B2(n_672), .Y(n_1036) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_846), .Y(n_1037) );
AOI22xp5_ASAP7_75t_L g1038 ( .A1(n_816), .A2(n_595), .B1(n_544), .B2(n_627), .Y(n_1038) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_846), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_818), .B(n_808), .Y(n_1040) );
BUFx3_ASAP7_75t_L g1041 ( .A(n_846), .Y(n_1041) );
OAI21xp5_ASAP7_75t_L g1042 ( .A1(n_783), .A2(n_728), .B(n_733), .Y(n_1042) );
AOI21xp5_ASAP7_75t_L g1043 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_816), .A2(n_544), .B1(n_538), .B2(n_672), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_804), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_816), .A2(n_835), .B1(n_812), .B2(n_858), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_846), .Y(n_1047) );
AOI21xp5_ASAP7_75t_L g1048 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_816), .A2(n_544), .B1(n_538), .B2(n_672), .Y(n_1049) );
AOI21xp5_ASAP7_75t_L g1050 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_862), .B(n_546), .Y(n_1051) );
INVx2_ASAP7_75t_L g1052 ( .A(n_804), .Y(n_1052) );
CKINVDCx6p67_ASAP7_75t_R g1053 ( .A(n_832), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_818), .B(n_808), .Y(n_1054) );
AOI21xp5_ASAP7_75t_L g1055 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_804), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_804), .Y(n_1057) );
AOI21xp5_ASAP7_75t_L g1058 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1058) );
AOI21xp33_ASAP7_75t_L g1059 ( .A1(n_816), .A2(n_835), .B(n_673), .Y(n_1059) );
INVxp67_ASAP7_75t_L g1060 ( .A(n_777), .Y(n_1060) );
NAND2xp5_ASAP7_75t_SL g1061 ( .A(n_858), .B(n_835), .Y(n_1061) );
AOI21xp5_ASAP7_75t_L g1062 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_816), .A2(n_544), .B1(n_538), .B2(n_672), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_862), .B(n_546), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_804), .Y(n_1065) );
AO22x1_ASAP7_75t_L g1066 ( .A1(n_858), .A2(n_869), .B1(n_870), .B2(n_849), .Y(n_1066) );
AOI21xp5_ASAP7_75t_L g1067 ( .A1(n_798), .A2(n_787), .B(n_825), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_1028), .A2(n_1049), .B1(n_1063), .B2(n_1044), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1069 ( .A(n_1001), .B(n_966), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_950), .Y(n_1070) );
OAI21xp5_ASAP7_75t_L g1071 ( .A1(n_992), .A2(n_1008), .B(n_1038), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1036), .B(n_1040), .Y(n_1072) );
AO21x2_ASAP7_75t_L g1073 ( .A1(n_1029), .A2(n_1043), .B(n_1034), .Y(n_1073) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_1020), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_951), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1054), .B(n_976), .Y(n_1076) );
OR2x6_ASAP7_75t_L g1077 ( .A(n_958), .B(n_971), .Y(n_1077) );
BUFx4f_ASAP7_75t_SL g1078 ( .A(n_944), .Y(n_1078) );
AND2x4_ASAP7_75t_L g1079 ( .A(n_970), .B(n_938), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1027), .Y(n_1080) );
OR2x6_ASAP7_75t_L g1081 ( .A(n_958), .B(n_1046), .Y(n_1081) );
INVxp67_ASAP7_75t_SL g1082 ( .A(n_1002), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_959), .B(n_975), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_980), .B(n_1035), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_930), .B(n_1030), .Y(n_1085) );
CKINVDCx20_ASAP7_75t_R g1086 ( .A(n_991), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_1035), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1052), .B(n_1065), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_942), .B(n_1045), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_993), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1056), .B(n_1057), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_994), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_1031), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_978), .B(n_948), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_977), .B(n_979), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1051), .B(n_1064), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1002), .B(n_954), .Y(n_1097) );
AO31x2_ASAP7_75t_L g1098 ( .A1(n_1021), .A2(n_1062), .A3(n_1058), .B(n_1055), .Y(n_1098) );
AO21x2_ASAP7_75t_L g1099 ( .A1(n_1048), .A2(n_1067), .B(n_1050), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_955), .B(n_961), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_936), .B(n_957), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1016), .Y(n_1102) );
OAI221xp5_ASAP7_75t_SL g1103 ( .A1(n_1025), .A2(n_995), .B1(n_958), .B2(n_982), .C(n_981), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1014), .B(n_1015), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_936), .B(n_957), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1106 ( .A1(n_1046), .A2(n_989), .B1(n_1059), .B2(n_1061), .Y(n_1106) );
OA21x2_ASAP7_75t_L g1107 ( .A1(n_1024), .A2(n_1022), .B(n_1023), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_970), .B(n_938), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_963), .B(n_1011), .Y(n_1109) );
OA21x2_ASAP7_75t_L g1110 ( .A1(n_1022), .A2(n_1019), .B(n_1026), .Y(n_1110) );
AND2x4_ASAP7_75t_L g1111 ( .A(n_938), .B(n_986), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_984), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_963), .B(n_1059), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1009), .B(n_1010), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_969), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_1033), .Y(n_1116) );
OA21x2_ASAP7_75t_L g1117 ( .A1(n_1042), .A2(n_967), .B(n_985), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1009), .B(n_1010), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_940), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_953), .B(n_981), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_940), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_972), .B(n_1060), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g1123 ( .A(n_999), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_982), .A2(n_1000), .B1(n_987), .B2(n_965), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g1125 ( .A1(n_935), .A2(n_1006), .B1(n_1039), .B2(n_1037), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_1003), .B(n_998), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1003), .B(n_973), .Y(n_1127) );
INVx3_ASAP7_75t_L g1128 ( .A(n_986), .Y(n_1128) );
OA21x2_ASAP7_75t_L g1129 ( .A1(n_968), .A2(n_929), .B(n_931), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_997), .B(n_943), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_943), .Y(n_1131) );
AO21x2_ASAP7_75t_L g1132 ( .A1(n_964), .A2(n_974), .B(n_990), .Y(n_1132) );
OAI21xp5_ASAP7_75t_L g1133 ( .A1(n_1018), .A2(n_1000), .B(n_1007), .Y(n_1133) );
INVxp67_ASAP7_75t_L g1134 ( .A(n_962), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_997), .B(n_937), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_1041), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1017), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_945), .B(n_1013), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1004), .B(n_1007), .Y(n_1139) );
BUFx3_ASAP7_75t_L g1140 ( .A(n_1047), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_941), .B(n_1005), .Y(n_1141) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_946), .B(n_1053), .Y(n_1142) );
OAI211xp5_ASAP7_75t_SL g1143 ( .A1(n_952), .A2(n_949), .B(n_996), .C(n_983), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_956), .B(n_1066), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1005), .B(n_933), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1005), .B(n_1017), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_935), .A2(n_988), .B1(n_1017), .B2(n_960), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_964), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_932), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1032), .B(n_947), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_1032), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1012), .Y(n_1152) );
INVx3_ASAP7_75t_L g1153 ( .A(n_1012), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_934), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1032), .Y(n_1155) );
OA21x2_ASAP7_75t_L g1156 ( .A1(n_1029), .A2(n_1043), .B(n_1034), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1157 ( .A(n_939), .B(n_950), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_930), .B(n_1030), .Y(n_1158) );
AO21x2_ASAP7_75t_L g1159 ( .A1(n_1029), .A2(n_1043), .B(n_1034), .Y(n_1159) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_1028), .A2(n_538), .B1(n_1038), .B2(n_1036), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1161 ( .A(n_939), .B(n_950), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_939), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_930), .B(n_1030), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_930), .B(n_1030), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1102), .Y(n_1165) );
AOI33xp33_ASAP7_75t_L g1166 ( .A1(n_1068), .A2(n_1124), .A3(n_1160), .B1(n_1139), .B2(n_1125), .B3(n_1100), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1109), .B(n_1113), .Y(n_1167) );
BUFx6f_ASAP7_75t_L g1168 ( .A(n_1111), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1109), .B(n_1113), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1102), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1090), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1070), .B(n_1075), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1070), .B(n_1075), .Y(n_1173) );
OAI21xp5_ASAP7_75t_L g1174 ( .A1(n_1071), .A2(n_1133), .B(n_1139), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1090), .Y(n_1175) );
INVxp67_ASAP7_75t_SL g1176 ( .A(n_1082), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1092), .Y(n_1177) );
BUFx2_ASAP7_75t_L g1178 ( .A(n_1074), .Y(n_1178) );
HB1xp67_ASAP7_75t_L g1179 ( .A(n_1126), .Y(n_1179) );
INVxp67_ASAP7_75t_SL g1180 ( .A(n_1074), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1162), .B(n_1157), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1157), .B(n_1161), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1157), .B(n_1161), .Y(n_1183) );
INVx1_ASAP7_75t_SL g1184 ( .A(n_1078), .Y(n_1184) );
NOR2xp67_ASAP7_75t_L g1185 ( .A(n_1106), .B(n_1137), .Y(n_1185) );
AND2x4_ASAP7_75t_L g1186 ( .A(n_1081), .B(n_1137), .Y(n_1186) );
AOI221xp5_ASAP7_75t_L g1187 ( .A1(n_1103), .A2(n_1069), .B1(n_1072), .B2(n_1076), .C(n_1084), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_1081), .A2(n_1138), .B1(n_1147), .B2(n_1077), .Y(n_1188) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_1081), .A2(n_1120), .B1(n_1131), .B2(n_1077), .Y(n_1189) );
INVx2_ASAP7_75t_SL g1190 ( .A(n_1079), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1161), .B(n_1095), .Y(n_1191) );
OAI33xp33_ASAP7_75t_L g1192 ( .A1(n_1083), .A2(n_1143), .A3(n_1096), .B1(n_1122), .B2(n_1120), .B3(n_1144), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1104), .Y(n_1193) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_1126), .Y(n_1194) );
BUFx6f_ASAP7_75t_L g1195 ( .A(n_1111), .Y(n_1195) );
INVx2_ASAP7_75t_SL g1196 ( .A(n_1079), .Y(n_1196) );
HB1xp67_ASAP7_75t_L g1197 ( .A(n_1116), .Y(n_1197) );
INVxp67_ASAP7_75t_L g1198 ( .A(n_1136), .Y(n_1198) );
AND2x4_ASAP7_75t_L g1199 ( .A(n_1081), .B(n_1146), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1107), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1097), .B(n_1100), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1087), .B(n_1127), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1095), .B(n_1085), .Y(n_1203) );
AND2x4_ASAP7_75t_L g1204 ( .A(n_1146), .B(n_1115), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1085), .B(n_1088), .Y(n_1205) );
OAI33xp33_ASAP7_75t_L g1206 ( .A1(n_1134), .A2(n_1155), .A3(n_1080), .B1(n_1127), .B2(n_1091), .B3(n_1148), .Y(n_1206) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1156), .Y(n_1207) );
NOR2x1_ASAP7_75t_L g1208 ( .A(n_1077), .B(n_1150), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1088), .B(n_1164), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1158), .B(n_1164), .Y(n_1210) );
INVxp67_ASAP7_75t_L g1211 ( .A(n_1140), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1097), .B(n_1089), .Y(n_1212) );
BUFx2_ASAP7_75t_L g1213 ( .A(n_1111), .Y(n_1213) );
AND2x2_ASAP7_75t_SL g1214 ( .A(n_1115), .B(n_1129), .Y(n_1214) );
BUFx2_ASAP7_75t_L g1215 ( .A(n_1077), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1216 ( .A(n_1158), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1163), .Y(n_1217) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_1140), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1094), .B(n_1138), .Y(n_1219) );
OAI33xp33_ASAP7_75t_L g1220 ( .A1(n_1155), .A2(n_1148), .A3(n_1093), .B1(n_1149), .B2(n_1131), .B3(n_1119), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1094), .B(n_1135), .Y(n_1221) );
INVx4_ASAP7_75t_L g1222 ( .A(n_1079), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1110), .B(n_1121), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1141), .B(n_1119), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1167), .B(n_1152), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1167), .B(n_1152), .Y(n_1226) );
OAI21xp5_ASAP7_75t_L g1227 ( .A1(n_1174), .A2(n_1123), .B(n_1121), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1178), .Y(n_1228) );
INVxp67_ASAP7_75t_L g1229 ( .A(n_1178), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1169), .B(n_1153), .Y(n_1230) );
AND2x4_ASAP7_75t_L g1231 ( .A(n_1186), .B(n_1098), .Y(n_1231) );
AND2x2_ASAP7_75t_SL g1232 ( .A(n_1214), .B(n_1129), .Y(n_1232) );
INVxp67_ASAP7_75t_SL g1233 ( .A(n_1176), .Y(n_1233) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_1180), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1165), .Y(n_1235) );
AND2x4_ASAP7_75t_L g1236 ( .A(n_1186), .B(n_1098), .Y(n_1236) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1169), .B(n_1098), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1223), .B(n_1117), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1165), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1223), .B(n_1117), .Y(n_1240) );
BUFx2_ASAP7_75t_L g1241 ( .A(n_1213), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1170), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_1187), .A2(n_1135), .B1(n_1101), .B2(n_1105), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1193), .B(n_1130), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1170), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1171), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1202), .B(n_1098), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1202), .B(n_1098), .Y(n_1248) );
AND2x4_ASAP7_75t_L g1249 ( .A(n_1186), .B(n_1132), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1172), .B(n_1130), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1179), .B(n_1073), .Y(n_1251) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1207), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1200), .B(n_1073), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1175), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1175), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1172), .B(n_1159), .Y(n_1256) );
AND2x4_ASAP7_75t_SL g1257 ( .A(n_1182), .B(n_1108), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1177), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1173), .B(n_1159), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1204), .B(n_1099), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1230), .B(n_1204), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1230), .B(n_1204), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1235), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1230), .B(n_1204), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1250), .B(n_1194), .Y(n_1265) );
AOI22xp5_ASAP7_75t_L g1266 ( .A1(n_1243), .A2(n_1192), .B1(n_1185), .B2(n_1188), .Y(n_1266) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1252), .Y(n_1267) );
OR2x2_ASAP7_75t_L g1268 ( .A(n_1250), .B(n_1219), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1244), .B(n_1216), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1225), .B(n_1191), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1235), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1244), .B(n_1217), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1225), .B(n_1203), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1239), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1225), .B(n_1203), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1239), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1242), .Y(n_1277) );
OAI21xp33_ASAP7_75t_L g1278 ( .A1(n_1237), .A2(n_1166), .B(n_1214), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1226), .B(n_1205), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1233), .B(n_1201), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1226), .B(n_1191), .Y(n_1281) );
OR2x6_ASAP7_75t_L g1282 ( .A(n_1227), .B(n_1208), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1242), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1233), .B(n_1212), .Y(n_1284) );
OAI21xp5_ASAP7_75t_SL g1285 ( .A1(n_1243), .A2(n_1151), .B(n_1189), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1226), .B(n_1205), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1245), .B(n_1209), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1245), .B(n_1209), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1237), .B(n_1210), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1237), .B(n_1210), .Y(n_1290) );
AND2x4_ASAP7_75t_L g1291 ( .A(n_1249), .B(n_1186), .Y(n_1291) );
INVx2_ASAP7_75t_SL g1292 ( .A(n_1257), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1246), .B(n_1197), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1238), .B(n_1214), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1247), .B(n_1224), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1234), .B(n_1224), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1238), .B(n_1181), .Y(n_1297) );
NAND2xp5_ASAP7_75t_SL g1298 ( .A(n_1227), .B(n_1185), .Y(n_1298) );
INVxp33_ASAP7_75t_L g1299 ( .A(n_1234), .Y(n_1299) );
INVx1_ASAP7_75t_SL g1300 ( .A(n_1257), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1247), .B(n_1221), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1254), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1294), .B(n_1260), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1263), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1289), .B(n_1248), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1271), .Y(n_1306) );
NOR2xp33_ASAP7_75t_L g1307 ( .A(n_1268), .B(n_1211), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1294), .B(n_1260), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1280), .B(n_1238), .Y(n_1309) );
AOI22xp5_ASAP7_75t_L g1310 ( .A1(n_1266), .A2(n_1189), .B1(n_1183), .B2(n_1182), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1297), .B(n_1260), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1297), .B(n_1240), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1284), .B(n_1240), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1273), .B(n_1240), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1274), .Y(n_1315) );
INVxp67_ASAP7_75t_L g1316 ( .A(n_1296), .Y(n_1316) );
INVxp67_ASAP7_75t_L g1317 ( .A(n_1293), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1270), .B(n_1231), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1265), .B(n_1218), .Y(n_1319) );
NAND4xp25_ASAP7_75t_L g1320 ( .A(n_1278), .B(n_1285), .C(n_1298), .D(n_1208), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1275), .B(n_1256), .Y(n_1321) );
NAND2xp5_ASAP7_75t_SL g1322 ( .A(n_1299), .B(n_1198), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1270), .B(n_1231), .Y(n_1323) );
AND2x2_ASAP7_75t_SL g1324 ( .A(n_1295), .B(n_1257), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1281), .B(n_1256), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1281), .B(n_1259), .Y(n_1326) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1290), .B(n_1248), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1276), .Y(n_1328) );
INVx2_ASAP7_75t_L g1329 ( .A(n_1267), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1277), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1261), .B(n_1231), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1283), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1261), .B(n_1231), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1301), .B(n_1259), .Y(n_1334) );
XOR2x2_ASAP7_75t_L g1335 ( .A(n_1292), .B(n_1184), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1302), .Y(n_1336) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_1310), .A2(n_1298), .B1(n_1291), .B2(n_1236), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1304), .Y(n_1338) );
NOR2xp33_ASAP7_75t_L g1339 ( .A(n_1317), .B(n_1299), .Y(n_1339) );
XNOR2xp5_ASAP7_75t_L g1340 ( .A(n_1335), .B(n_1086), .Y(n_1340) );
OAI21xp33_ASAP7_75t_L g1341 ( .A1(n_1320), .A2(n_1264), .B(n_1262), .Y(n_1341) );
INVx1_ASAP7_75t_SL g1342 ( .A(n_1335), .Y(n_1342) );
AO22x2_ASAP7_75t_L g1343 ( .A1(n_1322), .A2(n_1292), .B1(n_1255), .B2(n_1258), .Y(n_1343) );
CKINVDCx14_ASAP7_75t_R g1344 ( .A(n_1319), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1304), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1316), .B(n_1279), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1334), .B(n_1253), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1306), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1306), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1315), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1321), .B(n_1286), .Y(n_1351) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_1305), .B(n_1295), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1315), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1325), .B(n_1253), .Y(n_1354) );
OAI21xp33_ASAP7_75t_L g1355 ( .A1(n_1318), .A2(n_1264), .B(n_1262), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_1324), .A2(n_1231), .B1(n_1236), .B2(n_1249), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1307), .B(n_1287), .Y(n_1357) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1329), .Y(n_1358) );
AOI222xp33_ASAP7_75t_L g1359 ( .A1(n_1324), .A2(n_1272), .B1(n_1269), .B2(n_1313), .C1(n_1309), .C2(n_1229), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_1324), .A2(n_1236), .B1(n_1249), .B2(n_1199), .Y(n_1360) );
OAI211xp5_ASAP7_75t_L g1361 ( .A1(n_1342), .A2(n_1142), .B(n_1093), .C(n_1300), .Y(n_1361) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_1344), .B(n_1314), .Y(n_1362) );
NAND2xp33_ASAP7_75t_SL g1363 ( .A(n_1340), .B(n_1305), .Y(n_1363) );
OAI21xp5_ASAP7_75t_SL g1364 ( .A1(n_1356), .A2(n_1257), .B(n_1183), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1352), .Y(n_1365) );
INVx2_ASAP7_75t_SL g1366 ( .A(n_1343), .Y(n_1366) );
XNOR2x1_ASAP7_75t_L g1367 ( .A(n_1343), .B(n_1327), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1338), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1345), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1348), .Y(n_1370) );
AOI221xp5_ASAP7_75t_L g1371 ( .A1(n_1341), .A2(n_1303), .B1(n_1308), .B2(n_1326), .C(n_1318), .Y(n_1371) );
OAI211xp5_ASAP7_75t_L g1372 ( .A1(n_1337), .A2(n_1229), .B(n_1327), .C(n_1215), .Y(n_1372) );
NAND2xp5_ASAP7_75t_SL g1373 ( .A(n_1359), .B(n_1323), .Y(n_1373) );
AOI211xp5_ASAP7_75t_L g1374 ( .A1(n_1339), .A2(n_1291), .B(n_1248), .C(n_1236), .Y(n_1374) );
AOI21xp33_ASAP7_75t_L g1375 ( .A1(n_1343), .A2(n_1112), .B(n_1251), .Y(n_1375) );
NOR2xp33_ASAP7_75t_L g1376 ( .A(n_1357), .B(n_1331), .Y(n_1376) );
OAI221xp5_ASAP7_75t_SL g1377 ( .A1(n_1364), .A2(n_1360), .B1(n_1355), .B2(n_1282), .C(n_1346), .Y(n_1377) );
AOI211xp5_ASAP7_75t_L g1378 ( .A1(n_1361), .A2(n_1251), .B(n_1291), .C(n_1236), .Y(n_1378) );
NAND3xp33_ASAP7_75t_L g1379 ( .A(n_1366), .B(n_1349), .C(n_1350), .Y(n_1379) );
AOI222xp33_ASAP7_75t_L g1380 ( .A1(n_1363), .A2(n_1353), .B1(n_1351), .B2(n_1347), .C1(n_1354), .C2(n_1308), .Y(n_1380) );
A2O1A1Ixp33_ASAP7_75t_L g1381 ( .A1(n_1362), .A2(n_1323), .B(n_1333), .C(n_1331), .Y(n_1381) );
NAND3xp33_ASAP7_75t_L g1382 ( .A(n_1367), .B(n_1330), .C(n_1328), .Y(n_1382) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_1373), .A2(n_1347), .B1(n_1354), .B2(n_1303), .C(n_1336), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_1371), .A2(n_1249), .B1(n_1282), .B2(n_1199), .Y(n_1384) );
NAND2xp33_ASAP7_75t_R g1385 ( .A(n_1362), .B(n_1282), .Y(n_1385) );
INVxp67_ASAP7_75t_L g1386 ( .A(n_1376), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1365), .B(n_1311), .Y(n_1387) );
AOI21xp33_ASAP7_75t_L g1388 ( .A1(n_1385), .A2(n_1372), .B(n_1375), .Y(n_1388) );
NAND5xp2_ASAP7_75t_L g1389 ( .A(n_1377), .B(n_1374), .C(n_1376), .D(n_1215), .E(n_1141), .Y(n_1389) );
OAI211xp5_ASAP7_75t_L g1390 ( .A1(n_1380), .A2(n_1112), .B(n_1369), .C(n_1368), .Y(n_1390) );
OAI221xp5_ASAP7_75t_L g1391 ( .A1(n_1382), .A2(n_1370), .B1(n_1358), .B2(n_1336), .C(n_1332), .Y(n_1391) );
AND2x4_ASAP7_75t_L g1392 ( .A(n_1386), .B(n_1333), .Y(n_1392) );
AOI311xp33_ASAP7_75t_L g1393 ( .A1(n_1383), .A2(n_1332), .A3(n_1330), .B(n_1328), .C(n_1288), .Y(n_1393) );
NOR2x1_ASAP7_75t_L g1394 ( .A(n_1379), .B(n_1312), .Y(n_1394) );
NOR4xp25_ASAP7_75t_L g1395 ( .A(n_1384), .B(n_1312), .C(n_1154), .D(n_1311), .Y(n_1395) );
NAND3xp33_ASAP7_75t_SL g1396 ( .A(n_1390), .B(n_1378), .C(n_1381), .Y(n_1396) );
AND3x4_ASAP7_75t_L g1397 ( .A(n_1395), .B(n_1394), .C(n_1392), .Y(n_1397) );
AND2x4_ASAP7_75t_L g1398 ( .A(n_1392), .B(n_1387), .Y(n_1398) );
AND5x1_ASAP7_75t_L g1399 ( .A(n_1389), .B(n_1206), .C(n_1220), .D(n_1232), .E(n_1251), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1388), .B(n_1249), .Y(n_1400) );
XNOR2xp5_ASAP7_75t_L g1401 ( .A(n_1391), .B(n_1232), .Y(n_1401) );
INVx3_ASAP7_75t_L g1402 ( .A(n_1398), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1400), .Y(n_1403) );
AOI221xp5_ASAP7_75t_L g1404 ( .A1(n_1396), .A2(n_1393), .B1(n_1228), .B2(n_1241), .C(n_1253), .Y(n_1404) );
OAI22xp5_ASAP7_75t_SL g1405 ( .A1(n_1397), .A2(n_1232), .B1(n_1222), .B2(n_1228), .Y(n_1405) );
OA22x2_ASAP7_75t_L g1406 ( .A1(n_1402), .A2(n_1401), .B1(n_1399), .B2(n_1190), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1403), .Y(n_1407) );
OR2x2_ASAP7_75t_L g1408 ( .A(n_1405), .B(n_1401), .Y(n_1408) );
XNOR2x1_ASAP7_75t_L g1409 ( .A(n_1404), .B(n_1114), .Y(n_1409) );
NOR3xp33_ASAP7_75t_L g1410 ( .A(n_1407), .B(n_1128), .C(n_1154), .Y(n_1410) );
OAI22xp5_ASAP7_75t_SL g1411 ( .A1(n_1408), .A2(n_1232), .B1(n_1222), .B2(n_1149), .Y(n_1411) );
AOI22x1_ASAP7_75t_L g1412 ( .A1(n_1406), .A2(n_1101), .B1(n_1105), .B2(n_1118), .Y(n_1412) );
OAI21xp5_ASAP7_75t_L g1413 ( .A1(n_1412), .A2(n_1409), .B(n_1410), .Y(n_1413) );
OAI21xp5_ASAP7_75t_SL g1414 ( .A1(n_1411), .A2(n_1114), .B(n_1118), .Y(n_1414) );
AO221x1_ASAP7_75t_L g1415 ( .A1(n_1411), .A2(n_1241), .B1(n_1195), .B2(n_1168), .C(n_1128), .Y(n_1415) );
AOI21xp5_ASAP7_75t_L g1416 ( .A1(n_1413), .A2(n_1415), .B(n_1414), .Y(n_1416) );
OAI21xp5_ASAP7_75t_L g1417 ( .A1(n_1416), .A2(n_1108), .B(n_1145), .Y(n_1417) );
AOI22xp33_ASAP7_75t_SL g1418 ( .A1(n_1417), .A2(n_1222), .B1(n_1190), .B2(n_1196), .Y(n_1418) );
endmodule