module fake_ariane_2615_n_4638 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_913, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_878, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_850, n_908, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_906, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_864, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_897, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_891, n_737, n_137, n_885, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_870, n_87, n_714, n_279, n_905, n_702, n_207, n_790, n_857, n_898, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_900, n_154, n_883, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_871, n_315, n_903, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_879, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_855, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_858, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_901, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_894, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_868, n_326, n_681, n_778, n_227, n_48, n_874, n_188, n_323, n_550, n_635, n_707, n_330, n_914, n_400, n_689, n_694, n_884, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_859, n_636, n_427, n_108, n_587, n_497, n_693, n_863, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_899, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_887, n_661, n_488, n_775, n_667, n_300, n_533, n_904, n_505, n_14, n_163, n_88, n_869, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_889, n_579, n_844, n_459, n_685, n_221, n_321, n_911, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_861, n_175, n_711, n_877, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_907, n_235, n_881, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_910, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_371, n_845, n_888, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_865, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_860, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_851, n_255, n_560, n_450, n_890, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_896, n_409, n_171, n_519, n_902, n_384, n_468, n_853, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_872, n_13, n_27, n_254, n_596, n_912, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_915, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_862, n_110, n_304, n_895, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_875, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_880, n_793, n_852, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_873, n_51, n_496, n_739, n_76, n_342, n_866, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_892, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_882, n_317, n_867, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_856, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_876, n_618, n_411, n_484, n_712, n_849, n_909, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_893, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_854, n_471, n_351, n_886, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_4638);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_913;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_878;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_850;
input n_908;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_906;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_864;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_897;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_891;
input n_737;
input n_137;
input n_885;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_870;
input n_87;
input n_714;
input n_279;
input n_905;
input n_702;
input n_207;
input n_790;
input n_857;
input n_898;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_900;
input n_154;
input n_883;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_871;
input n_315;
input n_903;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_879;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_855;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_858;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_901;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_894;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_868;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_874;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_914;
input n_400;
input n_689;
input n_694;
input n_884;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_859;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_863;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_899;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_887;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_904;
input n_505;
input n_14;
input n_163;
input n_88;
input n_869;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_889;
input n_579;
input n_844;
input n_459;
input n_685;
input n_221;
input n_321;
input n_911;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_861;
input n_175;
input n_711;
input n_877;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_907;
input n_235;
input n_881;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_910;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_371;
input n_845;
input n_888;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_865;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_860;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_851;
input n_255;
input n_560;
input n_450;
input n_890;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_896;
input n_409;
input n_171;
input n_519;
input n_902;
input n_384;
input n_468;
input n_853;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_872;
input n_13;
input n_27;
input n_254;
input n_596;
input n_912;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_915;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_862;
input n_110;
input n_304;
input n_895;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_875;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_880;
input n_793;
input n_852;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_873;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_866;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_892;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_882;
input n_317;
input n_867;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_856;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_876;
input n_618;
input n_411;
input n_484;
input n_712;
input n_849;
input n_909;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_893;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_854;
input n_471;
input n_351;
input n_886;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_4638;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_4030;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_4586;
wire n_1469;
wire n_4342;
wire n_4557;
wire n_3056;
wire n_1353;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_4382;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_4259;
wire n_3264;
wire n_4475;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_3181;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_4403;
wire n_4602;
wire n_1713;
wire n_2818;
wire n_1436;
wire n_2407;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_1430;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_4626;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_1837;
wire n_924;
wire n_4178;
wire n_2013;
wire n_2786;
wire n_4547;
wire n_1566;
wire n_2837;
wire n_3765;
wire n_2006;
wire n_4058;
wire n_952;
wire n_4090;
wire n_2446;
wire n_1096;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_2461;
wire n_2207;
wire n_2702;
wire n_1706;
wire n_3719;
wire n_4363;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_3954;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_4103;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_4610;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_2278;
wire n_4028;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_4416;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4439;
wire n_2547;
wire n_4600;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_4575;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_4106;
wire n_4589;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_4581;
wire n_2960;
wire n_4260;
wire n_4625;
wire n_3270;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_4148;
wire n_1062;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_4512;
wire n_2342;
wire n_4590;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_4132;
wire n_4038;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_953;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_4500;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_2634;
wire n_3451;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_4515;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_2878;
wire n_1284;
wire n_1428;
wire n_1241;
wire n_3890;
wire n_3830;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_2782;
wire n_4136;
wire n_4604;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_4353;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_4567;
wire n_4176;
wire n_1207;
wire n_4124;
wire n_3606;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_3474;
wire n_2232;
wire n_4488;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_3552;
wire n_1542;
wire n_3756;
wire n_1314;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_1512;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_3412;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_4608;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_4597;
wire n_4560;
wire n_3482;
wire n_1900;
wire n_3948;
wire n_4621;
wire n_1074;
wire n_3230;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_4546;
wire n_1889;
wire n_1977;
wire n_2650;
wire n_1254;
wire n_3960;
wire n_4454;
wire n_4147;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_2332;
wire n_1703;
wire n_2391;
wire n_3828;
wire n_3975;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_4018;
wire n_4576;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_3003;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1560;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_4572;
wire n_4505;
wire n_2575;
wire n_2722;
wire n_3728;
wire n_3739;
wire n_1840;
wire n_1230;
wire n_2739;
wire n_1396;
wire n_3962;
wire n_1597;
wire n_4082;
wire n_4476;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_4541;
wire n_4360;
wire n_1544;
wire n_3271;
wire n_4540;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1790;
wire n_1354;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_4443;
wire n_1021;
wire n_1443;
wire n_4000;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_3458;
wire n_2727;
wire n_4593;
wire n_942;
wire n_4562;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_2909;
wire n_1378;
wire n_1121;
wire n_3554;
wire n_1416;
wire n_1461;
wire n_3012;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3850;
wire n_4529;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_4498;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_4432;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_4495;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_4357;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_4109;
wire n_3777;
wire n_4108;
wire n_4502;
wire n_4530;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_3588;
wire n_1108;
wire n_3692;
wire n_1590;
wire n_3280;
wire n_3234;
wire n_3413;
wire n_3900;
wire n_1351;
wire n_4115;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_4394;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_930;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_4513;
wire n_1179;
wire n_4311;
wire n_3284;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_2810;
wire n_1386;
wire n_3391;
wire n_3506;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_1253;
wire n_2791;
wire n_1468;
wire n_1661;
wire n_4378;
wire n_2683;
wire n_3212;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_4354;
wire n_4405;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_4459;
wire n_992;
wire n_966;
wire n_955;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_4594;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_4345;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_2398;
wire n_4233;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_1972;
wire n_1178;
wire n_2015;
wire n_2925;
wire n_1292;
wire n_3717;
wire n_3407;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_4029;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2930;
wire n_2871;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_1491;
wire n_931;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_967;
wire n_1083;
wire n_3937;
wire n_4130;
wire n_2161;
wire n_1418;
wire n_4175;
wire n_1357;
wire n_1079;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_4587;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_4456;
wire n_1312;
wire n_4508;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_1812;
wire n_3651;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_2224;
wire n_1226;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_3046;
wire n_2668;
wire n_2921;
wire n_1240;
wire n_1087;
wire n_4055;
wire n_3980;
wire n_4410;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_3741;
wire n_2388;
wire n_4352;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_976;
wire n_3567;
wire n_4003;
wire n_1832;
wire n_2795;
wire n_1392;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_4438;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_3884;
wire n_1731;
wire n_4433;
wire n_2829;
wire n_1147;
wire n_4367;
wire n_4492;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_965;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_3010;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_4445;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_4254;
wire n_4462;
wire n_2507;
wire n_4219;
wire n_4484;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_4043;
wire n_4336;
wire n_4451;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1234;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_3981;
wire n_1247;
wire n_4234;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_1255;
wire n_2632;
wire n_3179;
wire n_3031;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_4613;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_927;
wire n_2980;
wire n_1095;
wire n_3699;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3971;
wire n_4315;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_4442;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_4494;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_4201;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_2312;
wire n_2677;
wire n_4296;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_2812;
wire n_3660;
wire n_1592;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_4386;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_4049;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_4522;
wire n_2718;
wire n_4263;
wire n_926;
wire n_1943;
wire n_2687;
wire n_4426;
wire n_2296;
wire n_3876;
wire n_4588;
wire n_3615;
wire n_4362;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_3946;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_2640;
wire n_1163;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_4634;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4089;
wire n_1501;
wire n_4186;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3513;
wire n_3498;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_1198;
wire n_4096;
wire n_4506;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_1879;
wire n_1886;
wire n_4346;
wire n_4138;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_3968;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_2122;
wire n_3572;
wire n_1611;
wire n_2975;
wire n_3332;
wire n_4337;
wire n_2399;
wire n_4543;
wire n_1414;
wire n_2067;
wire n_1134;
wire n_3374;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_4555;
wire n_1901;
wire n_2055;
wire n_4486;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_4359;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_4072;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4441;
wire n_1906;
wire n_4323;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_3922;
wire n_4447;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_1467;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_4458;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_4523;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_3705;
wire n_3983;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3286;
wire n_4480;
wire n_3734;
wire n_3370;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_4583;
wire n_3788;
wire n_3939;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_3569;
wire n_2523;
wire n_1945;
wire n_3542;
wire n_3835;
wire n_3837;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_2496;
wire n_1162;
wire n_2031;
wire n_3260;
wire n_1614;
wire n_3349;
wire n_3761;
wire n_3819;
wire n_3996;
wire n_4292;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_4348;
wire n_4616;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_4374;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_3403;
wire n_4261;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4344;
wire n_4084;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_957;
wire n_1402;
wire n_1242;
wire n_3957;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_4580;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_4393;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_1431;
wire n_4389;
wire n_3995;
wire n_1119;
wire n_4460;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_4481;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4461;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_4615;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3501;
wire n_3492;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_3931;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2949;
wire n_2661;
wire n_1667;
wire n_2894;
wire n_2300;
wire n_3896;
wire n_4067;
wire n_2452;
wire n_1649;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_4551;
wire n_3214;
wire n_3551;
wire n_4521;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_4525;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1219;
wire n_1711;
wire n_4387;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_4369;
wire n_2124;
wire n_1894;
wire n_2594;
wire n_1239;
wire n_1460;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_4324;
wire n_3626;
wire n_1898;
wire n_4428;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_4598;
wire n_4464;
wire n_4463;
wire n_1793;
wire n_4446;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1975;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_2119;
wire n_1719;
wire n_2742;
wire n_1540;
wire n_3671;
wire n_4396;
wire n_4440;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_4425;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_4565;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_3065;
wire n_3016;
wire n_4114;
wire n_2460;
wire n_4552;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_4482;
wire n_2480;
wire n_951;
wire n_3024;
wire n_4528;
wire n_2772;
wire n_3564;
wire n_1700;
wire n_2637;
wire n_3795;
wire n_1332;
wire n_2306;
wire n_4328;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_3990;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_4400;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4568;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2916;
wire n_3617;
wire n_2576;
wire n_3459;
wire n_1394;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_4351;
wire n_4424;
wire n_3340;
wire n_4429;
wire n_4192;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_2468;
wire n_2171;
wire n_1243;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1527;
wire n_2581;
wire n_1513;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_4524;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_4436;
wire n_3197;
wire n_1993;
wire n_3586;
wire n_1545;
wire n_2629;
wire n_3369;
wire n_4035;
wire n_4160;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_4190;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_4545;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_4145;
wire n_3097;
wire n_4395;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_2492;
wire n_3864;
wire n_4385;
wire n_2939;
wire n_3425;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_4633;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_4050;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_4306;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_4558;
wire n_1318;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_4511;
wire n_4358;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1281;
wire n_4289;
wire n_1873;
wire n_1137;
wire n_1856;
wire n_1476;
wire n_2723;
wire n_1733;
wire n_1258;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_1524;
wire n_3925;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_2850;
wire n_1874;
wire n_3167;
wire n_1293;
wire n_3746;
wire n_961;
wire n_4537;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_4618;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3753;
wire n_3893;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_4076;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_2720;
wire n_1556;
wire n_2412;
wire n_1561;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_2064;
wire n_2353;
wire n_1429;
wire n_3543;
wire n_2528;
wire n_1778;
wire n_3640;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_1154;
wire n_3609;
wire n_1759;
wire n_1557;
wire n_1829;
wire n_2325;
wire n_4330;
wire n_1130;
wire n_4635;
wire n_1450;
wire n_4152;
wire n_3718;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_3879;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_4343;
wire n_2298;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2570;
wire n_2329;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_2546;
wire n_949;
wire n_2454;
wire n_2911;
wire n_2890;
wire n_3455;
wire n_3381;
wire n_1493;
wire n_3736;
wire n_4466;
wire n_3313;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3907;
wire n_4603;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_4419;
wire n_1151;
wire n_4595;
wire n_960;
wire n_4420;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_3605;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4404;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_4630;
wire n_4372;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_4377;
wire n_4617;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_4563;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4301;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_4561;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_3654;
wire n_4188;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_4399;
wire n_2413;
wire n_4008;
wire n_2610;
wire n_1593;
wire n_3715;
wire n_4140;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_2605;
wire n_1201;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_3982;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_2665;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_3973;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_3842;
wire n_4202;
wire n_4536;
wire n_2044;
wire n_4534;
wire n_928;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_3769;
wire n_4078;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_4437;
wire n_1192;
wire n_3738;
wire n_3098;
wire n_1380;
wire n_4503;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_4070;
wire n_2020;
wire n_3987;
wire n_2310;
wire n_4249;
wire n_4418;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_4139;
wire n_4582;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_4450;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_3967;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_1517;
wire n_2036;
wire n_4412;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_4368;
wire n_3444;
wire n_4370;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_4091;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_4184;
wire n_4430;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_4631;
wire n_2234;
wire n_1341;
wire n_1356;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1955;
wire n_1504;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_4538;
wire n_4544;
wire n_1370;
wire n_1603;
wire n_4191;
wire n_4478;
wire n_4409;
wire n_2935;
wire n_2401;
wire n_4246;
wire n_3822;
wire n_3255;
wire n_3818;
wire n_1549;
wire n_1066;
wire n_4355;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_4061;
wire n_2658;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_4601;
wire n_3344;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_4518;
wire n_4155;
wire n_3376;
wire n_4278;
wire n_4531;
wire n_1290;
wire n_1959;
wire n_3770;
wire n_3497;
wire n_4375;
wire n_4542;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_2121;
wire n_1559;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_4532;
wire n_2692;
wire n_3927;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_2553;
wire n_2645;
wire n_1420;
wire n_3790;
wire n_2749;
wire n_2592;
wire n_1454;
wire n_3490;
wire n_2459;
wire n_962;
wire n_4413;
wire n_941;
wire n_3396;
wire n_1210;
wire n_4241;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_3288;
wire n_3251;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_4341;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3904;
wire n_3887;
wire n_3195;
wire n_3008;
wire n_3242;
wire n_1695;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_4126;
wire n_4164;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_3836;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_3409;
wire n_1653;
wire n_1749;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4381;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_4469;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_4455;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_4384;
wire n_1584;
wire n_1157;
wire n_4366;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_1814;
wire n_4210;
wire n_4577;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_4208;
wire n_3972;
wire n_2054;
wire n_4623;
wire n_1857;
wire n_2315;
wire n_3926;
wire n_4209;
wire n_984;
wire n_1687;
wire n_4457;
wire n_2073;
wire n_2150;
wire n_4509;
wire n_4004;
wire n_1552;
wire n_2938;
wire n_3630;
wire n_2498;
wire n_1612;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_4350;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2602;
wire n_2444;
wire n_3354;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_3106;
wire n_2977;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_1100;
wire n_2455;
wire n_1617;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_2828;
wire n_4212;
wire n_4270;
wire n_1626;
wire n_3436;
wire n_4620;
wire n_4584;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_3751;
wire n_2299;
wire n_4388;
wire n_3402;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_4477;
wire n_1621;
wire n_4110;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_4411;
wire n_1221;
wire n_4217;
wire n_4585;
wire n_1785;
wire n_1262;
wire n_4271;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_4317;
wire n_4406;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_4605;
wire n_3301;
wire n_981;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_2503;
wire n_3873;
wire n_1758;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_2465;
wire n_3610;
wire n_1407;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_3100;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_4592;
wire n_1176;
wire n_3721;
wire n_3676;
wire n_1564;
wire n_2010;
wire n_3677;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_2356;
wire n_1361;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_1057;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_2941;
wire n_1509;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_3536;
wire n_2564;
wire n_1721;
wire n_3558;
wire n_3576;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_3034;
wire n_1317;
wire n_1445;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_4435;
wire n_4053;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_3091;
wire n_1024;
wire n_4496;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_4596;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_4628;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_4554;
wire n_2630;
wire n_4105;
wire n_4526;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_3114;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_3225;
wire n_2086;
wire n_1625;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_4578;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_2409;
wire n_2966;
wire n_1720;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_3360;
wire n_4470;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_1809;
wire n_2787;
wire n_4092;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_2215;
wire n_1530;
wire n_4057;
wire n_2770;
wire n_4550;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_4347;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3633;
wire n_3042;
wire n_1067;
wire n_968;
wire n_4144;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_4379;
wire n_3111;
wire n_2212;
wire n_3838;
wire n_1813;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_2268;
wire n_4434;
wire n_2835;
wire n_1452;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_4499;
wire n_2569;
wire n_4504;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_4339;
wire n_1322;
wire n_3273;
wire n_4497;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_4510;
wire n_3155;
wire n_4300;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4472;
wire n_4253;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_1710;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_2580;
wire n_2699;
wire n_1390;
wire n_1792;
wire n_4064;
wire n_3351;
wire n_2062;
wire n_4489;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_2153;
wire n_2324;
wire n_1459;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_4519;
wire n_1099;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_4197;
wire n_4564;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_3776;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_4566;
wire n_3970;
wire n_4371;
wire n_1619;
wire n_2351;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_4080;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_3898;
wire n_4414;
wire n_2541;
wire n_1643;
wire n_4185;
wire n_3188;
wire n_3232;
wire n_3001;
wire n_1320;
wire n_4448;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_2447;
wire n_4295;
wire n_3932;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_4579;
wire n_4507;
wire n_2104;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_2552;
wire n_1806;
wire n_3445;
wire n_1576;
wire n_1533;
wire n_1470;
wire n_4087;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_4473;
wire n_4619;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_4398;
wire n_3253;
wire n_4471;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_4392;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_4238;
wire n_4365;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_4349;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3966;
wire n_4397;
wire n_4449;
wire n_3285;
wire n_3824;
wire n_4607;
wire n_3825;
wire n_4198;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_1150;
wire n_4266;
wire n_977;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_3874;
wire n_4373;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_4407;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_4165;
wire n_4154;
wire n_4479;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_4390;
wire n_3845;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_3941;
wire n_1915;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_2240;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_2846;
wire n_4258;
wire n_3371;
wire n_1781;
wire n_4571;
wire n_2917;
wire n_3137;
wire n_4250;
wire n_2544;
wire n_3194;
wire n_3143;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_4415;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1477;
wire n_2097;
wire n_1982;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_939;
wire n_1410;
wire n_2297;
wire n_4276;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2957;
wire n_4408;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_4569;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_4483;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_4128;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_4036;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_4487;
wire n_4548;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_4539;
wire n_4574;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_3071;
wire n_3918;
wire n_4010;
wire n_4329;
wire n_1571;
wire n_4501;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_1946;
wire n_2148;
wire n_933;
wire n_3244;
wire n_4383;
wire n_3499;
wire n_4391;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1821;
wire n_1168;
wire n_4095;
wire n_4444;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3910;
wire n_3947;
wire n_4485;
wire n_4624;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_2585;
wire n_1591;
wire n_3293;
wire n_2995;
wire n_3361;
wire n_4287;
wire n_4533;
wire n_1229;
wire n_2582;
wire n_1683;
wire n_3228;
wire n_3327;
wire n_4356;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_2381;
wire n_1732;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_3707;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3779;
wire n_3895;
wire n_4627;
wire n_3149;
wire n_1063;
wire n_3934;
wire n_4556;
wire n_2205;
wire n_991;
wire n_2183;
wire n_2275;
wire n_4338;
wire n_2563;
wire n_3088;
wire n_1724;
wire n_4224;
wire n_4606;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_4573;
wire n_938;
wire n_1891;
wire n_4520;
wire n_1328;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_4042;
wire n_1581;
wire n_3849;
wire n_4244;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_2792;
wire n_1818;
wire n_1146;
wire n_3398;
wire n_3709;
wire n_1655;
wire n_4465;
wire n_4553;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_3557;
wire n_3592;
wire n_3725;
wire n_1598;
wire n_3986;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_3399;
wire n_3894;
wire n_1702;
wire n_4612;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1368;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_2891;
wire n_1725;
wire n_4335;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_4120;
wire n_4149;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_2361;
wire n_2819;
wire n_1115;
wire n_2229;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_1722;
wire n_3505;
wire n_4277;
wire n_1339;
wire n_4614;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_4629;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_4516;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_4599;
wire n_1010;
wire n_2830;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4622;
wire n_4222;
wire n_1871;
wire n_2514;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_3162;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_4591;
wire n_4046;
wire n_4467;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_4570;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_3041;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_4493;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_4376;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_2479;
wire n_3204;
wire n_1981;
wire n_1069;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_2345;
wire n_4417;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_457),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_456),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_5),
.Y(n_918)
);

BUFx10_ASAP7_75t_L g919 ( 
.A(n_279),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_186),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_631),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_272),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_336),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_894),
.Y(n_924)
);

BUFx10_ASAP7_75t_L g925 ( 
.A(n_534),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_852),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_795),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_459),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_93),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_624),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_682),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_791),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_310),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_864),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_74),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_691),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_273),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_611),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_9),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_898),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_126),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_142),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_354),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_849),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_767),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_629),
.Y(n_946)
);

INVx4_ASAP7_75t_R g947 ( 
.A(n_173),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_197),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_911),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_889),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_271),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_193),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_405),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_428),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_216),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_14),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_328),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_583),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_674),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_391),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_664),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_526),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_692),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_536),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_819),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_26),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_776),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_551),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_145),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_578),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_618),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_559),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_905),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_324),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_645),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_144),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_245),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_718),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_732),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_895),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_737),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_582),
.Y(n_982)
);

CKINVDCx11_ASAP7_75t_R g983 ( 
.A(n_681),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_37),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_803),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_736),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_263),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_676),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_666),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_503),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_427),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_638),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_284),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_588),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_486),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_541),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_591),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_641),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_466),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_476),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_302),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_415),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_822),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_568),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_743),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_106),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_346),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_476),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_283),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_670),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_443),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_274),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_233),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_815),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_883),
.Y(n_1015)
);

BUFx10_ASAP7_75t_L g1016 ( 
.A(n_205),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_237),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_366),
.Y(n_1018)
);

BUFx5_ASAP7_75t_L g1019 ( 
.A(n_521),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_751),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_299),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_711),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_338),
.Y(n_1023)
);

CKINVDCx14_ASAP7_75t_R g1024 ( 
.A(n_580),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_809),
.Y(n_1025)
);

BUFx10_ASAP7_75t_L g1026 ( 
.A(n_148),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_760),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_414),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_596),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_411),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_608),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_108),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_772),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_80),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_231),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_359),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_203),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_559),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_865),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_548),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_431),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_775),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_147),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_611),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_716),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_234),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_613),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_91),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_709),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_915),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_594),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_812),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_783),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_51),
.Y(n_1054)
);

BUFx5_ASAP7_75t_L g1055 ( 
.A(n_610),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_899),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_584),
.Y(n_1057)
);

BUFx10_ASAP7_75t_L g1058 ( 
.A(n_185),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_661),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_602),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_432),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_687),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_587),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_123),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_543),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_167),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_480),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_482),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_461),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_487),
.Y(n_1070)
);

CKINVDCx16_ASAP7_75t_R g1071 ( 
.A(n_486),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_519),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_801),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_222),
.Y(n_1074)
);

CKINVDCx16_ASAP7_75t_R g1075 ( 
.A(n_738),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_296),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_411),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_781),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_495),
.Y(n_1079)
);

CKINVDCx16_ASAP7_75t_R g1080 ( 
.A(n_373),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_335),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_734),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_712),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_412),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_722),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_818),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_546),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_256),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_552),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_621),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_527),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_490),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_42),
.Y(n_1093)
);

CKINVDCx16_ASAP7_75t_R g1094 ( 
.A(n_374),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_229),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_805),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_38),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_572),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_368),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_829),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_503),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_846),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_143),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_90),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_636),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_806),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_620),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_786),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_828),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_221),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_168),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_823),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_106),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_374),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_679),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_678),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_804),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_813),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_845),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_109),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_686),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_256),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_348),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_325),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_442),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_886),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_459),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_598),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_265),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_669),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_847),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_887),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_549),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_604),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_12),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_667),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_518),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_824),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_280),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_485),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_780),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_639),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_825),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_586),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_211),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_560),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_875),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_416),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_842),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_113),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_499),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_157),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_321),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_409),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_579),
.Y(n_1155)
);

BUFx10_ASAP7_75t_L g1156 ( 
.A(n_884),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_409),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_491),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_556),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_876),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_210),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_575),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_295),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_294),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_381),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_533),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_92),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_689),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_564),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_267),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_402),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_719),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_117),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_644),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_793),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_222),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_135),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_128),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_904),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_826),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_909),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_902),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_800),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_52),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_448),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_34),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_66),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_164),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_58),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_696),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_632),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_817),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_603),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_656),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_389),
.Y(n_1195)
);

BUFx8_ASAP7_75t_SL g1196 ( 
.A(n_51),
.Y(n_1196)
);

CKINVDCx16_ASAP7_75t_R g1197 ( 
.A(n_702),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_159),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_890),
.Y(n_1199)
);

INVxp67_ASAP7_75t_SL g1200 ( 
.A(n_382),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_385),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_548),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_555),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_537),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_545),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_480),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_810),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_489),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_833),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_285),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_768),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_201),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_893),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_605),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_592),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_386),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_148),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_727),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_649),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_272),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_184),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_196),
.Y(n_1222)
);

CKINVDCx14_ASAP7_75t_R g1223 ( 
.A(n_349),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_705),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_658),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_605),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_107),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_156),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_769),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_519),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_361),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_477),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_455),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_483),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_394),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_537),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_200),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_376),
.Y(n_1238)
);

CKINVDCx14_ASAP7_75t_R g1239 ( 
.A(n_617),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_530),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_642),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_27),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_814),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_619),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_197),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_421),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_700),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_699),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_502),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_758),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_797),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_654),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_342),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_445),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_173),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_579),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_471),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_44),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_129),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_520),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_610),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_139),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_311),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_126),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_592),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_901),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_891),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_713),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_167),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_693),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_526),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_301),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_855),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_39),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_478),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_609),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_216),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_187),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_908),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_860),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_426),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_697),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_569),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_282),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_209),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_623),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_417),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_637),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_488),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_133),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_146),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_176),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_594),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_34),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_532),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_892),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_862),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_332),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_897),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_291),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_635),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_164),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_47),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_573),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_245),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_888),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_774),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_640),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_315),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_715),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_668),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_460),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_102),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_914),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_602),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_749),
.Y(n_1316)
);

BUFx8_ASAP7_75t_SL g1317 ( 
.A(n_266),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_146),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_501),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_753),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_96),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_785),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_488),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_869),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_255),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_741),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_159),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_569),
.Y(n_1328)
);

BUFx10_ASAP7_75t_L g1329 ( 
.A(n_646),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_740),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_683),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_773),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_294),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_790),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_787),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_840),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_777),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_94),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_209),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_680),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_832),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_26),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_504),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_183),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_744),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_622),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_58),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_651),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_770),
.Y(n_1349)
);

INVxp33_ASAP7_75t_SL g1350 ( 
.A(n_484),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_730),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_778),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_119),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_188),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_866),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_528),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_399),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_903),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_746),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_235),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_728),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_614),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_432),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_574),
.Y(n_1364)
);

BUFx10_ASAP7_75t_L g1365 ( 
.A(n_858),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_80),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_870),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_220),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_37),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_421),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_75),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_566),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_85),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_405),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_83),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_342),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_428),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_671),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_648),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_871),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_839),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_485),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_95),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_584),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_600),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_684),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_392),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_707),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_354),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_708),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_657),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_550),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_567),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_688),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_325),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_851),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_907),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_867),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_81),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_529),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_874),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_607),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_276),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_565),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_514),
.Y(n_1405)
);

BUFx5_ASAP7_75t_L g1406 ( 
.A(n_698),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_739),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_853),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_759),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_748),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_137),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_228),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_539),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_19),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_516),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_655),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_54),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_15),
.Y(n_1418)
);

BUFx8_ASAP7_75t_SL g1419 ( 
.A(n_588),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_150),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_44),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_192),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_61),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_162),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_525),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_451),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_238),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_400),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_583),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_357),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_571),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_163),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_558),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_281),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_820),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_531),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_28),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_74),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_284),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_717),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_690),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_473),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_784),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_764),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_122),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_418),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_900),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_585),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_521),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_454),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_333),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_752),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_422),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_761),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_102),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_896),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_872),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_750),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_762),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_576),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_326),
.Y(n_1461)
);

BUFx10_ASAP7_75t_L g1462 ( 
.A(n_913),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_82),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_580),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_113),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_338),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_305),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_504),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_549),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_835),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_130),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_218),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_48),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_157),
.Y(n_1474)
);

BUFx5_ASAP7_75t_L g1475 ( 
.A(n_831),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_779),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_425),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_575),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_124),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_841),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_295),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_742),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_675),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_906),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_19),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_808),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_437),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_378),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_706),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_601),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_789),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_721),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_843),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_230),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_141),
.Y(n_1495)
);

CKINVDCx14_ASAP7_75t_R g1496 ( 
.A(n_633),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_387),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_581),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_838),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_314),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_494),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_375),
.Y(n_1502)
);

CKINVDCx16_ASAP7_75t_R g1503 ( 
.A(n_171),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_512),
.Y(n_1504)
);

BUFx10_ASAP7_75t_L g1505 ( 
.A(n_673),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_628),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_756),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_391),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_547),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_379),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_520),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_393),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_880),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_227),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_912),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_827),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_910),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_418),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_27),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_576),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_10),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_287),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_821),
.Y(n_1523)
);

BUFx10_ASAP7_75t_L g1524 ( 
.A(n_685),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_599),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_878),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_182),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_850),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_369),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_177),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_178),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_16),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_208),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_885),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_86),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_608),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_310),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_652),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_609),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_723),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_299),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_231),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_593),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_442),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_647),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_726),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_703),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_46),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_547),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_448),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_334),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_626),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_771),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_109),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_221),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_399),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_101),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_861),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_517),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_757),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_881),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_392),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_395),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_498),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_293),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_724),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_474),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_280),
.Y(n_1568)
);

CKINVDCx16_ASAP7_75t_R g1569 ( 
.A(n_528),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_794),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_558),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_349),
.Y(n_1572)
);

BUFx10_ASAP7_75t_L g1573 ( 
.A(n_36),
.Y(n_1573)
);

BUFx5_ASAP7_75t_L g1574 ( 
.A(n_440),
.Y(n_1574)
);

BUFx8_ASAP7_75t_SL g1575 ( 
.A(n_115),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_177),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_144),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_97),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_856),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_538),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_731),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_201),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_306),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_788),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_417),
.Y(n_1585)
);

BUFx8_ASAP7_75t_SL g1586 ( 
.A(n_59),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_138),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_190),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_695),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_782),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_515),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_747),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_176),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_363),
.Y(n_1594)
);

BUFx10_ASAP7_75t_L g1595 ( 
.A(n_848),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_799),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_792),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_754),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_258),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_25),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_616),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_606),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_577),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_554),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_165),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_61),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_289),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_242),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_375),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_663),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_653),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_816),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_765),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_535),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_672),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_720),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_561),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_466),
.Y(n_1618)
);

CKINVDCx16_ASAP7_75t_R g1619 ( 
.A(n_598),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_612),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_560),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_114),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_868),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_184),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_271),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_543),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_20),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_328),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_125),
.Y(n_1629)
);

BUFx10_ASAP7_75t_L g1630 ( 
.A(n_21),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_590),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_524),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_830),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_389),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_193),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_304),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_857),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_589),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_811),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_229),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_729),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_701),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_553),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_93),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_477),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_14),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_38),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_677),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_710),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_877),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_599),
.Y(n_1651)
);

BUFx10_ASAP7_75t_L g1652 ( 
.A(n_98),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_83),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_402),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_704),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_151),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_444),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_226),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_542),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_443),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_627),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_562),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_394),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_763),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_66),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_873),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_615),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_286),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_136),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_254),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_334),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_285),
.Y(n_1672)
);

BUFx5_ASAP7_75t_L g1673 ( 
.A(n_807),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_95),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_441),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_802),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_189),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_181),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_834),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_643),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_438),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_694),
.Y(n_1682)
);

BUFx2_ASAP7_75t_SL g1683 ( 
.A(n_650),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_15),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_324),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_603),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_625),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_578),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_597),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_220),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_219),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_269),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_665),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_317),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_725),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_116),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_31),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_379),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_187),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_660),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_401),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_755),
.Y(n_1704)
);

BUFx10_ASAP7_75t_L g1705 ( 
.A(n_563),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_455),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_388),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_530),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_733),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_9),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_662),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_837),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_882),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_863),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_403),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_587),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_156),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_714),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_199),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_798),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_854),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_320),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_879),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_458),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_582),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_395),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_326),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_255),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_254),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_4),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_659),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_451),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_844),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_336),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_544),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_398),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_276),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_423),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_317),
.Y(n_1739)
);

CKINVDCx16_ASAP7_75t_R g1740 ( 
.A(n_297),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_183),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_607),
.Y(n_1742)
);

CKINVDCx20_ASAP7_75t_R g1743 ( 
.A(n_212),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_484),
.Y(n_1744)
);

CKINVDCx20_ASAP7_75t_R g1745 ( 
.A(n_630),
.Y(n_1745)
);

BUFx10_ASAP7_75t_L g1746 ( 
.A(n_571),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_203),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_275),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_570),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_33),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_595),
.Y(n_1751)
);

CKINVDCx16_ASAP7_75t_R g1752 ( 
.A(n_469),
.Y(n_1752)
);

CKINVDCx16_ASAP7_75t_R g1753 ( 
.A(n_796),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_149),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_28),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_836),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_557),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_859),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_502),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_233),
.Y(n_1760)
);

INVxp33_ASAP7_75t_L g1761 ( 
.A(n_735),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_360),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_541),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_766),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_540),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_745),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_634),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_318),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_49),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_957),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1024),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1029),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1029),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1196),
.Y(n_1774)
);

INVxp67_ASAP7_75t_SL g1775 ( 
.A(n_1255),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1255),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_922),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_1024),
.Y(n_1778)
);

INVxp67_ASAP7_75t_SL g1779 ( 
.A(n_922),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1065),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1019),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_962),
.Y(n_1782)
);

INVxp33_ASAP7_75t_L g1783 ( 
.A(n_1317),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1419),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1575),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1019),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_962),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_993),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_993),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1185),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1256),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1185),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1186),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1186),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1257),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1257),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1290),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1290),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1294),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1090),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1019),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1294),
.Y(n_1802)
);

INVxp33_ASAP7_75t_L g1803 ( 
.A(n_1586),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1343),
.Y(n_1804)
);

CKINVDCx16_ASAP7_75t_R g1805 ( 
.A(n_1223),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1343),
.Y(n_1806)
);

INVxp33_ASAP7_75t_L g1807 ( 
.A(n_1467),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1412),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1412),
.Y(n_1809)
);

CKINVDCx20_ASAP7_75t_R g1810 ( 
.A(n_1223),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1439),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1439),
.Y(n_1812)
);

INVxp33_ASAP7_75t_SL g1813 ( 
.A(n_1536),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1549),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1607),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1019),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1549),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1651),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1651),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1675),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_983),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1675),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1717),
.Y(n_1823)
);

CKINVDCx20_ASAP7_75t_R g1824 ( 
.A(n_1039),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1717),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1019),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1019),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1055),
.Y(n_1828)
);

CKINVDCx20_ASAP7_75t_R g1829 ( 
.A(n_1119),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1071),
.Y(n_1830)
);

CKINVDCx16_ASAP7_75t_R g1831 ( 
.A(n_1080),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1055),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1073),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1055),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1055),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1055),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1055),
.Y(n_1837)
);

INVxp67_ASAP7_75t_SL g1838 ( 
.A(n_918),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1678),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1574),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1574),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1574),
.Y(n_1842)
);

CKINVDCx16_ASAP7_75t_R g1843 ( 
.A(n_1094),
.Y(n_1843)
);

INVxp33_ASAP7_75t_L g1844 ( 
.A(n_1004),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1126),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1574),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1574),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_918),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1574),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_918),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_920),
.Y(n_1851)
);

INVxp33_ASAP7_75t_SL g1852 ( 
.A(n_916),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_918),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1350),
.B(n_2),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_941),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_964),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_951),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_952),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_958),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_970),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_974),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_964),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1164),
.Y(n_1863)
);

INVxp67_ASAP7_75t_SL g1864 ( 
.A(n_964),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1338),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_982),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_984),
.Y(n_1867)
);

INVxp33_ASAP7_75t_SL g1868 ( 
.A(n_917),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_995),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_964),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1141),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1006),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1031),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1153),
.Y(n_1874)
);

CKINVDCx16_ASAP7_75t_R g1875 ( 
.A(n_1503),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1034),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1036),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1038),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_938),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_1199),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1054),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1048),
.Y(n_1882)
);

INVxp67_ASAP7_75t_SL g1883 ( 
.A(n_1153),
.Y(n_1883)
);

INVxp67_ASAP7_75t_SL g1884 ( 
.A(n_1153),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1060),
.Y(n_1885)
);

INVxp67_ASAP7_75t_SL g1886 ( 
.A(n_1153),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1569),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1067),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1170),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1068),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1088),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1089),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1219),
.B(n_2),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1091),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1619),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_1213),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1127),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1638),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1128),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1740),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1129),
.Y(n_1901)
);

CKINVDCx20_ASAP7_75t_R g1902 ( 
.A(n_1247),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1135),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1139),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1144),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1145),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1752),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1148),
.Y(n_1908)
);

CKINVDCx20_ASAP7_75t_R g1909 ( 
.A(n_1252),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1151),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1267),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1155),
.Y(n_1912)
);

INVxp33_ASAP7_75t_L g1913 ( 
.A(n_1275),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_969),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1158),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1166),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1299),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1330),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1167),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1359),
.Y(n_1920)
);

CKINVDCx16_ASAP7_75t_R g1921 ( 
.A(n_1049),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1169),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1189),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1278),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_997),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1204),
.Y(n_1926)
);

INVxp67_ASAP7_75t_SL g1927 ( 
.A(n_1189),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1205),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1216),
.Y(n_1929)
);

INVxp67_ASAP7_75t_SL g1930 ( 
.A(n_1189),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1217),
.Y(n_1931)
);

INVxp67_ASAP7_75t_L g1932 ( 
.A(n_1302),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1232),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1233),
.Y(n_1934)
);

INVxp67_ASAP7_75t_SL g1935 ( 
.A(n_1189),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1237),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1238),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1253),
.Y(n_1938)
);

CKINVDCx20_ASAP7_75t_R g1939 ( 
.A(n_1362),
.Y(n_1939)
);

CKINVDCx14_ASAP7_75t_R g1940 ( 
.A(n_1239),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1291),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1380),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1249),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1249),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1295),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1421),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_1441),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1298),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1300),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1488),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1456),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1249),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1312),
.Y(n_1953)
);

CKINVDCx20_ASAP7_75t_R g1954 ( 
.A(n_1458),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1319),
.Y(n_1955)
);

INVxp33_ASAP7_75t_SL g1956 ( 
.A(n_923),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1491),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1249),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1325),
.Y(n_1959)
);

CKINVDCx14_ASAP7_75t_R g1960 ( 
.A(n_1239),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1333),
.Y(n_1961)
);

INVxp67_ASAP7_75t_SL g1962 ( 
.A(n_1339),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1342),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1073),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1838),
.Y(n_1965)
);

BUFx2_ASAP7_75t_L g1966 ( 
.A(n_1830),
.Y(n_1966)
);

INVx5_ASAP7_75t_L g1967 ( 
.A(n_1805),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1781),
.A2(n_930),
.B(n_921),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1940),
.B(n_1266),
.Y(n_1969)
);

OAI22x1_ASAP7_75t_R g1970 ( 
.A1(n_1774),
.A2(n_1011),
.B1(n_1041),
.B2(n_1002),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1960),
.B(n_1492),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1786),
.A2(n_950),
.B(n_940),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1850),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1848),
.Y(n_1974)
);

AND2x6_ASAP7_75t_L g1975 ( 
.A(n_1800),
.B(n_932),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1833),
.Y(n_1976)
);

AND2x6_ASAP7_75t_L g1977 ( 
.A(n_1871),
.B(n_932),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1853),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1856),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1813),
.A2(n_1780),
.B1(n_1791),
.B2(n_1770),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1862),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1817),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1864),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1817),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1870),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1779),
.B(n_1712),
.Y(n_1986)
);

OAI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1801),
.A2(n_971),
.B(n_967),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1874),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1883),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1921),
.A2(n_1511),
.B1(n_1104),
.B2(n_1146),
.Y(n_1990)
);

BUFx2_ASAP7_75t_L g1991 ( 
.A(n_1863),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1821),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1884),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1826),
.A2(n_959),
.B(n_949),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1943),
.Y(n_1995)
);

INVx5_ASAP7_75t_L g1996 ( 
.A(n_1831),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1886),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1819),
.B(n_1674),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1923),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1775),
.B(n_1895),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1815),
.B(n_1839),
.Y(n_2001)
);

CKINVDCx6p67_ASAP7_75t_R g2002 ( 
.A(n_1771),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1833),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1927),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1865),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1930),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1777),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1833),
.Y(n_2008)
);

INVx3_ASAP7_75t_L g2009 ( 
.A(n_1782),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1852),
.B(n_1761),
.Y(n_2010)
);

OAI22x1_ASAP7_75t_SL g2011 ( 
.A1(n_1784),
.A2(n_1123),
.B1(n_1152),
.B2(n_1150),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1911),
.Y(n_2012)
);

OA21x2_ASAP7_75t_L g2013 ( 
.A1(n_1828),
.A2(n_959),
.B(n_949),
.Y(n_2013)
);

BUFx8_ASAP7_75t_L g2014 ( 
.A(n_1787),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1920),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1879),
.B(n_1328),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1944),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1788),
.Y(n_2018)
);

OA21x2_ASAP7_75t_L g2019 ( 
.A1(n_1832),
.A2(n_1082),
.B(n_989),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1935),
.B(n_1075),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1887),
.Y(n_2021)
);

OAI22x1_ASAP7_75t_L g2022 ( 
.A1(n_1914),
.A2(n_968),
.B1(n_1124),
.B2(n_937),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1964),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1952),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1964),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1962),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1958),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1898),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1900),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1882),
.B(n_1276),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1789),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1964),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1772),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1816),
.Y(n_2034)
);

CKINVDCx16_ASAP7_75t_R g2035 ( 
.A(n_1843),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1827),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1834),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_1807),
.A2(n_1173),
.B1(n_1715),
.B2(n_1202),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1773),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1835),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1907),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1844),
.B(n_1496),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1790),
.B(n_1197),
.Y(n_2043)
);

AND2x6_ASAP7_75t_L g2044 ( 
.A(n_1792),
.B(n_945),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1776),
.Y(n_2045)
);

CKINVDCx20_ASAP7_75t_R g2046 ( 
.A(n_1824),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1836),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1837),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1840),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1793),
.B(n_1753),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1875),
.B(n_1344),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1794),
.B(n_1496),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_SL g2053 ( 
.A(n_1785),
.B(n_1778),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1841),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1842),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1846),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1795),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_1847),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1913),
.B(n_1156),
.Y(n_2059)
);

CKINVDCx8_ASAP7_75t_R g2060 ( 
.A(n_1942),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1868),
.B(n_1288),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_1925),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_1810),
.Y(n_2063)
);

BUFx2_ASAP7_75t_L g2064 ( 
.A(n_1951),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1889),
.B(n_1315),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1849),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1851),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1796),
.Y(n_2068)
);

BUFx6f_ASAP7_75t_L g2069 ( 
.A(n_1855),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1797),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1857),
.Y(n_2071)
);

AND2x6_ASAP7_75t_L g2072 ( 
.A(n_1798),
.B(n_945),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1957),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1924),
.B(n_1156),
.Y(n_2074)
);

INVx3_ASAP7_75t_L g2075 ( 
.A(n_1799),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1802),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1932),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_1829),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_SL g2079 ( 
.A(n_1956),
.B(n_1499),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1893),
.B(n_1349),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1804),
.B(n_975),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1806),
.B(n_978),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_1845),
.Y(n_2083)
);

OA21x2_ASAP7_75t_L g2084 ( 
.A1(n_1808),
.A2(n_1082),
.B(n_989),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1858),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1809),
.B(n_1811),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1812),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_1946),
.B(n_1321),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1814),
.Y(n_2089)
);

OA21x2_ASAP7_75t_L g2090 ( 
.A1(n_1818),
.A2(n_1398),
.B(n_1096),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1950),
.B(n_1280),
.Y(n_2091)
);

BUFx3_ASAP7_75t_L g2092 ( 
.A(n_1820),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1822),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1823),
.B(n_1280),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1859),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_SL g2096 ( 
.A(n_1783),
.B(n_1507),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1880),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_1896),
.Y(n_2098)
);

INVx6_ASAP7_75t_L g2099 ( 
.A(n_1803),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1825),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1860),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1861),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1866),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1867),
.B(n_1354),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1869),
.B(n_1872),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1873),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1876),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1877),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1878),
.B(n_986),
.Y(n_2109)
);

INVx6_ASAP7_75t_L g2110 ( 
.A(n_1881),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1885),
.Y(n_2111)
);

OA21x2_ASAP7_75t_L g2112 ( 
.A1(n_1888),
.A2(n_1398),
.B(n_1096),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1890),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1963),
.B(n_998),
.Y(n_2114)
);

AND2x6_ASAP7_75t_L g2115 ( 
.A(n_1891),
.B(n_979),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1892),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1894),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1897),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1899),
.Y(n_2119)
);

BUFx6f_ASAP7_75t_L g2120 ( 
.A(n_1901),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_1903),
.B(n_1372),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_1904),
.B(n_1729),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1905),
.B(n_1329),
.Y(n_2123)
);

OA21x2_ASAP7_75t_L g2124 ( 
.A1(n_1906),
.A2(n_1025),
.B(n_1014),
.Y(n_2124)
);

OAI21x1_ASAP7_75t_L g2125 ( 
.A1(n_1908),
.A2(n_1042),
.B(n_1027),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_1910),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1912),
.Y(n_2127)
);

BUFx3_ASAP7_75t_L g2128 ( 
.A(n_1915),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_1916),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1854),
.A2(n_1187),
.B1(n_1264),
.B2(n_1231),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1919),
.Y(n_2131)
);

BUFx12f_ASAP7_75t_L g2132 ( 
.A(n_1902),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_1922),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1926),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1928),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1929),
.B(n_1953),
.Y(n_2136)
);

BUFx8_ASAP7_75t_L g2137 ( 
.A(n_1931),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1933),
.B(n_1329),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1934),
.Y(n_2139)
);

OA21x2_ASAP7_75t_L g2140 ( 
.A1(n_1936),
.A2(n_1047),
.B(n_1045),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1937),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1938),
.B(n_1059),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1941),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_SL g2144 ( 
.A1(n_1909),
.A2(n_1269),
.B1(n_1272),
.B2(n_1265),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1945),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1948),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1949),
.B(n_1100),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_1955),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_1961),
.B(n_1959),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_1917),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1918),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1939),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1947),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1954),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1838),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1833),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1911),
.Y(n_2157)
);

OAI22x1_ASAP7_75t_R g2158 ( 
.A1(n_1774),
.A2(n_1287),
.B1(n_1304),
.B2(n_1283),
.Y(n_2158)
);

OAI22x1_ASAP7_75t_R g2159 ( 
.A1(n_1774),
.A2(n_1313),
.B1(n_1377),
.B2(n_1309),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1770),
.A2(n_1404),
.B1(n_1418),
.B2(n_1389),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1838),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_1817),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1838),
.Y(n_2163)
);

INVx5_ASAP7_75t_L g2164 ( 
.A(n_1805),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_1833),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_1911),
.Y(n_2166)
);

BUFx8_ASAP7_75t_L g2167 ( 
.A(n_1800),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1838),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1940),
.B(n_1106),
.Y(n_2169)
);

OAI21x1_ASAP7_75t_L g2170 ( 
.A1(n_1781),
.A2(n_1136),
.B(n_1132),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1838),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1850),
.Y(n_2172)
);

INVx4_ASAP7_75t_L g2173 ( 
.A(n_1821),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_1895),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1850),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_1770),
.A2(n_1532),
.B1(n_1622),
.B2(n_1434),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1833),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1850),
.Y(n_2178)
);

INVxp33_ASAP7_75t_SL g2179 ( 
.A(n_1821),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_1813),
.A2(n_1681),
.B1(n_1685),
.B2(n_1654),
.Y(n_2180)
);

INVx5_ASAP7_75t_L g2181 ( 
.A(n_1805),
.Y(n_2181)
);

CKINVDCx11_ASAP7_75t_R g2182 ( 
.A(n_1824),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1817),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1850),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_1800),
.B(n_1084),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1805),
.B(n_1365),
.Y(n_2186)
);

OA21x2_ASAP7_75t_L g2187 ( 
.A1(n_1826),
.A2(n_1160),
.B(n_1142),
.Y(n_2187)
);

AOI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_1813),
.A2(n_1728),
.B1(n_1743),
.B2(n_1590),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_1833),
.Y(n_2189)
);

NAND2xp33_ASAP7_75t_L g2190 ( 
.A(n_1821),
.B(n_1339),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1838),
.Y(n_2191)
);

INVx5_ASAP7_75t_L g2192 ( 
.A(n_1805),
.Y(n_2192)
);

INVxp33_ASAP7_75t_SL g2193 ( 
.A(n_1821),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1850),
.Y(n_2194)
);

CKINVDCx11_ASAP7_75t_R g2195 ( 
.A(n_1824),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1850),
.Y(n_2196)
);

BUFx3_ASAP7_75t_L g2197 ( 
.A(n_1817),
.Y(n_2197)
);

BUFx6f_ASAP7_75t_L g2198 ( 
.A(n_1833),
.Y(n_2198)
);

OA21x2_ASAP7_75t_L g2199 ( 
.A1(n_1826),
.A2(n_1179),
.B(n_1175),
.Y(n_2199)
);

OA21x2_ASAP7_75t_L g2200 ( 
.A1(n_1826),
.A2(n_1192),
.B(n_1182),
.Y(n_2200)
);

OA21x2_ASAP7_75t_L g2201 ( 
.A1(n_1826),
.A2(n_1211),
.B(n_1194),
.Y(n_2201)
);

CKINVDCx16_ASAP7_75t_R g2202 ( 
.A(n_1805),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1838),
.Y(n_2203)
);

OAI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_1770),
.A2(n_1203),
.B1(n_1242),
.B2(n_1161),
.Y(n_2204)
);

CKINVDCx20_ASAP7_75t_R g2205 ( 
.A(n_1824),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_SL g2206 ( 
.A1(n_1771),
.A2(n_1360),
.B1(n_1403),
.B2(n_1289),
.Y(n_2206)
);

OA21x2_ASAP7_75t_L g2207 ( 
.A1(n_1826),
.A2(n_1248),
.B(n_1244),
.Y(n_2207)
);

CKINVDCx11_ASAP7_75t_R g2208 ( 
.A(n_1824),
.Y(n_2208)
);

OA21x2_ASAP7_75t_L g2209 ( 
.A1(n_1826),
.A2(n_1296),
.B(n_1273),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1813),
.A2(n_1610),
.B1(n_1613),
.B2(n_1566),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_SL g2211 ( 
.A1(n_1771),
.A2(n_1537),
.B1(n_1644),
.B2(n_1519),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1838),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1838),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1838),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1850),
.Y(n_2215)
);

INVx3_ASAP7_75t_L g2216 ( 
.A(n_1817),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1838),
.Y(n_2217)
);

BUFx3_ASAP7_75t_L g2218 ( 
.A(n_1817),
.Y(n_2218)
);

AOI22x1_ASAP7_75t_SL g2219 ( 
.A1(n_1824),
.A2(n_1007),
.B1(n_1017),
.B2(n_933),
.Y(n_2219)
);

BUFx2_ASAP7_75t_L g2220 ( 
.A(n_1830),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_1800),
.B(n_1230),
.Y(n_2221)
);

BUFx3_ASAP7_75t_L g2222 ( 
.A(n_1817),
.Y(n_2222)
);

BUFx2_ASAP7_75t_L g2223 ( 
.A(n_1830),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1850),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1805),
.B(n_1365),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1838),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1805),
.B(n_1462),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_1833),
.Y(n_2228)
);

INVx6_ASAP7_75t_L g2229 ( 
.A(n_1831),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1838),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1838),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_1770),
.A2(n_1689),
.B1(n_929),
.B2(n_935),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_1805),
.B(n_1311),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1850),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1817),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_1830),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_1895),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1850),
.Y(n_2238)
);

OAI21x1_ASAP7_75t_L g2239 ( 
.A1(n_1781),
.A2(n_1322),
.B(n_1316),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1940),
.B(n_1336),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1940),
.B(n_1340),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1850),
.Y(n_2242)
);

INVx4_ASAP7_75t_L g2243 ( 
.A(n_1821),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1850),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1850),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1838),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1850),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1850),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1838),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1911),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1838),
.Y(n_2251)
);

OA21x2_ASAP7_75t_L g2252 ( 
.A1(n_1826),
.A2(n_1378),
.B(n_1352),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1850),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1838),
.Y(n_2254)
);

BUFx6f_ASAP7_75t_L g2255 ( 
.A(n_1833),
.Y(n_2255)
);

INVx2_ASAP7_75t_SL g2256 ( 
.A(n_1800),
.Y(n_2256)
);

OAI22x1_ASAP7_75t_SL g2257 ( 
.A1(n_1813),
.A2(n_939),
.B1(n_942),
.B2(n_928),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1838),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1838),
.Y(n_2259)
);

AOI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_1813),
.A2(n_1682),
.B1(n_1711),
.B2(n_1642),
.Y(n_2260)
);

INVx4_ASAP7_75t_L g2261 ( 
.A(n_1821),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_1805),
.B(n_1462),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1850),
.Y(n_2263)
);

AND2x6_ASAP7_75t_L g2264 ( 
.A(n_1800),
.B(n_979),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1838),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1850),
.Y(n_2266)
);

INVx5_ASAP7_75t_L g2267 ( 
.A(n_1805),
.Y(n_2267)
);

BUFx6f_ASAP7_75t_L g2268 ( 
.A(n_1833),
.Y(n_2268)
);

AOI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_1813),
.A2(n_1745),
.B1(n_943),
.B2(n_976),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1800),
.B(n_1230),
.Y(n_2270)
);

NAND2xp33_ASAP7_75t_SL g2271 ( 
.A(n_1807),
.B(n_1339),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1850),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1850),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1805),
.B(n_1505),
.Y(n_2274)
);

OAI21x1_ASAP7_75t_L g2275 ( 
.A1(n_1781),
.A2(n_1381),
.B(n_1379),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1940),
.B(n_1409),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1940),
.B(n_1410),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1838),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1838),
.Y(n_2279)
);

AOI22x1_ASAP7_75t_SL g2280 ( 
.A1(n_1824),
.A2(n_994),
.B1(n_1009),
.B2(n_960),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_1833),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1850),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_1833),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1838),
.Y(n_2284)
);

NAND2x1p5_ASAP7_75t_L g2285 ( 
.A(n_1817),
.B(n_961),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1838),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1833),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1838),
.Y(n_2288)
);

OA21x2_ASAP7_75t_L g2289 ( 
.A1(n_1826),
.A2(n_1476),
.B(n_1457),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1838),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1850),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1850),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_1895),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1940),
.B(n_1480),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_1817),
.Y(n_2295)
);

BUFx6f_ASAP7_75t_L g2296 ( 
.A(n_1833),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_1833),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_1833),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_1911),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1940),
.B(n_1484),
.Y(n_2300)
);

HB1xp67_ASAP7_75t_L g2301 ( 
.A(n_1895),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_1895),
.Y(n_2302)
);

AND2x6_ASAP7_75t_L g2303 ( 
.A(n_1800),
.B(n_1108),
.Y(n_2303)
);

INVx3_ASAP7_75t_L g2304 ( 
.A(n_1817),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2036),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_2012),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_2015),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_2036),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_2157),
.Y(n_2309)
);

BUFx10_ASAP7_75t_L g2310 ( 
.A(n_2229),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_2166),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_2250),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_1976),
.Y(n_2313)
);

BUFx10_ASAP7_75t_L g2314 ( 
.A(n_2099),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1973),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2033),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_2299),
.Y(n_2317)
);

HB1xp67_ASAP7_75t_L g2318 ( 
.A(n_2174),
.Y(n_2318)
);

CKINVDCx20_ASAP7_75t_R g2319 ( 
.A(n_2046),
.Y(n_2319)
);

CKINVDCx20_ASAP7_75t_R g2320 ( 
.A(n_2205),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_1976),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_2182),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2039),
.Y(n_2323)
);

INVx3_ASAP7_75t_L g2324 ( 
.A(n_2003),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_2003),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_R g2326 ( 
.A(n_2060),
.B(n_924),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2045),
.Y(n_2327)
);

INVx4_ASAP7_75t_L g2328 ( 
.A(n_1967),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2068),
.Y(n_2329)
);

INVx8_ASAP7_75t_L g2330 ( 
.A(n_1967),
.Y(n_2330)
);

BUFx2_ASAP7_75t_L g2331 ( 
.A(n_2062),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_R g2332 ( 
.A(n_2035),
.B(n_926),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2070),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_2008),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2195),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2123),
.B(n_1200),
.Y(n_2336)
);

BUFx2_ASAP7_75t_L g2337 ( 
.A(n_1966),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2076),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_2208),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_2078),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_2097),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_2179),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_2193),
.Y(n_2343)
);

CKINVDCx20_ASAP7_75t_R g2344 ( 
.A(n_2202),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1978),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_2008),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2089),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_2132),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_R g2349 ( 
.A(n_1992),
.B(n_927),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_2064),
.Y(n_2350)
);

BUFx3_ASAP7_75t_L g2351 ( 
.A(n_2197),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2093),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_2150),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2106),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_2002),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2108),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_1991),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_2237),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_R g2359 ( 
.A(n_2053),
.B(n_931),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_2029),
.Y(n_2360)
);

OAI22xp5_ASAP7_75t_SL g2361 ( 
.A1(n_2144),
.A2(n_953),
.B1(n_1008),
.B2(n_991),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2220),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_2223),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2134),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_R g2365 ( 
.A(n_2079),
.B(n_934),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_2236),
.Y(n_2366)
);

BUFx2_ASAP7_75t_L g2367 ( 
.A(n_2293),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2141),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1979),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_R g2370 ( 
.A(n_2096),
.B(n_936),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2083),
.Y(n_2371)
);

NAND2xp33_ASAP7_75t_R g2372 ( 
.A(n_2063),
.B(n_948),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_1981),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_2098),
.Y(n_2374)
);

NOR2xp67_ASAP7_75t_L g2375 ( 
.A(n_1996),
.B(n_992),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_2173),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2243),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_1995),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2261),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2042),
.B(n_1020),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2017),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2095),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2101),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_2073),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_R g2385 ( 
.A(n_2164),
.B(n_944),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2024),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2167),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_R g2388 ( 
.A(n_2164),
.B(n_946),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2059),
.B(n_919),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_1996),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2027),
.Y(n_2391)
);

AND3x2_ASAP7_75t_L g2392 ( 
.A(n_2010),
.B(n_1671),
.C(n_1051),
.Y(n_2392)
);

CKINVDCx20_ASAP7_75t_R g2393 ( 
.A(n_2005),
.Y(n_2393)
);

OAI22xp33_ASAP7_75t_L g2394 ( 
.A1(n_2269),
.A2(n_1023),
.B1(n_1040),
.B2(n_966),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2103),
.Y(n_2395)
);

CKINVDCx16_ASAP7_75t_R g2396 ( 
.A(n_1970),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2301),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_2021),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_R g2399 ( 
.A(n_2181),
.B(n_2192),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2107),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2111),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_R g2402 ( 
.A(n_2181),
.B(n_963),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_2028),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2302),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_L g2405 ( 
.A(n_2080),
.B(n_1486),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_2041),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_2160),
.Y(n_2407)
);

CKINVDCx20_ASAP7_75t_R g2408 ( 
.A(n_2192),
.Y(n_2408)
);

NOR2xp67_ASAP7_75t_L g2409 ( 
.A(n_2267),
.B(n_1306),
.Y(n_2409)
);

INVxp67_ASAP7_75t_L g2410 ( 
.A(n_2077),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_R g2411 ( 
.A(n_2267),
.B(n_965),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2176),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2172),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2113),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2116),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2117),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_2218),
.Y(n_2417)
);

BUFx10_ASAP7_75t_L g2418 ( 
.A(n_2061),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2256),
.B(n_919),
.Y(n_2419)
);

CKINVDCx20_ASAP7_75t_R g2420 ( 
.A(n_2210),
.Y(n_2420)
);

NAND2xp33_ASAP7_75t_R g2421 ( 
.A(n_2001),
.B(n_954),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_2260),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2175),
.Y(n_2423)
);

NOR2xp67_ASAP7_75t_L g2424 ( 
.A(n_1980),
.B(n_1331),
.Y(n_2424)
);

HB1xp67_ASAP7_75t_L g2425 ( 
.A(n_2000),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_2222),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_1975),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_1975),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_1977),
.Y(n_2429)
);

NAND2xp33_ASAP7_75t_R g2430 ( 
.A(n_2186),
.B(n_955),
.Y(n_2430)
);

BUFx3_ASAP7_75t_L g2431 ( 
.A(n_2110),
.Y(n_2431)
);

CKINVDCx5p33_ASAP7_75t_R g2432 ( 
.A(n_1977),
.Y(n_2432)
);

NOR2xp67_ASAP7_75t_L g2433 ( 
.A(n_2148),
.B(n_1982),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2118),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_R g2435 ( 
.A(n_2271),
.B(n_973),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2178),
.Y(n_2436)
);

CKINVDCx20_ASAP7_75t_R g2437 ( 
.A(n_2188),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2119),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_2264),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_2264),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_2303),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_2303),
.Y(n_2442)
);

CKINVDCx20_ASAP7_75t_R g2443 ( 
.A(n_1990),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_2219),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2280),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_2130),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_2018),
.Y(n_2447)
);

AOI21x1_ASAP7_75t_L g2448 ( 
.A1(n_2125),
.A2(n_1516),
.B(n_1515),
.Y(n_2448)
);

CKINVDCx5p33_ASAP7_75t_R g2449 ( 
.A(n_2057),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2225),
.B(n_925),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2127),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_R g2452 ( 
.A(n_1984),
.B(n_980),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2131),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_2162),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_2092),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2227),
.B(n_925),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2139),
.Y(n_2457)
);

AND2x6_ASAP7_75t_L g2458 ( 
.A(n_2138),
.B(n_1108),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_2151),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2184),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_2153),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_2154),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2143),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2146),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_R g2465 ( 
.A(n_2183),
.B(n_2216),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2067),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2067),
.Y(n_2467)
);

XOR2xp5_ASAP7_75t_L g2468 ( 
.A(n_2180),
.B(n_956),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2137),
.Y(n_2469)
);

BUFx3_ASAP7_75t_L g2470 ( 
.A(n_2235),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2069),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2152),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_2257),
.Y(n_2473)
);

BUFx10_ASAP7_75t_L g2474 ( 
.A(n_2233),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2102),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_2128),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2274),
.B(n_1016),
.Y(n_2477)
);

CKINVDCx20_ASAP7_75t_R g2478 ( 
.A(n_2038),
.Y(n_2478)
);

BUFx10_ASAP7_75t_L g2479 ( 
.A(n_1986),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2129),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_2014),
.Y(n_2481)
);

INVx4_ASAP7_75t_L g2482 ( 
.A(n_2295),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2069),
.Y(n_2483)
);

NOR2xp67_ASAP7_75t_L g2484 ( 
.A(n_2304),
.B(n_1397),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2071),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2071),
.Y(n_2486)
);

INVx2_ASAP7_75t_SL g2487 ( 
.A(n_2074),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2011),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2085),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2085),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_2120),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2120),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2126),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2126),
.Y(n_2494)
);

CKINVDCx20_ASAP7_75t_R g2495 ( 
.A(n_2158),
.Y(n_2495)
);

BUFx10_ASAP7_75t_L g2496 ( 
.A(n_1998),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2133),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2133),
.Y(n_2498)
);

CKINVDCx5p33_ASAP7_75t_R g2499 ( 
.A(n_2135),
.Y(n_2499)
);

NAND2xp33_ASAP7_75t_R g2500 ( 
.A(n_2051),
.B(n_972),
.Y(n_2500)
);

CKINVDCx5p33_ASAP7_75t_R g2501 ( 
.A(n_2135),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_2145),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2145),
.Y(n_2503)
);

AND3x2_ASAP7_75t_L g2504 ( 
.A(n_2091),
.B(n_1051),
.C(n_1037),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_R g2505 ( 
.A(n_2007),
.B(n_981),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2232),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_R g2507 ( 
.A(n_2009),
.B(n_985),
.Y(n_2507)
);

AO21x2_ASAP7_75t_L g2508 ( 
.A1(n_1968),
.A2(n_1987),
.B(n_1972),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_2206),
.Y(n_2509)
);

CKINVDCx20_ASAP7_75t_R g2510 ( 
.A(n_2159),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_2211),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_1965),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_1969),
.Y(n_2513)
);

CKINVDCx20_ASAP7_75t_R g2514 ( 
.A(n_2262),
.Y(n_2514)
);

CKINVDCx20_ASAP7_75t_R g2515 ( 
.A(n_1971),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_2031),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_1974),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_2075),
.Y(n_2518)
);

CKINVDCx20_ASAP7_75t_R g2519 ( 
.A(n_2094),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2087),
.Y(n_2520)
);

AND2x6_ASAP7_75t_L g2521 ( 
.A(n_2105),
.B(n_1174),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_2100),
.Y(n_2522)
);

CKINVDCx5p33_ASAP7_75t_R g2523 ( 
.A(n_2169),
.Y(n_2523)
);

BUFx10_ASAP7_75t_L g2524 ( 
.A(n_2016),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_2240),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2300),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_1983),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2194),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_R g2529 ( 
.A(n_2190),
.B(n_988),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2047),
.B(n_1105),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2196),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2241),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_1985),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_2043),
.Y(n_2534)
);

CKINVDCx20_ASAP7_75t_R g2535 ( 
.A(n_2050),
.Y(n_2535)
);

CKINVDCx20_ASAP7_75t_R g2536 ( 
.A(n_2020),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_2276),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2215),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_R g2539 ( 
.A(n_1988),
.B(n_1003),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_2277),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_2204),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2294),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_1989),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_1993),
.Y(n_2544)
);

INVxp67_ASAP7_75t_L g2545 ( 
.A(n_2149),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_1997),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_1999),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2004),
.Y(n_2548)
);

CKINVDCx20_ASAP7_75t_R g2549 ( 
.A(n_2052),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_2006),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2026),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2155),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2161),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2163),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_R g2555 ( 
.A(n_2168),
.B(n_1005),
.Y(n_2555)
);

CKINVDCx20_ASAP7_75t_R g2556 ( 
.A(n_2171),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2191),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_2203),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2212),
.Y(n_2559)
);

NAND2xp33_ASAP7_75t_R g2560 ( 
.A(n_2187),
.B(n_977),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2213),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2214),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2217),
.Y(n_2563)
);

BUFx10_ASAP7_75t_L g2564 ( 
.A(n_2185),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2226),
.B(n_1517),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_2230),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2231),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_2246),
.Y(n_2568)
);

CKINVDCx20_ASAP7_75t_R g2569 ( 
.A(n_2249),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_L g2570 ( 
.A(n_2251),
.B(n_2254),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_2258),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2259),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2265),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_R g2574 ( 
.A(n_2278),
.B(n_1015),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2048),
.B(n_1367),
.Y(n_2575)
);

NAND2xp33_ASAP7_75t_SL g2576 ( 
.A(n_2136),
.B(n_987),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2279),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2284),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2030),
.Y(n_2579)
);

CKINVDCx20_ASAP7_75t_R g2580 ( 
.A(n_2286),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_R g2581 ( 
.A(n_2288),
.B(n_1022),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2290),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_2086),
.Y(n_2583)
);

CKINVDCx5p33_ASAP7_75t_R g2584 ( 
.A(n_2115),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2115),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_R g2586 ( 
.A(n_2049),
.B(n_1033),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2040),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_R g2588 ( 
.A(n_2109),
.B(n_1050),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2044),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_2142),
.Y(n_2590)
);

OAI22xp5_ASAP7_75t_SL g2591 ( 
.A1(n_2022),
.A2(n_1035),
.B1(n_1057),
.B2(n_1013),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_2044),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2224),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_R g2594 ( 
.A(n_2147),
.B(n_1052),
.Y(n_2594)
);

XNOR2xp5_ASAP7_75t_L g2595 ( 
.A(n_2285),
.B(n_990),
.Y(n_2595)
);

CKINVDCx20_ASAP7_75t_R g2596 ( 
.A(n_2124),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2072),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2037),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2072),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_2221),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_2270),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_2040),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2054),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2055),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_2056),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2066),
.Y(n_2606)
);

BUFx6f_ASAP7_75t_L g2607 ( 
.A(n_2023),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2034),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2234),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_R g2610 ( 
.A(n_2081),
.B(n_1053),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2512),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_SL g2612 ( 
.A(n_2376),
.B(n_2056),
.Y(n_2612)
);

BUFx3_ASAP7_75t_L g2613 ( 
.A(n_2314),
.Y(n_2613)
);

BUFx6f_ASAP7_75t_SL g2614 ( 
.A(n_2314),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2405),
.B(n_2058),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2517),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2315),
.Y(n_2617)
);

AOI22xp33_ASAP7_75t_L g2618 ( 
.A1(n_2407),
.A2(n_2140),
.B1(n_2200),
.B2(n_2199),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2310),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2310),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2545),
.B(n_2058),
.Y(n_2621)
);

HB1xp67_ASAP7_75t_L g2622 ( 
.A(n_2367),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2527),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2345),
.Y(n_2624)
);

INVx4_ASAP7_75t_L g2625 ( 
.A(n_2330),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2319),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_L g2627 ( 
.A1(n_2446),
.A2(n_2201),
.B1(n_2209),
.B2(n_2207),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2533),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2513),
.B(n_2082),
.Y(n_2629)
);

INVx2_ASAP7_75t_SL g2630 ( 
.A(n_2331),
.Y(n_2630)
);

INVx4_ASAP7_75t_L g2631 ( 
.A(n_2330),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2431),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2583),
.B(n_2114),
.Y(n_2633)
);

INVx3_ASAP7_75t_L g2634 ( 
.A(n_2351),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2551),
.Y(n_2635)
);

BUFx2_ASAP7_75t_L g2636 ( 
.A(n_2320),
.Y(n_2636)
);

BUFx3_ASAP7_75t_L g2637 ( 
.A(n_2330),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2523),
.B(n_996),
.Y(n_2638)
);

INVx4_ASAP7_75t_L g2639 ( 
.A(n_2353),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2525),
.B(n_2252),
.Y(n_2640)
);

INVx4_ASAP7_75t_L g2641 ( 
.A(n_2306),
.Y(n_2641)
);

INVx4_ASAP7_75t_L g2642 ( 
.A(n_2307),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2526),
.B(n_2289),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2553),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_2532),
.B(n_999),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2554),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2369),
.Y(n_2647)
);

INVx1_ASAP7_75t_SL g2648 ( 
.A(n_2337),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2373),
.Y(n_2649)
);

OR2x2_ASAP7_75t_L g2650 ( 
.A(n_2318),
.B(n_2065),
.Y(n_2650)
);

BUFx6f_ASAP7_75t_L g2651 ( 
.A(n_2587),
.Y(n_2651)
);

BUFx3_ASAP7_75t_L g2652 ( 
.A(n_2340),
.Y(n_2652)
);

BUFx6f_ASAP7_75t_L g2653 ( 
.A(n_2417),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2537),
.B(n_2112),
.Y(n_2654)
);

INVx4_ASAP7_75t_L g2655 ( 
.A(n_2309),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2540),
.B(n_1994),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2377),
.B(n_1000),
.Y(n_2657)
);

BUFx3_ASAP7_75t_L g2658 ( 
.A(n_2341),
.Y(n_2658)
);

AND2x4_ASAP7_75t_L g2659 ( 
.A(n_2344),
.B(n_2104),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_L g2660 ( 
.A(n_2542),
.B(n_1001),
.Y(n_2660)
);

AND2x6_ASAP7_75t_L g2661 ( 
.A(n_2419),
.B(n_1174),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2418),
.B(n_1012),
.Y(n_2662)
);

INVx4_ASAP7_75t_L g2663 ( 
.A(n_2311),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2378),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2381),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2557),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2559),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2386),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2418),
.B(n_1018),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2325),
.Y(n_2670)
);

NAND2x1p5_ASAP7_75t_L g2671 ( 
.A(n_2328),
.B(n_2121),
.Y(n_2671)
);

BUFx4f_ASAP7_75t_L g2672 ( 
.A(n_2336),
.Y(n_2672)
);

BUFx3_ASAP7_75t_L g2673 ( 
.A(n_2312),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2562),
.Y(n_2674)
);

OAI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2506),
.A2(n_1074),
.B1(n_1084),
.B2(n_1037),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2458),
.B(n_2013),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2572),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_SL g2678 ( 
.A(n_2379),
.B(n_1021),
.Y(n_2678)
);

NAND2xp33_ASAP7_75t_L g2679 ( 
.A(n_2317),
.B(n_1339),
.Y(n_2679)
);

INVx2_ASAP7_75t_SL g2680 ( 
.A(n_2479),
.Y(n_2680)
);

INVx2_ASAP7_75t_SL g2681 ( 
.A(n_2479),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2425),
.B(n_2088),
.Y(n_2682)
);

OR2x6_ASAP7_75t_L g2683 ( 
.A(n_2328),
.B(n_2122),
.Y(n_2683)
);

AND2x2_ASAP7_75t_SL g2684 ( 
.A(n_2396),
.B(n_1184),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2408),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2573),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2410),
.B(n_1028),
.Y(n_2687)
);

OR2x6_ASAP7_75t_L g2688 ( 
.A(n_2579),
.B(n_1074),
.Y(n_2688)
);

INVx4_ASAP7_75t_L g2689 ( 
.A(n_2490),
.Y(n_2689)
);

INVxp67_ASAP7_75t_SL g2690 ( 
.A(n_2433),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2578),
.Y(n_2691)
);

CKINVDCx20_ASAP7_75t_R g2692 ( 
.A(n_2342),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_L g2693 ( 
.A(n_2487),
.B(n_1030),
.Y(n_2693)
);

BUFx4f_ASAP7_75t_L g2694 ( 
.A(n_2336),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2357),
.B(n_1347),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2582),
.Y(n_2696)
);

INVx4_ASAP7_75t_L g2697 ( 
.A(n_2491),
.Y(n_2697)
);

NAND2xp33_ASAP7_75t_L g2698 ( 
.A(n_2349),
.B(n_1368),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_2475),
.B(n_1032),
.Y(n_2699)
);

NAND2xp33_ASAP7_75t_L g2700 ( 
.A(n_2521),
.B(n_1368),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2371),
.Y(n_2701)
);

BUFx2_ASAP7_75t_L g2702 ( 
.A(n_2374),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2382),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2391),
.Y(n_2704)
);

INVx3_ASAP7_75t_L g2705 ( 
.A(n_2564),
.Y(n_2705)
);

AND2x4_ASAP7_75t_L g2706 ( 
.A(n_2360),
.B(n_1357),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2383),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_2325),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2395),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_L g2710 ( 
.A(n_2325),
.Y(n_2710)
);

CKINVDCx11_ASAP7_75t_R g2711 ( 
.A(n_2393),
.Y(n_2711)
);

CKINVDCx20_ASAP7_75t_R g2712 ( 
.A(n_2343),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2400),
.Y(n_2713)
);

OR2x6_ASAP7_75t_L g2714 ( 
.A(n_2450),
.B(n_1254),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2401),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2496),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2458),
.B(n_2019),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2413),
.Y(n_2718)
);

AO21x2_ASAP7_75t_L g2719 ( 
.A1(n_2448),
.A2(n_2239),
.B(n_2170),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2564),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2414),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2394),
.A2(n_2521),
.B1(n_2412),
.B2(n_2416),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2423),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2458),
.B(n_2084),
.Y(n_2724)
);

INVx4_ASAP7_75t_L g2725 ( 
.A(n_2493),
.Y(n_2725)
);

INVx3_ASAP7_75t_L g2726 ( 
.A(n_2497),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2415),
.Y(n_2727)
);

AND2x4_ASAP7_75t_L g2728 ( 
.A(n_2362),
.B(n_1363),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2363),
.B(n_1366),
.Y(n_2729)
);

BUFx6f_ASAP7_75t_L g2730 ( 
.A(n_2334),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2366),
.B(n_1016),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2399),
.Y(n_2732)
);

AND2x4_ASAP7_75t_SL g2733 ( 
.A(n_2524),
.B(n_1026),
.Y(n_2733)
);

AND2x4_ASAP7_75t_L g2734 ( 
.A(n_2350),
.B(n_1383),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_L g2735 ( 
.A(n_2474),
.B(n_1043),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2458),
.B(n_2090),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2474),
.B(n_2534),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2434),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2438),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2600),
.Y(n_2740)
);

CKINVDCx16_ASAP7_75t_R g2741 ( 
.A(n_2332),
.Y(n_2741)
);

BUFx8_ASAP7_75t_SL g2742 ( 
.A(n_2322),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2451),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2436),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2453),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2380),
.B(n_2238),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2460),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2456),
.B(n_1026),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2457),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2528),
.Y(n_2750)
);

AO22x2_ASAP7_75t_L g2751 ( 
.A1(n_2468),
.A2(n_1387),
.B1(n_1395),
.B2(n_1393),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2463),
.Y(n_2752)
);

BUFx3_ASAP7_75t_L g2753 ( 
.A(n_2476),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2464),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2316),
.Y(n_2755)
);

BUFx6f_ASAP7_75t_L g2756 ( 
.A(n_2334),
.Y(n_2756)
);

BUFx2_ASAP7_75t_L g2757 ( 
.A(n_2358),
.Y(n_2757)
);

AND2x6_ASAP7_75t_L g2758 ( 
.A(n_2477),
.B(n_1401),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2531),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2535),
.B(n_1044),
.Y(n_2760)
);

INVx1_ASAP7_75t_SL g2761 ( 
.A(n_2601),
.Y(n_2761)
);

INVx5_ASAP7_75t_L g2762 ( 
.A(n_2524),
.Y(n_2762)
);

BUFx3_ASAP7_75t_L g2763 ( 
.A(n_2480),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2323),
.Y(n_2764)
);

BUFx3_ASAP7_75t_L g2765 ( 
.A(n_2335),
.Y(n_2765)
);

INVx3_ASAP7_75t_L g2766 ( 
.A(n_2498),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_L g2767 ( 
.A(n_2482),
.B(n_1046),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_2339),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2516),
.B(n_1061),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2538),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_L g2771 ( 
.A(n_2482),
.B(n_1063),
.Y(n_2771)
);

AND2x4_ASAP7_75t_L g2772 ( 
.A(n_2355),
.B(n_1400),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2570),
.B(n_2242),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2327),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_2326),
.Y(n_2775)
);

INVxp67_ASAP7_75t_SL g2776 ( 
.A(n_2308),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2499),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2454),
.B(n_1405),
.Y(n_2778)
);

BUFx4f_ASAP7_75t_L g2779 ( 
.A(n_2389),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2334),
.Y(n_2780)
);

NOR2xp33_ASAP7_75t_L g2781 ( 
.A(n_2536),
.B(n_1064),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2530),
.B(n_2575),
.Y(n_2782)
);

NAND2x1p5_ASAP7_75t_L g2783 ( 
.A(n_2470),
.B(n_2244),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_2348),
.B(n_1411),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2521),
.A2(n_2291),
.B1(n_2292),
.B2(n_2282),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2329),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2333),
.Y(n_2787)
);

BUFx6f_ASAP7_75t_L g2788 ( 
.A(n_2607),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2593),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2397),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_SL g2791 ( 
.A(n_2518),
.B(n_1066),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2338),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2347),
.Y(n_2793)
);

INVx4_ASAP7_75t_L g2794 ( 
.A(n_2501),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2609),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2354),
.B(n_2245),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2352),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2356),
.B(n_2247),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2364),
.B(n_2248),
.Y(n_2799)
);

AND2x4_ASAP7_75t_L g2800 ( 
.A(n_2502),
.B(n_1417),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2543),
.B(n_1069),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2398),
.B(n_1058),
.Y(n_2802)
);

AND2x2_ASAP7_75t_SL g2803 ( 
.A(n_2404),
.B(n_1274),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_SL g2804 ( 
.A(n_2520),
.B(n_1072),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2403),
.B(n_2406),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2496),
.B(n_1058),
.Y(n_2806)
);

INVx4_ASAP7_75t_L g2807 ( 
.A(n_2503),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2544),
.B(n_1076),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2384),
.B(n_1438),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2368),
.B(n_2253),
.Y(n_2810)
);

AND2x6_ASAP7_75t_L g2811 ( 
.A(n_2466),
.B(n_1401),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2546),
.B(n_2263),
.Y(n_2812)
);

INVx4_ASAP7_75t_L g2813 ( 
.A(n_2602),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2598),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2521),
.A2(n_2273),
.B1(n_2272),
.B2(n_2266),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2603),
.Y(n_2816)
);

INVx6_ASAP7_75t_L g2817 ( 
.A(n_2607),
.Y(n_2817)
);

INVx4_ASAP7_75t_L g2818 ( 
.A(n_2605),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2608),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2604),
.Y(n_2820)
);

OR2x2_ASAP7_75t_L g2821 ( 
.A(n_2422),
.B(n_1442),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2607),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2606),
.Y(n_2823)
);

OR2x6_ASAP7_75t_L g2824 ( 
.A(n_2361),
.B(n_1184),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2467),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_2359),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2308),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2471),
.Y(n_2828)
);

BUFx2_ASAP7_75t_L g2829 ( 
.A(n_2519),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2588),
.B(n_2594),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2483),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2522),
.B(n_1077),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2485),
.Y(n_2833)
);

AND2x6_ASAP7_75t_L g2834 ( 
.A(n_2486),
.B(n_1696),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_SL g2835 ( 
.A(n_2426),
.B(n_1079),
.Y(n_2835)
);

CKINVDCx5p33_ASAP7_75t_R g2836 ( 
.A(n_2390),
.Y(n_2836)
);

CKINVDCx5p33_ASAP7_75t_R g2837 ( 
.A(n_2387),
.Y(n_2837)
);

INVx4_ASAP7_75t_L g2838 ( 
.A(n_2447),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2449),
.B(n_1070),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2489),
.Y(n_2840)
);

INVx4_ASAP7_75t_L g2841 ( 
.A(n_2455),
.Y(n_2841)
);

INVx1_ASAP7_75t_SL g2842 ( 
.A(n_2472),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2547),
.B(n_1440),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_SL g2844 ( 
.A(n_2586),
.B(n_1081),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2492),
.Y(n_2845)
);

BUFx6f_ASAP7_75t_L g2846 ( 
.A(n_2305),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_2313),
.Y(n_2847)
);

INVx2_ASAP7_75t_SL g2848 ( 
.A(n_2465),
.Y(n_2848)
);

BUFx3_ASAP7_75t_L g2849 ( 
.A(n_2494),
.Y(n_2849)
);

BUFx2_ASAP7_75t_L g2850 ( 
.A(n_2590),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2313),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2321),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2321),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2324),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2469),
.Y(n_2855)
);

AND2x4_ASAP7_75t_L g2856 ( 
.A(n_2556),
.B(n_1432),
.Y(n_2856)
);

BUFx3_ASAP7_75t_L g2857 ( 
.A(n_2620),
.Y(n_2857)
);

OR2x6_ASAP7_75t_SL g2858 ( 
.A(n_2775),
.B(n_2481),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2805),
.B(n_2648),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2611),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2616),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2623),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2628),
.Y(n_2863)
);

OAI221xp5_ASAP7_75t_L g2864 ( 
.A1(n_2801),
.A2(n_2500),
.B1(n_2430),
.B2(n_2595),
.C(n_2421),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2630),
.B(n_2548),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2635),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2629),
.B(n_2550),
.Y(n_2867)
);

NOR2xp33_ASAP7_75t_L g2868 ( 
.A(n_2633),
.B(n_2515),
.Y(n_2868)
);

AND2x4_ASAP7_75t_L g2869 ( 
.A(n_2620),
.B(n_2569),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2644),
.Y(n_2870)
);

CKINVDCx5p33_ASAP7_75t_R g2871 ( 
.A(n_2742),
.Y(n_2871)
);

AND2x4_ASAP7_75t_L g2872 ( 
.A(n_2613),
.B(n_2580),
.Y(n_2872)
);

OA22x2_ASAP7_75t_L g2873 ( 
.A1(n_2842),
.A2(n_2511),
.B1(n_2509),
.B2(n_2591),
.Y(n_2873)
);

AND2x2_ASAP7_75t_SL g2874 ( 
.A(n_2684),
.B(n_2370),
.Y(n_2874)
);

INVx5_ASAP7_75t_L g2875 ( 
.A(n_2619),
.Y(n_2875)
);

OAI221xp5_ASAP7_75t_L g2876 ( 
.A1(n_2808),
.A2(n_2424),
.B1(n_2372),
.B2(n_2461),
.C(n_2459),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2782),
.B(n_2571),
.Y(n_2877)
);

AND2x4_ASAP7_75t_L g2878 ( 
.A(n_2637),
.B(n_2427),
.Y(n_2878)
);

AO22x1_ASAP7_75t_L g2879 ( 
.A1(n_2737),
.A2(n_2429),
.B1(n_2432),
.B2(n_2428),
.Y(n_2879)
);

AOI22xp33_ASAP7_75t_L g2880 ( 
.A1(n_2803),
.A2(n_2541),
.B1(n_2420),
.B2(n_2437),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2646),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2615),
.B(n_2552),
.Y(n_2882)
);

AO22x2_ASAP7_75t_L g2883 ( 
.A1(n_2821),
.A2(n_2478),
.B1(n_2443),
.B2(n_2495),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2617),
.Y(n_2884)
);

OR2x2_ASAP7_75t_SL g2885 ( 
.A(n_2741),
.B(n_2510),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2672),
.B(n_2558),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2624),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2694),
.B(n_2561),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2843),
.B(n_2567),
.Y(n_2889)
);

AO22x2_ASAP7_75t_L g2890 ( 
.A1(n_2856),
.A2(n_2560),
.B1(n_2514),
.B2(n_2596),
.Y(n_2890)
);

NAND2x1p5_ASAP7_75t_L g2891 ( 
.A(n_2689),
.B(n_2324),
.Y(n_2891)
);

NAND3xp33_ASAP7_75t_SL g2892 ( 
.A(n_2692),
.B(n_2365),
.C(n_2462),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2621),
.A2(n_2549),
.B1(n_2566),
.B2(n_2563),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2647),
.Y(n_2894)
);

INVx1_ASAP7_75t_SL g2895 ( 
.A(n_2622),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2666),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2667),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_SL g2898 ( 
.A(n_2779),
.B(n_2838),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2674),
.Y(n_2899)
);

CKINVDCx5p33_ASAP7_75t_R g2900 ( 
.A(n_2712),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2677),
.Y(n_2901)
);

NAND2x1p5_ASAP7_75t_L g2902 ( 
.A(n_2697),
.B(n_2725),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2757),
.Y(n_2903)
);

OAI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2703),
.A2(n_2577),
.B1(n_2568),
.B2(n_2440),
.Y(n_2904)
);

AND2x4_ASAP7_75t_L g2905 ( 
.A(n_2762),
.B(n_2626),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2686),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2691),
.B(n_2565),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2748),
.B(n_2439),
.Y(n_2908)
);

INVx4_ASAP7_75t_L g2909 ( 
.A(n_2614),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2696),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2707),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2709),
.Y(n_2912)
);

AND2x4_ASAP7_75t_L g2913 ( 
.A(n_2762),
.B(n_2441),
.Y(n_2913)
);

OR2x2_ASAP7_75t_SL g2914 ( 
.A(n_2809),
.B(n_2473),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_L g2915 ( 
.A(n_2638),
.B(n_2442),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2713),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2715),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2711),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2721),
.Y(n_2919)
);

INVx2_ASAP7_75t_SL g2920 ( 
.A(n_2636),
.Y(n_2920)
);

BUFx2_ASAP7_75t_L g2921 ( 
.A(n_2850),
.Y(n_2921)
);

AND2x4_ASAP7_75t_L g2922 ( 
.A(n_2753),
.B(n_2763),
.Y(n_2922)
);

INVxp67_ASAP7_75t_L g2923 ( 
.A(n_2790),
.Y(n_2923)
);

A2O1A1Ixp33_ASAP7_75t_L g2924 ( 
.A1(n_2767),
.A2(n_2576),
.B(n_2484),
.C(n_2275),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2727),
.Y(n_2925)
);

INVxp67_ASAP7_75t_L g2926 ( 
.A(n_2701),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2649),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2771),
.B(n_2589),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2664),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2738),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_2837),
.Y(n_2931)
);

INVx1_ASAP7_75t_SL g2932 ( 
.A(n_2702),
.Y(n_2932)
);

AO22x2_ASAP7_75t_L g2933 ( 
.A1(n_2751),
.A2(n_2488),
.B1(n_1201),
.B2(n_1245),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2739),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2743),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_R g2936 ( 
.A(n_2732),
.B(n_2584),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2645),
.B(n_2592),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2665),
.Y(n_2938)
);

BUFx3_ASAP7_75t_L g2939 ( 
.A(n_2673),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2745),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2749),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2752),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2754),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2668),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2755),
.Y(n_2945)
);

NAND2xp33_ASAP7_75t_L g2946 ( 
.A(n_2836),
.B(n_2597),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2704),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2764),
.Y(n_2948)
);

HB1xp67_ASAP7_75t_L g2949 ( 
.A(n_2829),
.Y(n_2949)
);

AND2x4_ASAP7_75t_L g2950 ( 
.A(n_2794),
.B(n_2585),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2774),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2786),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2718),
.Y(n_2953)
);

INVxp67_ASAP7_75t_L g2954 ( 
.A(n_2650),
.Y(n_2954)
);

INVxp67_ASAP7_75t_L g2955 ( 
.A(n_2652),
.Y(n_2955)
);

INVxp67_ASAP7_75t_L g2956 ( 
.A(n_2658),
.Y(n_2956)
);

OAI221xp5_ASAP7_75t_L g2957 ( 
.A1(n_2660),
.A2(n_2409),
.B1(n_2375),
.B2(n_1453),
.C(n_1463),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2625),
.Y(n_2958)
);

AND2x4_ASAP7_75t_L g2959 ( 
.A(n_2807),
.B(n_2599),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2781),
.B(n_2385),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2787),
.Y(n_2961)
);

BUFx8_ASAP7_75t_L g2962 ( 
.A(n_2855),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2792),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2723),
.Y(n_2964)
);

NAND2x1p5_ASAP7_75t_L g2965 ( 
.A(n_2813),
.B(n_2346),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_2760),
.B(n_2392),
.Y(n_2966)
);

INVxp67_ASAP7_75t_L g2967 ( 
.A(n_2740),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2773),
.B(n_2539),
.Y(n_2968)
);

NAND2x1p5_ASAP7_75t_L g2969 ( 
.A(n_2818),
.B(n_2346),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2744),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2793),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2797),
.Y(n_2972)
);

OR2x2_ASAP7_75t_L g2973 ( 
.A(n_2761),
.B(n_2444),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2814),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_SL g2975 ( 
.A(n_2841),
.B(n_2610),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2747),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2639),
.B(n_2504),
.Y(n_2977)
);

NAND3xp33_ASAP7_75t_L g2978 ( 
.A(n_2662),
.B(n_1162),
.C(n_1099),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2714),
.B(n_2445),
.Y(n_2979)
);

AND2x4_ASAP7_75t_L g2980 ( 
.A(n_2726),
.B(n_2508),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2816),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2750),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2669),
.B(n_2555),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_SL g2984 ( 
.A(n_2722),
.B(n_2505),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2823),
.Y(n_2985)
);

BUFx8_ASAP7_75t_L g2986 ( 
.A(n_2765),
.Y(n_2986)
);

AOI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2735),
.A2(n_1528),
.B1(n_1534),
.B2(n_1523),
.Y(n_2987)
);

NAND2x1p5_ASAP7_75t_L g2988 ( 
.A(n_2766),
.B(n_2023),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2661),
.B(n_2574),
.Y(n_2989)
);

BUFx8_ASAP7_75t_L g2990 ( 
.A(n_2768),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2796),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2661),
.B(n_2581),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2759),
.Y(n_2993)
);

BUFx3_ASAP7_75t_L g2994 ( 
.A(n_2632),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2661),
.B(n_2507),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2798),
.Y(n_2996)
);

CKINVDCx5p33_ASAP7_75t_R g2997 ( 
.A(n_2826),
.Y(n_2997)
);

AND2x4_ASAP7_75t_L g2998 ( 
.A(n_2777),
.B(n_2508),
.Y(n_2998)
);

OAI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2693),
.A2(n_2687),
.B1(n_2640),
.B2(n_2643),
.Y(n_2999)
);

OA22x2_ASAP7_75t_L g3000 ( 
.A1(n_2659),
.A2(n_1113),
.B1(n_1122),
.B2(n_1101),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2746),
.B(n_2452),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2770),
.Y(n_3002)
);

CKINVDCx5p33_ASAP7_75t_R g3003 ( 
.A(n_2641),
.Y(n_3003)
);

INVxp67_ASAP7_75t_L g3004 ( 
.A(n_2695),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2802),
.B(n_2388),
.Y(n_3005)
);

AND2x4_ASAP7_75t_L g3006 ( 
.A(n_2631),
.B(n_1433),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2799),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2685),
.B(n_1448),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2789),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2642),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2810),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2820),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2819),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2795),
.Y(n_3014)
);

OAI22x1_ASAP7_75t_L g3015 ( 
.A1(n_2800),
.A2(n_1221),
.B1(n_1263),
.B2(n_1208),
.Y(n_3015)
);

CKINVDCx5p33_ASAP7_75t_R g3016 ( 
.A(n_2655),
.Y(n_3016)
);

INVxp67_ASAP7_75t_L g3017 ( 
.A(n_2706),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2825),
.Y(n_3018)
);

A2O1A1Ixp33_ASAP7_75t_L g3019 ( 
.A1(n_2679),
.A2(n_1584),
.B(n_1601),
.C(n_1547),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2663),
.B(n_1087),
.Y(n_3020)
);

BUFx3_ASAP7_75t_L g3021 ( 
.A(n_2653),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2828),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2831),
.Y(n_3023)
);

AND2x4_ASAP7_75t_L g3024 ( 
.A(n_2848),
.B(n_1449),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2839),
.B(n_2402),
.Y(n_3025)
);

AND2x4_ASAP7_75t_L g3026 ( 
.A(n_2705),
.B(n_1465),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2833),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2812),
.B(n_2758),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2840),
.Y(n_3029)
);

AO22x2_ASAP7_75t_L g3030 ( 
.A1(n_2845),
.A2(n_2729),
.B1(n_2734),
.B2(n_2728),
.Y(n_3030)
);

NOR2x1p5_ASAP7_75t_L g3031 ( 
.A(n_2720),
.B(n_2411),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2758),
.B(n_2529),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2827),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2851),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2853),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2854),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2776),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2849),
.Y(n_3038)
);

OAI22x1_ASAP7_75t_L g3039 ( 
.A1(n_2772),
.A2(n_1133),
.B1(n_1154),
.B2(n_1103),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2846),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2847),
.Y(n_3041)
);

AO22x2_ASAP7_75t_L g3042 ( 
.A1(n_2654),
.A2(n_1201),
.B1(n_1254),
.B2(n_1234),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2852),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2731),
.B(n_1092),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_SL g3045 ( 
.A(n_2830),
.B(n_2435),
.Y(n_3045)
);

INVx3_ASAP7_75t_L g3046 ( 
.A(n_2653),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2846),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2783),
.Y(n_3048)
);

CKINVDCx16_ASAP7_75t_R g3049 ( 
.A(n_2680),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2670),
.Y(n_3050)
);

AND2x4_ASAP7_75t_L g3051 ( 
.A(n_2681),
.B(n_1473),
.Y(n_3051)
);

AND2x4_ASAP7_75t_L g3052 ( 
.A(n_2716),
.B(n_1487),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2670),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2708),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2708),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2710),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2710),
.Y(n_3057)
);

A2O1A1Ixp33_ASAP7_75t_L g3058 ( 
.A1(n_2698),
.A2(n_1615),
.B(n_1637),
.C(n_1612),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2867),
.B(n_2806),
.Y(n_3059)
);

AOI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2907),
.A2(n_2700),
.B(n_2676),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2928),
.A2(n_2717),
.B(n_2690),
.Y(n_3061)
);

OAI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2999),
.A2(n_2656),
.B(n_2627),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_3022),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2877),
.B(n_2889),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_3001),
.A2(n_2736),
.B(n_2724),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2882),
.B(n_2758),
.Y(n_3066)
);

OAI321xp33_ASAP7_75t_L g3067 ( 
.A1(n_2864),
.A2(n_2675),
.A3(n_2824),
.B1(n_1500),
.B2(n_1495),
.C(n_1504),
.Y(n_3067)
);

AOI21xp5_ASAP7_75t_L g3068 ( 
.A1(n_2968),
.A2(n_2719),
.B(n_2612),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2865),
.B(n_2651),
.Y(n_3069)
);

NOR3xp33_ASAP7_75t_L g3070 ( 
.A(n_2892),
.B(n_2844),
.C(n_2832),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2983),
.B(n_2682),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2915),
.B(n_2834),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2860),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2868),
.B(n_2834),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2937),
.B(n_2834),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2991),
.B(n_2811),
.Y(n_3076)
);

NOR2x1_ASAP7_75t_L g3077 ( 
.A(n_2939),
.B(n_2634),
.Y(n_3077)
);

INVxp67_ASAP7_75t_L g3078 ( 
.A(n_2903),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2861),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2924),
.A2(n_2791),
.B(n_2769),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2996),
.B(n_2811),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2893),
.B(n_2876),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_3007),
.B(n_2811),
.Y(n_3083)
);

OAI21xp33_ASAP7_75t_L g3084 ( 
.A1(n_3044),
.A2(n_2678),
.B(n_2657),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_3011),
.B(n_2904),
.Y(n_3085)
);

OAI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_3035),
.A2(n_2618),
.B(n_2804),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_2922),
.B(n_2651),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2886),
.B(n_2730),
.Y(n_3088)
);

NOR2x1_ASAP7_75t_L g3089 ( 
.A(n_3031),
.B(n_2683),
.Y(n_3089)
);

AOI22xp5_ASAP7_75t_L g3090 ( 
.A1(n_2859),
.A2(n_2784),
.B1(n_2699),
.B2(n_2733),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2984),
.A2(n_3028),
.B(n_2998),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2980),
.A2(n_2835),
.B(n_2785),
.Y(n_3092)
);

OAI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_3036),
.A2(n_2815),
.B(n_2778),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2975),
.A2(n_2756),
.B(n_2730),
.Y(n_3094)
);

OAI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_2952),
.A2(n_2671),
.B(n_1667),
.Y(n_3095)
);

A2O1A1Ixp33_ASAP7_75t_L g3096 ( 
.A1(n_2987),
.A2(n_1650),
.B(n_1713),
.C(n_1676),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2857),
.Y(n_3097)
);

INVxp67_ASAP7_75t_L g3098 ( 
.A(n_2895),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2888),
.B(n_2756),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_3029),
.Y(n_3100)
);

NAND2xp33_ASAP7_75t_L g3101 ( 
.A(n_3003),
.B(n_2780),
.Y(n_3101)
);

AOI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2932),
.A2(n_2688),
.B1(n_2817),
.B2(n_2788),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2960),
.B(n_1070),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_SL g3104 ( 
.A(n_3005),
.B(n_2780),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_3012),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2862),
.B(n_2788),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2863),
.B(n_2822),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2866),
.Y(n_3108)
);

AOI22xp5_ASAP7_75t_L g3109 ( 
.A1(n_3004),
.A2(n_2822),
.B1(n_1095),
.B2(n_1097),
.Y(n_3109)
);

AOI21x1_ASAP7_75t_L g3110 ( 
.A1(n_3042),
.A2(n_1733),
.B(n_1714),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2874),
.B(n_1195),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2995),
.A2(n_1623),
.B(n_1447),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2870),
.B(n_1093),
.Y(n_3113)
);

BUFx2_ASAP7_75t_L g3114 ( 
.A(n_2921),
.Y(n_3114)
);

AO32x1_ASAP7_75t_L g3115 ( 
.A1(n_3013),
.A2(n_1508),
.A3(n_1512),
.B1(n_1498),
.B2(n_1494),
.Y(n_3115)
);

O2A1O1Ixp5_ASAP7_75t_L g3116 ( 
.A1(n_3045),
.A2(n_1245),
.B(n_1274),
.C(n_1234),
.Y(n_3116)
);

OAI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2961),
.A2(n_1756),
.B(n_1518),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2954),
.B(n_1195),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_2926),
.B(n_1098),
.Y(n_3119)
);

INVxp67_ASAP7_75t_L g3120 ( 
.A(n_2949),
.Y(n_3120)
);

O2A1O1Ixp33_ASAP7_75t_L g3121 ( 
.A1(n_2923),
.A2(n_1514),
.B(n_1535),
.C(n_1521),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2881),
.A2(n_1109),
.B(n_1010),
.Y(n_3122)
);

INVx3_ASAP7_75t_L g3123 ( 
.A(n_2986),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2896),
.B(n_1110),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2897),
.B(n_1111),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2899),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2901),
.A2(n_1307),
.B(n_1147),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_2906),
.A2(n_1346),
.B(n_1341),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2910),
.A2(n_1721),
.B(n_1062),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_2911),
.A2(n_1078),
.B(n_1056),
.Y(n_3130)
);

OAI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_2912),
.A2(n_1120),
.B1(n_1125),
.B2(n_1114),
.Y(n_3131)
);

OAI22xp5_ASAP7_75t_L g3132 ( 
.A1(n_2916),
.A2(n_1134),
.B1(n_1140),
.B2(n_1137),
.Y(n_3132)
);

BUFx2_ASAP7_75t_SL g3133 ( 
.A(n_2909),
.Y(n_3133)
);

AOI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2917),
.A2(n_1085),
.B(n_1083),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2919),
.Y(n_3135)
);

AOI21xp5_ASAP7_75t_L g3136 ( 
.A1(n_2925),
.A2(n_1102),
.B(n_1086),
.Y(n_3136)
);

AOI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_2930),
.A2(n_2935),
.B(n_2934),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2940),
.A2(n_1112),
.B(n_1107),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2941),
.Y(n_3139)
);

OAI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_2963),
.A2(n_1548),
.B(n_1543),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2942),
.A2(n_1116),
.B(n_1115),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2943),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2945),
.A2(n_1118),
.B(n_1117),
.Y(n_3143)
);

NOR3xp33_ASAP7_75t_L g3144 ( 
.A(n_3020),
.B(n_1555),
.C(n_1550),
.Y(n_3144)
);

INVx3_ASAP7_75t_L g3145 ( 
.A(n_2990),
.Y(n_3145)
);

AOI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_2948),
.A2(n_1130),
.B(n_1121),
.Y(n_3146)
);

AOI21x1_ASAP7_75t_L g3147 ( 
.A1(n_3042),
.A2(n_1559),
.B(n_1556),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_2962),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2951),
.B(n_1157),
.Y(n_3149)
);

BUFx2_ASAP7_75t_L g3150 ( 
.A(n_2869),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_L g3151 ( 
.A1(n_3037),
.A2(n_1138),
.B(n_1131),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2884),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_2971),
.A2(n_1163),
.B1(n_1165),
.B2(n_1159),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2972),
.B(n_1171),
.Y(n_3154)
);

INVx3_ASAP7_75t_L g3155 ( 
.A(n_2900),
.Y(n_3155)
);

HB1xp67_ASAP7_75t_L g3156 ( 
.A(n_2920),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2978),
.A2(n_1149),
.B(n_1143),
.Y(n_3157)
);

CKINVDCx10_ASAP7_75t_R g3158 ( 
.A(n_3049),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2974),
.B(n_1176),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2981),
.B(n_2985),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2908),
.B(n_3025),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2887),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2989),
.A2(n_1180),
.B(n_1172),
.Y(n_3163)
);

NOR2xp33_ASAP7_75t_L g3164 ( 
.A(n_2967),
.B(n_1177),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_2872),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2992),
.A2(n_1183),
.B(n_1181),
.Y(n_3166)
);

O2A1O1Ixp33_ASAP7_75t_L g3167 ( 
.A1(n_2898),
.A2(n_1565),
.B(n_1568),
.C(n_1562),
.Y(n_3167)
);

OAI321xp33_ASAP7_75t_L g3168 ( 
.A1(n_2957),
.A2(n_1572),
.A3(n_1591),
.B1(n_1602),
.B2(n_1594),
.C(n_1578),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2879),
.B(n_1178),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2880),
.B(n_1188),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2875),
.B(n_1193),
.Y(n_3171)
);

OAI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_3018),
.A2(n_1608),
.B(n_1606),
.Y(n_3172)
);

O2A1O1Ixp33_ASAP7_75t_L g3173 ( 
.A1(n_2955),
.A2(n_1617),
.B(n_1618),
.C(n_1609),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_3023),
.B(n_1198),
.Y(n_3174)
);

AOI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_3032),
.A2(n_1191),
.B(n_1190),
.Y(n_3175)
);

A2O1A1Ixp33_ASAP7_75t_L g3176 ( 
.A1(n_3019),
.A2(n_1541),
.B(n_1563),
.C(n_1392),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2875),
.B(n_1206),
.Y(n_3177)
);

OAI22xp5_ASAP7_75t_L g3178 ( 
.A1(n_3027),
.A2(n_1212),
.B1(n_1215),
.B2(n_1210),
.Y(n_3178)
);

INVx2_ASAP7_75t_SL g3179 ( 
.A(n_2931),
.Y(n_3179)
);

A2O1A1Ixp33_ASAP7_75t_L g3180 ( 
.A1(n_3058),
.A2(n_1541),
.B(n_1563),
.C(n_1392),
.Y(n_3180)
);

OA21x2_ASAP7_75t_L g3181 ( 
.A1(n_3014),
.A2(n_1626),
.B(n_1620),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_SL g3182 ( 
.A(n_2956),
.B(n_1220),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_3038),
.B(n_1222),
.Y(n_3183)
);

INVx1_ASAP7_75t_SL g3184 ( 
.A(n_2936),
.Y(n_3184)
);

OR2x6_ASAP7_75t_L g3185 ( 
.A(n_2905),
.B(n_1742),
.Y(n_3185)
);

BUFx2_ASAP7_75t_L g3186 ( 
.A(n_3017),
.Y(n_3186)
);

AND2x4_ASAP7_75t_L g3187 ( 
.A(n_2950),
.B(n_1627),
.Y(n_3187)
);

AOI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2966),
.A2(n_1226),
.B1(n_1235),
.B2(n_1227),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_3041),
.A2(n_1209),
.B(n_1207),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_3043),
.A2(n_1225),
.B(n_1224),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_3033),
.A2(n_1241),
.B(n_1229),
.Y(n_3191)
);

A2O1A1Ixp33_ASAP7_75t_L g3192 ( 
.A1(n_3034),
.A2(n_1754),
.B(n_1742),
.C(n_1720),
.Y(n_3192)
);

AOI21x1_ASAP7_75t_L g3193 ( 
.A1(n_3053),
.A2(n_1647),
.B(n_1631),
.Y(n_3193)
);

AOI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_2894),
.A2(n_1251),
.B(n_1250),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_3016),
.B(n_1236),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_SL g3196 ( 
.A(n_3010),
.B(n_1240),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2959),
.B(n_1246),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3030),
.B(n_3024),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_L g3199 ( 
.A(n_2997),
.B(n_1258),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2927),
.B(n_1259),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2929),
.A2(n_1270),
.B(n_1268),
.Y(n_3201)
);

BUFx12f_ASAP7_75t_L g3202 ( 
.A(n_2871),
.Y(n_3202)
);

BUFx6f_ASAP7_75t_L g3203 ( 
.A(n_3021),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_2938),
.A2(n_1282),
.B(n_1279),
.Y(n_3204)
);

BUFx12f_ASAP7_75t_L g3205 ( 
.A(n_2918),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2944),
.B(n_1260),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2994),
.Y(n_3207)
);

OAI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_2947),
.A2(n_2964),
.B(n_2953),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_2970),
.A2(n_1297),
.B(n_1286),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3073),
.Y(n_3210)
);

BUFx10_ASAP7_75t_L g3211 ( 
.A(n_3087),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_3059),
.B(n_3064),
.Y(n_3212)
);

AOI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_3060),
.A2(n_2946),
.B(n_3054),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_3063),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_L g3215 ( 
.A(n_3161),
.B(n_2973),
.Y(n_3215)
);

AOI22xp33_ASAP7_75t_L g3216 ( 
.A1(n_3198),
.A2(n_2883),
.B1(n_2933),
.B2(n_2873),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_R g3217 ( 
.A(n_3158),
.B(n_2958),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3071),
.B(n_3103),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_3080),
.A2(n_3057),
.B(n_3055),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_3098),
.B(n_3030),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3079),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_3100),
.Y(n_3222)
);

OR2x6_ASAP7_75t_SL g3223 ( 
.A(n_3088),
.B(n_2979),
.Y(n_3223)
);

AOI21x1_ASAP7_75t_L g3224 ( 
.A1(n_3068),
.A2(n_3047),
.B(n_3040),
.Y(n_3224)
);

OAI21x1_ASAP7_75t_L g3225 ( 
.A1(n_3091),
.A2(n_2988),
.B(n_2982),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_3061),
.A2(n_3056),
.B(n_3050),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3085),
.B(n_3078),
.Y(n_3227)
);

BUFx6f_ASAP7_75t_L g3228 ( 
.A(n_3097),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_3065),
.A2(n_2993),
.B(n_2976),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3108),
.Y(n_3230)
);

OAI22xp5_ASAP7_75t_L g3231 ( 
.A1(n_3082),
.A2(n_2902),
.B1(n_2965),
.B2(n_2891),
.Y(n_3231)
);

NOR3xp33_ASAP7_75t_L g3232 ( 
.A(n_3144),
.B(n_1747),
.C(n_1693),
.Y(n_3232)
);

O2A1O1Ixp5_ASAP7_75t_L g3233 ( 
.A1(n_3116),
.A2(n_3026),
.B(n_3006),
.C(n_3051),
.Y(n_3233)
);

CKINVDCx11_ASAP7_75t_R g3234 ( 
.A(n_3205),
.Y(n_3234)
);

BUFx6f_ASAP7_75t_L g3235 ( 
.A(n_3097),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_3072),
.B(n_3074),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_3087),
.Y(n_3237)
);

INVx8_ASAP7_75t_L g3238 ( 
.A(n_3202),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3062),
.A2(n_3009),
.B(n_3002),
.Y(n_3239)
);

OAI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_3120),
.A2(n_2969),
.B1(n_3052),
.B2(n_2858),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_SL g3241 ( 
.A(n_3095),
.B(n_2913),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3075),
.A2(n_3048),
.B(n_3015),
.Y(n_3242)
);

OAI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_3067),
.A2(n_3039),
.B1(n_3000),
.B2(n_3046),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3137),
.A2(n_2890),
.B(n_2977),
.Y(n_3244)
);

NOR2xp33_ASAP7_75t_SL g3245 ( 
.A(n_3184),
.B(n_2878),
.Y(n_3245)
);

BUFx8_ASAP7_75t_SL g3246 ( 
.A(n_3123),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3160),
.B(n_3111),
.Y(n_3247)
);

NOR2xp33_ASAP7_75t_L g3248 ( 
.A(n_3114),
.B(n_3008),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3164),
.B(n_2883),
.Y(n_3249)
);

INVx2_ASAP7_75t_SL g3250 ( 
.A(n_3097),
.Y(n_3250)
);

OAI22xp5_ASAP7_75t_L g3251 ( 
.A1(n_3084),
.A2(n_2890),
.B1(n_2914),
.B2(n_2933),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3140),
.B(n_1261),
.Y(n_3252)
);

OAI21xp33_ASAP7_75t_L g3253 ( 
.A1(n_3117),
.A2(n_3199),
.B(n_3172),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3066),
.A2(n_1754),
.B(n_1168),
.Y(n_3254)
);

AOI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_3092),
.A2(n_1168),
.B(n_1073),
.Y(n_3255)
);

BUFx6f_ASAP7_75t_L g3256 ( 
.A(n_3203),
.Y(n_3256)
);

NOR3xp33_ASAP7_75t_SL g3257 ( 
.A(n_3197),
.B(n_1271),
.C(n_1262),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_3099),
.B(n_2885),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3105),
.Y(n_3259)
);

BUFx2_ASAP7_75t_L g3260 ( 
.A(n_3156),
.Y(n_3260)
);

A2O1A1Ixp33_ASAP7_75t_SL g3261 ( 
.A1(n_3070),
.A2(n_3155),
.B(n_3167),
.C(n_3166),
.Y(n_3261)
);

O2A1O1Ixp33_ASAP7_75t_L g3262 ( 
.A1(n_3121),
.A2(n_1670),
.B(n_1688),
.C(n_1665),
.Y(n_3262)
);

OAI22xp5_ASAP7_75t_L g3263 ( 
.A1(n_3113),
.A2(n_1277),
.B1(n_1285),
.B2(n_1284),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3126),
.B(n_1281),
.Y(n_3264)
);

O2A1O1Ixp33_ASAP7_75t_L g3265 ( 
.A1(n_3173),
.A2(n_1692),
.B(n_1699),
.C(n_1690),
.Y(n_3265)
);

NOR2xp33_ASAP7_75t_L g3266 ( 
.A(n_3179),
.B(n_3165),
.Y(n_3266)
);

AOI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3090),
.A2(n_1293),
.B1(n_1303),
.B2(n_1292),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3152),
.Y(n_3268)
);

INVx1_ASAP7_75t_SL g3269 ( 
.A(n_3150),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3162),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_L g3271 ( 
.A1(n_3170),
.A2(n_1214),
.B1(n_1573),
.B2(n_1228),
.Y(n_3271)
);

AOI33xp33_ASAP7_75t_L g3272 ( 
.A1(n_3188),
.A2(n_1722),
.A3(n_1707),
.B1(n_1725),
.B2(n_1719),
.B3(n_1703),
.Y(n_3272)
);

BUFx6f_ASAP7_75t_L g3273 ( 
.A(n_3203),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_3086),
.A2(n_3081),
.B(n_3076),
.Y(n_3274)
);

AND2x4_ASAP7_75t_L g3275 ( 
.A(n_3089),
.B(n_1726),
.Y(n_3275)
);

AOI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_3083),
.A2(n_1168),
.B(n_1073),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_L g3277 ( 
.A1(n_3187),
.A2(n_1214),
.B1(n_1573),
.B2(n_1228),
.Y(n_3277)
);

NOR2xp33_ASAP7_75t_L g3278 ( 
.A(n_3186),
.B(n_1305),
.Y(n_3278)
);

INVx3_ASAP7_75t_L g3279 ( 
.A(n_3203),
.Y(n_3279)
);

BUFx2_ASAP7_75t_L g3280 ( 
.A(n_3185),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_3135),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_3102),
.B(n_1505),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_3094),
.A2(n_3112),
.B(n_3093),
.Y(n_3283)
);

OR2x6_ASAP7_75t_L g3284 ( 
.A(n_3133),
.B(n_1683),
.Y(n_3284)
);

O2A1O1Ixp33_ASAP7_75t_L g3285 ( 
.A1(n_3096),
.A2(n_1737),
.B(n_1750),
.C(n_1734),
.Y(n_3285)
);

CKINVDCx11_ASAP7_75t_R g3286 ( 
.A(n_3185),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_3106),
.A2(n_3107),
.B(n_3139),
.Y(n_3287)
);

AO22x1_ASAP7_75t_L g3288 ( 
.A1(n_3145),
.A2(n_1318),
.B1(n_1451),
.B2(n_1374),
.Y(n_3288)
);

O2A1O1Ixp33_ASAP7_75t_L g3289 ( 
.A1(n_3168),
.A2(n_1757),
.B(n_1759),
.C(n_1751),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_3207),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3142),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3104),
.A2(n_1218),
.B(n_1168),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_3181),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3118),
.B(n_1323),
.Y(n_3294)
);

BUFx12f_ASAP7_75t_L g3295 ( 
.A(n_3187),
.Y(n_3295)
);

OAI22xp5_ASAP7_75t_L g3296 ( 
.A1(n_3124),
.A2(n_1353),
.B1(n_1356),
.B2(n_1327),
.Y(n_3296)
);

CKINVDCx8_ASAP7_75t_R g3297 ( 
.A(n_3181),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3193),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_3175),
.A2(n_1243),
.B(n_1218),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3101),
.B(n_1364),
.Y(n_3300)
);

INVxp67_ASAP7_75t_L g3301 ( 
.A(n_3069),
.Y(n_3301)
);

A2O1A1Ixp33_ASAP7_75t_SL g3302 ( 
.A1(n_3163),
.A2(n_1768),
.B(n_1765),
.C(n_1369),
.Y(n_3302)
);

A2O1A1Ixp33_ASAP7_75t_L g3303 ( 
.A1(n_3129),
.A2(n_1720),
.B(n_1696),
.C(n_1370),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3077),
.B(n_1371),
.Y(n_3304)
);

BUFx6f_ASAP7_75t_L g3305 ( 
.A(n_3148),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3208),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3200),
.Y(n_3307)
);

BUFx2_ASAP7_75t_L g3308 ( 
.A(n_3169),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3147),
.Y(n_3309)
);

BUFx2_ASAP7_75t_L g3310 ( 
.A(n_3109),
.Y(n_3310)
);

CKINVDCx16_ASAP7_75t_R g3311 ( 
.A(n_3131),
.Y(n_3311)
);

OAI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_3125),
.A2(n_1375),
.B1(n_1376),
.B2(n_1373),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3206),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3151),
.A2(n_1243),
.B(n_1218),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3149),
.Y(n_3315)
);

OAI21xp5_ASAP7_75t_L g3316 ( 
.A1(n_3130),
.A2(n_1384),
.B(n_1382),
.Y(n_3316)
);

O2A1O1Ixp33_ASAP7_75t_L g3317 ( 
.A1(n_3132),
.A2(n_1630),
.B(n_1705),
.C(n_1652),
.Y(n_3317)
);

AOI21xp5_ASAP7_75t_L g3318 ( 
.A1(n_3191),
.A2(n_3201),
.B(n_3194),
.Y(n_3318)
);

BUFx6f_ASAP7_75t_SL g3319 ( 
.A(n_3195),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3110),
.Y(n_3320)
);

AO32x2_ASAP7_75t_L g3321 ( 
.A1(n_3153),
.A2(n_1652),
.A3(n_1746),
.B1(n_1705),
.B2(n_1630),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3154),
.A2(n_1385),
.B1(n_1402),
.B2(n_1399),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_R g3323 ( 
.A(n_3183),
.B(n_1746),
.Y(n_3323)
);

OR2x6_ASAP7_75t_L g3324 ( 
.A(n_3171),
.B(n_1368),
.Y(n_3324)
);

OAI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_3159),
.A2(n_1413),
.B1(n_1420),
.B2(n_1414),
.Y(n_3325)
);

BUFx2_ASAP7_75t_L g3326 ( 
.A(n_3174),
.Y(n_3326)
);

O2A1O1Ixp33_ASAP7_75t_L g3327 ( 
.A1(n_3178),
.A2(n_947),
.B(n_1422),
.C(n_1415),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3119),
.B(n_1425),
.Y(n_3328)
);

A2O1A1Ixp33_ASAP7_75t_L g3329 ( 
.A1(n_3122),
.A2(n_1427),
.B(n_1429),
.C(n_1428),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3182),
.B(n_1426),
.Y(n_3330)
);

INVx3_ASAP7_75t_L g3331 ( 
.A(n_3177),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3196),
.B(n_3134),
.Y(n_3332)
);

INVx1_ASAP7_75t_SL g3333 ( 
.A(n_3127),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3204),
.A2(n_1243),
.B(n_1218),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_SL g3335 ( 
.A(n_3136),
.B(n_1524),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_3192),
.Y(n_3336)
);

O2A1O1Ixp33_ASAP7_75t_L g3337 ( 
.A1(n_3176),
.A2(n_1431),
.B(n_1436),
.C(n_1430),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3180),
.B(n_1437),
.Y(n_3338)
);

OAI21xp33_ASAP7_75t_SL g3339 ( 
.A1(n_3138),
.A2(n_0),
.B(n_3),
.Y(n_3339)
);

O2A1O1Ixp5_ASAP7_75t_L g3340 ( 
.A1(n_3157),
.A2(n_1423),
.B(n_1424),
.C(n_1368),
.Y(n_3340)
);

INVx6_ASAP7_75t_L g3341 ( 
.A(n_3128),
.Y(n_3341)
);

BUFx6f_ASAP7_75t_L g3342 ( 
.A(n_3115),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3115),
.Y(n_3343)
);

OAI21x1_ASAP7_75t_L g3344 ( 
.A1(n_3209),
.A2(n_1475),
.B(n_1406),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_3141),
.B(n_1524),
.Y(n_3345)
);

HB1xp67_ASAP7_75t_L g3346 ( 
.A(n_3143),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3146),
.B(n_1445),
.Y(n_3347)
);

NOR2x1_ASAP7_75t_L g3348 ( 
.A(n_3189),
.B(n_2025),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3190),
.Y(n_3349)
);

BUFx6f_ASAP7_75t_L g3350 ( 
.A(n_3228),
.Y(n_3350)
);

INVx1_ASAP7_75t_SL g3351 ( 
.A(n_3286),
.Y(n_3351)
);

INVx1_ASAP7_75t_SL g3352 ( 
.A(n_3269),
.Y(n_3352)
);

NAND2x1p5_ASAP7_75t_L g3353 ( 
.A(n_3228),
.B(n_2025),
.Y(n_3353)
);

BUFx4f_ASAP7_75t_L g3354 ( 
.A(n_3238),
.Y(n_3354)
);

INVx1_ASAP7_75t_SL g3355 ( 
.A(n_3217),
.Y(n_3355)
);

CKINVDCx5p33_ASAP7_75t_R g3356 ( 
.A(n_3234),
.Y(n_3356)
);

INVxp67_ASAP7_75t_SL g3357 ( 
.A(n_3227),
.Y(n_3357)
);

INVx5_ASAP7_75t_L g3358 ( 
.A(n_3235),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3212),
.B(n_1446),
.Y(n_3359)
);

BUFx2_ASAP7_75t_SL g3360 ( 
.A(n_3319),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3281),
.Y(n_3361)
);

BUFx3_ASAP7_75t_L g3362 ( 
.A(n_3235),
.Y(n_3362)
);

BUFx2_ASAP7_75t_L g3363 ( 
.A(n_3260),
.Y(n_3363)
);

INVx2_ASAP7_75t_SL g3364 ( 
.A(n_3256),
.Y(n_3364)
);

BUFx5_ASAP7_75t_L g3365 ( 
.A(n_3349),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3259),
.Y(n_3366)
);

BUFx4_ASAP7_75t_SL g3367 ( 
.A(n_3284),
.Y(n_3367)
);

NAND2x1p5_ASAP7_75t_L g3368 ( 
.A(n_3256),
.B(n_2032),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3218),
.B(n_1450),
.Y(n_3369)
);

BUFx2_ASAP7_75t_L g3370 ( 
.A(n_3279),
.Y(n_3370)
);

AOI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_3253),
.A2(n_3311),
.B1(n_3215),
.B2(n_3310),
.Y(n_3371)
);

INVx3_ASAP7_75t_L g3372 ( 
.A(n_3273),
.Y(n_3372)
);

BUFx6f_ASAP7_75t_L g3373 ( 
.A(n_3273),
.Y(n_3373)
);

INVx3_ASAP7_75t_L g3374 ( 
.A(n_3211),
.Y(n_3374)
);

BUFx3_ASAP7_75t_L g3375 ( 
.A(n_3305),
.Y(n_3375)
);

CKINVDCx11_ASAP7_75t_R g3376 ( 
.A(n_3238),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3291),
.Y(n_3377)
);

INVx3_ASAP7_75t_L g3378 ( 
.A(n_3237),
.Y(n_3378)
);

INVx2_ASAP7_75t_SL g3379 ( 
.A(n_3250),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3210),
.Y(n_3380)
);

BUFx3_ASAP7_75t_L g3381 ( 
.A(n_3305),
.Y(n_3381)
);

BUFx3_ASAP7_75t_L g3382 ( 
.A(n_3295),
.Y(n_3382)
);

BUFx3_ASAP7_75t_L g3383 ( 
.A(n_3290),
.Y(n_3383)
);

BUFx3_ASAP7_75t_L g3384 ( 
.A(n_3246),
.Y(n_3384)
);

BUFx2_ASAP7_75t_L g3385 ( 
.A(n_3284),
.Y(n_3385)
);

INVx6_ASAP7_75t_L g3386 ( 
.A(n_3275),
.Y(n_3386)
);

BUFx4f_ASAP7_75t_SL g3387 ( 
.A(n_3331),
.Y(n_3387)
);

INVx1_ASAP7_75t_SL g3388 ( 
.A(n_3280),
.Y(n_3388)
);

BUFx3_ASAP7_75t_L g3389 ( 
.A(n_3266),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3221),
.Y(n_3390)
);

BUFx12f_ASAP7_75t_L g3391 ( 
.A(n_3326),
.Y(n_3391)
);

INVx1_ASAP7_75t_SL g3392 ( 
.A(n_3245),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3230),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3214),
.Y(n_3394)
);

INVx4_ASAP7_75t_L g3395 ( 
.A(n_3324),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3222),
.Y(n_3396)
);

INVx2_ASAP7_75t_SL g3397 ( 
.A(n_3323),
.Y(n_3397)
);

INVx1_ASAP7_75t_SL g3398 ( 
.A(n_3223),
.Y(n_3398)
);

BUFx2_ASAP7_75t_L g3399 ( 
.A(n_3247),
.Y(n_3399)
);

HB1xp67_ASAP7_75t_L g3400 ( 
.A(n_3220),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3268),
.Y(n_3401)
);

BUFx10_ASAP7_75t_L g3402 ( 
.A(n_3248),
.Y(n_3402)
);

INVx5_ASAP7_75t_L g3403 ( 
.A(n_3324),
.Y(n_3403)
);

INVx6_ASAP7_75t_SL g3404 ( 
.A(n_3240),
.Y(n_3404)
);

BUFx2_ASAP7_75t_L g3405 ( 
.A(n_3301),
.Y(n_3405)
);

HB1xp67_ASAP7_75t_L g3406 ( 
.A(n_3287),
.Y(n_3406)
);

INVx5_ASAP7_75t_L g3407 ( 
.A(n_3308),
.Y(n_3407)
);

INVx4_ASAP7_75t_L g3408 ( 
.A(n_3341),
.Y(n_3408)
);

INVx5_ASAP7_75t_L g3409 ( 
.A(n_3342),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3270),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3307),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3315),
.B(n_1455),
.Y(n_3412)
);

BUFx3_ASAP7_75t_L g3413 ( 
.A(n_3258),
.Y(n_3413)
);

INVx1_ASAP7_75t_SL g3414 ( 
.A(n_3249),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3306),
.Y(n_3415)
);

BUFx5_ASAP7_75t_L g3416 ( 
.A(n_3313),
.Y(n_3416)
);

BUFx2_ASAP7_75t_L g3417 ( 
.A(n_3231),
.Y(n_3417)
);

INVx2_ASAP7_75t_SL g3418 ( 
.A(n_3241),
.Y(n_3418)
);

BUFx6f_ASAP7_75t_L g3419 ( 
.A(n_3304),
.Y(n_3419)
);

BUFx4_ASAP7_75t_SL g3420 ( 
.A(n_3343),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3298),
.Y(n_3421)
);

BUFx3_ASAP7_75t_L g3422 ( 
.A(n_3278),
.Y(n_3422)
);

INVx4_ASAP7_75t_L g3423 ( 
.A(n_3338),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3272),
.B(n_3243),
.Y(n_3424)
);

INVx2_ASAP7_75t_SL g3425 ( 
.A(n_3282),
.Y(n_3425)
);

BUFx6f_ASAP7_75t_L g3426 ( 
.A(n_3300),
.Y(n_3426)
);

BUFx3_ASAP7_75t_L g3427 ( 
.A(n_3225),
.Y(n_3427)
);

NAND2x1p5_ASAP7_75t_L g3428 ( 
.A(n_3348),
.B(n_2032),
.Y(n_3428)
);

BUFx6f_ASAP7_75t_L g3429 ( 
.A(n_3294),
.Y(n_3429)
);

INVxp67_ASAP7_75t_SL g3430 ( 
.A(n_3239),
.Y(n_3430)
);

INVx3_ASAP7_75t_L g3431 ( 
.A(n_3336),
.Y(n_3431)
);

BUFx2_ASAP7_75t_L g3432 ( 
.A(n_3346),
.Y(n_3432)
);

INVx2_ASAP7_75t_SL g3433 ( 
.A(n_3288),
.Y(n_3433)
);

INVxp67_ASAP7_75t_SL g3434 ( 
.A(n_3309),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3293),
.Y(n_3435)
);

INVx1_ASAP7_75t_SL g3436 ( 
.A(n_3244),
.Y(n_3436)
);

BUFx3_ASAP7_75t_L g3437 ( 
.A(n_3264),
.Y(n_3437)
);

NAND2x1p5_ASAP7_75t_L g3438 ( 
.A(n_3236),
.B(n_2156),
.Y(n_3438)
);

BUFx3_ASAP7_75t_L g3439 ( 
.A(n_3330),
.Y(n_3439)
);

BUFx6f_ASAP7_75t_L g3440 ( 
.A(n_3321),
.Y(n_3440)
);

INVx4_ASAP7_75t_L g3441 ( 
.A(n_3342),
.Y(n_3441)
);

BUFx2_ASAP7_75t_SL g3442 ( 
.A(n_3242),
.Y(n_3442)
);

BUFx6f_ASAP7_75t_L g3443 ( 
.A(n_3321),
.Y(n_3443)
);

INVx2_ASAP7_75t_SL g3444 ( 
.A(n_3328),
.Y(n_3444)
);

INVx3_ASAP7_75t_L g3445 ( 
.A(n_3224),
.Y(n_3445)
);

NAND2x1p5_ASAP7_75t_L g3446 ( 
.A(n_3335),
.B(n_3345),
.Y(n_3446)
);

AND2x4_ASAP7_75t_L g3447 ( 
.A(n_3257),
.B(n_2156),
.Y(n_3447)
);

BUFx3_ASAP7_75t_L g3448 ( 
.A(n_3332),
.Y(n_3448)
);

INVx2_ASAP7_75t_SL g3449 ( 
.A(n_3251),
.Y(n_3449)
);

NAND2x1p5_ASAP7_75t_L g3450 ( 
.A(n_3333),
.B(n_2165),
.Y(n_3450)
);

BUFx6f_ASAP7_75t_L g3451 ( 
.A(n_3297),
.Y(n_3451)
);

NAND2x1p5_ASAP7_75t_L g3452 ( 
.A(n_3213),
.B(n_2165),
.Y(n_3452)
);

INVx1_ASAP7_75t_SL g3453 ( 
.A(n_3347),
.Y(n_3453)
);

CKINVDCx20_ASAP7_75t_R g3454 ( 
.A(n_3267),
.Y(n_3454)
);

BUFx3_ASAP7_75t_L g3455 ( 
.A(n_3320),
.Y(n_3455)
);

INVx3_ASAP7_75t_SL g3456 ( 
.A(n_3261),
.Y(n_3456)
);

BUFx8_ASAP7_75t_L g3457 ( 
.A(n_3277),
.Y(n_3457)
);

INVx3_ASAP7_75t_L g3458 ( 
.A(n_3344),
.Y(n_3458)
);

INVx4_ASAP7_75t_L g3459 ( 
.A(n_3233),
.Y(n_3459)
);

NAND2x1p5_ASAP7_75t_L g3460 ( 
.A(n_3219),
.B(n_2177),
.Y(n_3460)
);

OAI21x1_ASAP7_75t_L g3461 ( 
.A1(n_3452),
.A2(n_3255),
.B(n_3283),
.Y(n_3461)
);

INVx4_ASAP7_75t_L g3462 ( 
.A(n_3354),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3366),
.Y(n_3463)
);

OAI211xp5_ASAP7_75t_SL g3464 ( 
.A1(n_3359),
.A2(n_3316),
.B(n_3317),
.C(n_3339),
.Y(n_3464)
);

HB1xp67_ASAP7_75t_L g3465 ( 
.A(n_3432),
.Y(n_3465)
);

INVxp67_ASAP7_75t_L g3466 ( 
.A(n_3389),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_3363),
.B(n_3216),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3380),
.Y(n_3468)
);

AOI21x1_ASAP7_75t_L g3469 ( 
.A1(n_3406),
.A2(n_3254),
.B(n_3274),
.Y(n_3469)
);

HB1xp67_ASAP7_75t_L g3470 ( 
.A(n_3357),
.Y(n_3470)
);

CKINVDCx8_ASAP7_75t_R g3471 ( 
.A(n_3360),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3390),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3422),
.B(n_1460),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3399),
.B(n_3232),
.Y(n_3474)
);

INVx3_ASAP7_75t_L g3475 ( 
.A(n_3350),
.Y(n_3475)
);

AO21x2_ASAP7_75t_L g3476 ( 
.A1(n_3421),
.A2(n_3276),
.B(n_3226),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_SL g3477 ( 
.A(n_3371),
.B(n_3252),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3393),
.Y(n_3478)
);

NOR2xp67_ASAP7_75t_L g3479 ( 
.A(n_3407),
.B(n_3292),
.Y(n_3479)
);

AOI221xp5_ASAP7_75t_L g3480 ( 
.A1(n_3424),
.A2(n_3262),
.B1(n_3265),
.B2(n_3312),
.C(n_3289),
.Y(n_3480)
);

BUFx6f_ASAP7_75t_L g3481 ( 
.A(n_3373),
.Y(n_3481)
);

BUFx8_ASAP7_75t_L g3482 ( 
.A(n_3384),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_3387),
.B(n_1461),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3361),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3377),
.Y(n_3485)
);

OR2x6_ASAP7_75t_L g3486 ( 
.A(n_3386),
.B(n_3327),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3411),
.B(n_1464),
.Y(n_3487)
);

OAI21x1_ASAP7_75t_L g3488 ( 
.A1(n_3460),
.A2(n_3229),
.B(n_3340),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3400),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3415),
.Y(n_3490)
);

INVx3_ASAP7_75t_L g3491 ( 
.A(n_3362),
.Y(n_3491)
);

INVxp67_ASAP7_75t_L g3492 ( 
.A(n_3437),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3449),
.A2(n_3271),
.B1(n_1595),
.B2(n_3318),
.Y(n_3493)
);

AND2x4_ASAP7_75t_L g3494 ( 
.A(n_3407),
.B(n_3303),
.Y(n_3494)
);

AO31x2_ASAP7_75t_L g3495 ( 
.A1(n_3459),
.A2(n_3334),
.A3(n_3299),
.B(n_3314),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3394),
.Y(n_3496)
);

BUFx3_ASAP7_75t_L g3497 ( 
.A(n_3375),
.Y(n_3497)
);

OAI21x1_ASAP7_75t_L g3498 ( 
.A1(n_3458),
.A2(n_3337),
.B(n_3285),
.Y(n_3498)
);

OAI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3412),
.A2(n_3329),
.B(n_3296),
.Y(n_3499)
);

OAI21x1_ASAP7_75t_L g3500 ( 
.A1(n_3445),
.A2(n_3322),
.B(n_3263),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3396),
.Y(n_3501)
);

AO21x2_ASAP7_75t_L g3502 ( 
.A1(n_3434),
.A2(n_3302),
.B(n_3325),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3401),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3352),
.B(n_1466),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3440),
.B(n_1423),
.Y(n_3505)
);

AO21x2_ASAP7_75t_L g3506 ( 
.A1(n_3430),
.A2(n_1595),
.B(n_1475),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_3417),
.A2(n_1424),
.B(n_1423),
.Y(n_3507)
);

CKINVDCx5p33_ASAP7_75t_R g3508 ( 
.A(n_3376),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3453),
.A2(n_1424),
.B1(n_1576),
.B2(n_1423),
.Y(n_3509)
);

BUFx12f_ASAP7_75t_L g3510 ( 
.A(n_3356),
.Y(n_3510)
);

OAI22xp5_ASAP7_75t_L g3511 ( 
.A1(n_3454),
.A2(n_1485),
.B1(n_1509),
.B2(n_1474),
.Y(n_3511)
);

OR2x2_ASAP7_75t_L g3512 ( 
.A(n_3414),
.B(n_1424),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3410),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3435),
.Y(n_3514)
);

BUFx10_ASAP7_75t_L g3515 ( 
.A(n_3397),
.Y(n_3515)
);

OAI21x1_ASAP7_75t_L g3516 ( 
.A1(n_3450),
.A2(n_1475),
.B(n_1406),
.Y(n_3516)
);

OR2x6_ASAP7_75t_L g3517 ( 
.A(n_3391),
.B(n_1576),
.Y(n_3517)
);

AOI21x1_ASAP7_75t_L g3518 ( 
.A1(n_3405),
.A2(n_2189),
.B(n_2177),
.Y(n_3518)
);

AND2x6_ASAP7_75t_L g3519 ( 
.A(n_3436),
.B(n_1576),
.Y(n_3519)
);

OA21x2_ASAP7_75t_L g3520 ( 
.A1(n_3398),
.A2(n_1469),
.B(n_1468),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3455),
.Y(n_3521)
);

OR2x6_ASAP7_75t_L g3522 ( 
.A(n_3382),
.B(n_1576),
.Y(n_3522)
);

CKINVDCx6p67_ASAP7_75t_R g3523 ( 
.A(n_3355),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3443),
.A2(n_1701),
.B1(n_1472),
.B2(n_1477),
.Y(n_3524)
);

AOI22xp5_ASAP7_75t_L g3525 ( 
.A1(n_3433),
.A2(n_1478),
.B1(n_1479),
.B2(n_1471),
.Y(n_3525)
);

OAI21xp5_ASAP7_75t_SL g3526 ( 
.A1(n_3351),
.A2(n_1701),
.B(n_0),
.Y(n_3526)
);

OAI21x1_ASAP7_75t_L g3527 ( 
.A1(n_3428),
.A2(n_1475),
.B(n_1406),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3416),
.Y(n_3528)
);

AND2x4_ASAP7_75t_L g3529 ( 
.A(n_3388),
.B(n_2189),
.Y(n_3529)
);

AOI22x1_ASAP7_75t_L g3530 ( 
.A1(n_3456),
.A2(n_1490),
.B1(n_1497),
.B2(n_1481),
.Y(n_3530)
);

INVx8_ASAP7_75t_L g3531 ( 
.A(n_3358),
.Y(n_3531)
);

OAI21x1_ASAP7_75t_L g3532 ( 
.A1(n_3431),
.A2(n_1475),
.B(n_1406),
.Y(n_3532)
);

OR2x2_ASAP7_75t_L g3533 ( 
.A(n_3413),
.B(n_1701),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3448),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3416),
.Y(n_3535)
);

INVx4_ASAP7_75t_L g3536 ( 
.A(n_3358),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3465),
.B(n_3383),
.Y(n_3537)
);

AOI22xp33_ASAP7_75t_L g3538 ( 
.A1(n_3477),
.A2(n_3429),
.B1(n_3419),
.B2(n_3423),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3501),
.Y(n_3539)
);

HB1xp67_ASAP7_75t_L g3540 ( 
.A(n_3470),
.Y(n_3540)
);

INVx3_ASAP7_75t_L g3541 ( 
.A(n_3531),
.Y(n_3541)
);

OA21x2_ASAP7_75t_L g3542 ( 
.A1(n_3532),
.A2(n_3370),
.B(n_3385),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3484),
.Y(n_3543)
);

BUFx3_ASAP7_75t_L g3544 ( 
.A(n_3497),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3466),
.B(n_3402),
.Y(n_3545)
);

INVx2_ASAP7_75t_SL g3546 ( 
.A(n_3491),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_3485),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3490),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_SL g3549 ( 
.A1(n_3519),
.A2(n_3442),
.B1(n_3403),
.B2(n_3457),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3489),
.Y(n_3550)
);

CKINVDCx5p33_ASAP7_75t_R g3551 ( 
.A(n_3508),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3468),
.Y(n_3552)
);

CKINVDCx11_ASAP7_75t_R g3553 ( 
.A(n_3471),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_L g3554 ( 
.A1(n_3480),
.A2(n_3404),
.B1(n_3426),
.B2(n_3439),
.Y(n_3554)
);

INVx3_ASAP7_75t_L g3555 ( 
.A(n_3531),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3472),
.Y(n_3556)
);

BUFx4f_ASAP7_75t_L g3557 ( 
.A(n_3523),
.Y(n_3557)
);

HB1xp67_ASAP7_75t_L g3558 ( 
.A(n_3534),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3496),
.Y(n_3559)
);

BUFx3_ASAP7_75t_L g3560 ( 
.A(n_3482),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3478),
.Y(n_3561)
);

INVx3_ASAP7_75t_L g3562 ( 
.A(n_3536),
.Y(n_3562)
);

INVxp67_ASAP7_75t_SL g3563 ( 
.A(n_3535),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3503),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3513),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3514),
.Y(n_3566)
);

HB1xp67_ASAP7_75t_L g3567 ( 
.A(n_3521),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_3463),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3505),
.Y(n_3569)
);

OAI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_3526),
.A2(n_3403),
.B1(n_3395),
.B2(n_3418),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3512),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3528),
.Y(n_3572)
);

AOI21x1_ASAP7_75t_L g3573 ( 
.A1(n_3518),
.A2(n_3447),
.B(n_3369),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3467),
.B(n_3381),
.Y(n_3574)
);

AOI22xp33_ASAP7_75t_L g3575 ( 
.A1(n_3464),
.A2(n_3444),
.B1(n_3392),
.B2(n_3451),
.Y(n_3575)
);

AND2x4_ASAP7_75t_L g3576 ( 
.A(n_3492),
.B(n_3408),
.Y(n_3576)
);

INVx3_ASAP7_75t_L g3577 ( 
.A(n_3481),
.Y(n_3577)
);

INVx2_ASAP7_75t_SL g3578 ( 
.A(n_3481),
.Y(n_3578)
);

BUFx2_ASAP7_75t_L g3579 ( 
.A(n_3461),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3533),
.Y(n_3580)
);

HB1xp67_ASAP7_75t_L g3581 ( 
.A(n_3474),
.Y(n_3581)
);

OAI21x1_ASAP7_75t_L g3582 ( 
.A1(n_3469),
.A2(n_3438),
.B(n_3446),
.Y(n_3582)
);

INVx5_ASAP7_75t_L g3583 ( 
.A(n_3519),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3476),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3506),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3529),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3519),
.Y(n_3587)
);

BUFx6f_ASAP7_75t_L g3588 ( 
.A(n_3515),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3487),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_3494),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3500),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3502),
.Y(n_3592)
);

OAI21xp5_ASAP7_75t_SL g3593 ( 
.A1(n_3499),
.A2(n_3420),
.B(n_3367),
.Y(n_3593)
);

NOR2x1p5_ASAP7_75t_L g3594 ( 
.A(n_3560),
.B(n_3510),
.Y(n_3594)
);

OAI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3593),
.A2(n_3493),
.B1(n_3524),
.B2(n_3509),
.Y(n_3595)
);

AND2x4_ASAP7_75t_L g3596 ( 
.A(n_3590),
.B(n_3409),
.Y(n_3596)
);

AND2x4_ASAP7_75t_L g3597 ( 
.A(n_3590),
.B(n_3409),
.Y(n_3597)
);

OR2x2_ASAP7_75t_L g3598 ( 
.A(n_3581),
.B(n_3441),
.Y(n_3598)
);

INVxp33_ASAP7_75t_SL g3599 ( 
.A(n_3551),
.Y(n_3599)
);

NAND2xp33_ASAP7_75t_SL g3600 ( 
.A(n_3588),
.B(n_3462),
.Y(n_3600)
);

AOI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3589),
.A2(n_3520),
.B1(n_3486),
.B2(n_3425),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3548),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3552),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3540),
.B(n_3475),
.Y(n_3604)
);

HB1xp67_ASAP7_75t_L g3605 ( 
.A(n_3558),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3543),
.Y(n_3606)
);

OAI22xp5_ASAP7_75t_L g3607 ( 
.A1(n_3570),
.A2(n_3525),
.B1(n_3473),
.B2(n_3507),
.Y(n_3607)
);

CKINVDCx20_ASAP7_75t_R g3608 ( 
.A(n_3553),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3550),
.B(n_3416),
.Y(n_3609)
);

NOR2xp33_ASAP7_75t_R g3610 ( 
.A(n_3557),
.B(n_3483),
.Y(n_3610)
);

CKINVDCx5p33_ASAP7_75t_R g3611 ( 
.A(n_3544),
.Y(n_3611)
);

NAND3xp33_ASAP7_75t_SL g3612 ( 
.A(n_3575),
.B(n_3538),
.C(n_3549),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3537),
.B(n_3365),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3547),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_SL g3615 ( 
.A1(n_3588),
.A2(n_3517),
.B1(n_3522),
.B2(n_3511),
.Y(n_3615)
);

XOR2x2_ASAP7_75t_SL g3616 ( 
.A(n_3576),
.B(n_3504),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3567),
.B(n_3545),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3559),
.Y(n_3618)
);

HB1xp67_ASAP7_75t_L g3619 ( 
.A(n_3556),
.Y(n_3619)
);

AND2x4_ASAP7_75t_L g3620 ( 
.A(n_3569),
.B(n_3378),
.Y(n_3620)
);

CKINVDCx14_ASAP7_75t_R g3621 ( 
.A(n_3574),
.Y(n_3621)
);

HB1xp67_ASAP7_75t_L g3622 ( 
.A(n_3561),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3565),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3564),
.Y(n_3624)
);

CKINVDCx5p33_ASAP7_75t_R g3625 ( 
.A(n_3588),
.Y(n_3625)
);

CKINVDCx16_ASAP7_75t_R g3626 ( 
.A(n_3576),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3566),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3563),
.B(n_3365),
.Y(n_3628)
);

NAND2xp33_ASAP7_75t_R g3629 ( 
.A(n_3541),
.B(n_3372),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3546),
.B(n_3365),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3572),
.B(n_3379),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3539),
.Y(n_3632)
);

INVx2_ASAP7_75t_SL g3633 ( 
.A(n_3578),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3568),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3580),
.Y(n_3635)
);

CKINVDCx5p33_ASAP7_75t_R g3636 ( 
.A(n_3577),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3562),
.B(n_3364),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3571),
.Y(n_3638)
);

BUFx12f_ASAP7_75t_L g3639 ( 
.A(n_3583),
.Y(n_3639)
);

INVx4_ASAP7_75t_L g3640 ( 
.A(n_3555),
.Y(n_3640)
);

OAI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_3582),
.A2(n_3530),
.B(n_3498),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3591),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3586),
.B(n_3427),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3587),
.B(n_1701),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3592),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_R g3646 ( 
.A(n_3554),
.B(n_3374),
.Y(n_3646)
);

NAND3xp33_ASAP7_75t_L g3647 ( 
.A(n_3584),
.B(n_3479),
.C(n_1502),
.Y(n_3647)
);

OAI222xp33_ASAP7_75t_L g3648 ( 
.A1(n_3583),
.A2(n_1522),
.B1(n_1510),
.B2(n_1525),
.C1(n_1520),
.C2(n_1501),
.Y(n_3648)
);

NOR3xp33_ASAP7_75t_SL g3649 ( 
.A(n_3579),
.B(n_1529),
.C(n_1527),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3585),
.Y(n_3650)
);

CKINVDCx8_ASAP7_75t_R g3651 ( 
.A(n_3583),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3579),
.B(n_3495),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3626),
.B(n_3542),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3645),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3617),
.B(n_3542),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3605),
.B(n_3573),
.Y(n_3656)
);

HB1xp67_ASAP7_75t_L g3657 ( 
.A(n_3619),
.Y(n_3657)
);

INVx1_ASAP7_75t_SL g3658 ( 
.A(n_3608),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3606),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3622),
.Y(n_3660)
);

NAND2x1p5_ASAP7_75t_L g3661 ( 
.A(n_3594),
.B(n_3573),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3614),
.Y(n_3662)
);

BUFx6f_ASAP7_75t_L g3663 ( 
.A(n_3639),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3602),
.Y(n_3664)
);

BUFx6f_ASAP7_75t_L g3665 ( 
.A(n_3625),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3635),
.B(n_3495),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3618),
.Y(n_3667)
);

INVx3_ASAP7_75t_L g3668 ( 
.A(n_3640),
.Y(n_3668)
);

HB1xp67_ASAP7_75t_L g3669 ( 
.A(n_3603),
.Y(n_3669)
);

OR2x6_ASAP7_75t_L g3670 ( 
.A(n_3596),
.B(n_3597),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3624),
.B(n_3488),
.Y(n_3671)
);

OAI22xp33_ASAP7_75t_L g3672 ( 
.A1(n_3607),
.A2(n_3368),
.B1(n_3353),
.B2(n_1531),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3627),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3623),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3604),
.B(n_3621),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3613),
.B(n_3516),
.Y(n_3676)
);

INVx3_ASAP7_75t_L g3677 ( 
.A(n_3611),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3598),
.B(n_3527),
.Y(n_3678)
);

OR2x6_ASAP7_75t_L g3679 ( 
.A(n_3596),
.B(n_1243),
.Y(n_3679)
);

AOI33xp33_ASAP7_75t_L g3680 ( 
.A1(n_3601),
.A2(n_1542),
.A3(n_1533),
.B1(n_1544),
.B2(n_1539),
.B3(n_1530),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3634),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3642),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3652),
.B(n_1406),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3597),
.B(n_3),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_3599),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3630),
.B(n_3633),
.Y(n_3686)
);

HB1xp67_ASAP7_75t_L g3687 ( 
.A(n_3657),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3682),
.Y(n_3688)
);

HB1xp67_ASAP7_75t_L g3689 ( 
.A(n_3656),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3670),
.B(n_3675),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3670),
.B(n_3637),
.Y(n_3691)
);

OAI21xp33_ASAP7_75t_L g3692 ( 
.A1(n_3655),
.A2(n_3609),
.B(n_3628),
.Y(n_3692)
);

AOI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_3683),
.A2(n_3600),
.B(n_3641),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3666),
.A2(n_3612),
.B(n_3644),
.Y(n_3694)
);

HB1xp67_ASAP7_75t_L g3695 ( 
.A(n_3669),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3660),
.Y(n_3696)
);

A2O1A1Ixp33_ASAP7_75t_L g3697 ( 
.A1(n_3653),
.A2(n_3649),
.B(n_3647),
.C(n_3595),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3664),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3674),
.A2(n_3678),
.B1(n_3662),
.B2(n_3667),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3673),
.Y(n_3700)
);

AOI221xp5_ASAP7_75t_L g3701 ( 
.A1(n_3672),
.A2(n_3648),
.B1(n_1554),
.B2(n_1564),
.C(n_1557),
.Y(n_3701)
);

BUFx3_ASAP7_75t_L g3702 ( 
.A(n_3665),
.Y(n_3702)
);

A2O1A1Ixp33_ASAP7_75t_L g3703 ( 
.A1(n_3680),
.A2(n_3616),
.B(n_3631),
.C(n_3643),
.Y(n_3703)
);

OAI211xp5_ASAP7_75t_L g3704 ( 
.A1(n_3684),
.A2(n_3610),
.B(n_3646),
.C(n_3651),
.Y(n_3704)
);

BUFx2_ASAP7_75t_L g3705 ( 
.A(n_3665),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3654),
.Y(n_3706)
);

OA21x2_ASAP7_75t_L g3707 ( 
.A1(n_3659),
.A2(n_3650),
.B(n_3632),
.Y(n_3707)
);

AO31x2_ASAP7_75t_L g3708 ( 
.A1(n_3681),
.A2(n_3638),
.A3(n_3661),
.B(n_3679),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3671),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3671),
.Y(n_3710)
);

AO31x2_ASAP7_75t_L g3711 ( 
.A1(n_3679),
.A2(n_3629),
.A3(n_3636),
.B(n_3615),
.Y(n_3711)
);

AO31x2_ASAP7_75t_L g3712 ( 
.A1(n_3663),
.A2(n_3620),
.A3(n_1475),
.B(n_1673),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3676),
.Y(n_3713)
);

AOI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3686),
.A2(n_1567),
.B1(n_1571),
.B2(n_1551),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3668),
.B(n_1406),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3663),
.Y(n_3716)
);

HB1xp67_ASAP7_75t_L g3717 ( 
.A(n_3677),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3658),
.B(n_4),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3685),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_L g3720 ( 
.A(n_3704),
.B(n_5),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3695),
.B(n_1577),
.Y(n_3721)
);

INVxp67_ASAP7_75t_SL g3722 ( 
.A(n_3693),
.Y(n_3722)
);

INVx2_ASAP7_75t_SL g3723 ( 
.A(n_3690),
.Y(n_3723)
);

AND2x4_ASAP7_75t_L g3724 ( 
.A(n_3691),
.B(n_6),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3698),
.Y(n_3725)
);

AOI222xp33_ASAP7_75t_L g3726 ( 
.A1(n_3697),
.A2(n_1583),
.B1(n_1580),
.B2(n_1587),
.C1(n_1585),
.C2(n_1582),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3717),
.B(n_6),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3689),
.B(n_7),
.Y(n_3728)
);

AND2x4_ASAP7_75t_SL g3729 ( 
.A(n_3719),
.B(n_1345),
.Y(n_3729)
);

INVx3_ASAP7_75t_L g3730 ( 
.A(n_3702),
.Y(n_3730)
);

OR2x2_ASAP7_75t_L g3731 ( 
.A(n_3687),
.B(n_7),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3707),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3696),
.B(n_3700),
.Y(n_3733)
);

AND2x2_ASAP7_75t_L g3734 ( 
.A(n_3713),
.B(n_8),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3694),
.A2(n_1673),
.B1(n_1345),
.B2(n_1593),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3708),
.Y(n_3736)
);

AO21x2_ASAP7_75t_L g3737 ( 
.A1(n_3715),
.A2(n_1673),
.B(n_8),
.Y(n_3737)
);

O2A1O1Ixp5_ASAP7_75t_L g3738 ( 
.A1(n_3709),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3708),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3688),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3710),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3712),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_3705),
.B(n_11),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3716),
.B(n_13),
.Y(n_3744)
);

AO21x2_ASAP7_75t_L g3745 ( 
.A1(n_3714),
.A2(n_1673),
.B(n_13),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3703),
.B(n_1588),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3692),
.B(n_16),
.Y(n_3747)
);

BUFx2_ASAP7_75t_L g3748 ( 
.A(n_3711),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3699),
.B(n_17),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3718),
.B(n_17),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3712),
.B(n_1599),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3706),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3711),
.Y(n_3753)
);

AOI221xp5_ASAP7_75t_L g3754 ( 
.A1(n_3701),
.A2(n_1603),
.B1(n_1605),
.B2(n_1604),
.C(n_1600),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3730),
.B(n_18),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3733),
.Y(n_3756)
);

AND2x2_ASAP7_75t_SL g3757 ( 
.A(n_3748),
.B(n_1345),
.Y(n_3757)
);

AND2x4_ASAP7_75t_L g3758 ( 
.A(n_3730),
.B(n_18),
.Y(n_3758)
);

AND2x2_ASAP7_75t_L g3759 ( 
.A(n_3723),
.B(n_20),
.Y(n_3759)
);

BUFx2_ASAP7_75t_L g3760 ( 
.A(n_3722),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3736),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3728),
.B(n_21),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3725),
.Y(n_3763)
);

OR2x2_ASAP7_75t_L g3764 ( 
.A(n_3741),
.B(n_22),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3727),
.B(n_3724),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3724),
.B(n_22),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3743),
.B(n_23),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3741),
.B(n_23),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3747),
.B(n_24),
.Y(n_3769)
);

INVxp67_ASAP7_75t_L g3770 ( 
.A(n_3720),
.Y(n_3770)
);

AND2x4_ASAP7_75t_L g3771 ( 
.A(n_3734),
.B(n_3753),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3731),
.Y(n_3772)
);

AND2x4_ASAP7_75t_L g3773 ( 
.A(n_3737),
.B(n_24),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3740),
.Y(n_3774)
);

OR2x2_ASAP7_75t_L g3775 ( 
.A(n_3721),
.B(n_25),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3740),
.Y(n_3776)
);

AND2x4_ASAP7_75t_L g3777 ( 
.A(n_3750),
.B(n_29),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3744),
.B(n_29),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3752),
.Y(n_3779)
);

NOR3xp33_ASAP7_75t_L g3780 ( 
.A(n_3738),
.B(n_1621),
.C(n_1614),
.Y(n_3780)
);

OR2x2_ASAP7_75t_L g3781 ( 
.A(n_3749),
.B(n_30),
.Y(n_3781)
);

HB1xp67_ASAP7_75t_L g3782 ( 
.A(n_3751),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3729),
.B(n_30),
.Y(n_3783)
);

AND2x2_ASAP7_75t_L g3784 ( 
.A(n_3742),
.B(n_31),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3745),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3732),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3726),
.B(n_32),
.Y(n_3787)
);

AND2x4_ASAP7_75t_SL g3788 ( 
.A(n_3765),
.B(n_3739),
.Y(n_3788)
);

INVxp67_ASAP7_75t_L g3789 ( 
.A(n_3760),
.Y(n_3789)
);

OR2x2_ASAP7_75t_L g3790 ( 
.A(n_3760),
.B(n_3746),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3774),
.Y(n_3791)
);

INVx1_ASAP7_75t_SL g3792 ( 
.A(n_3767),
.Y(n_3792)
);

INVx1_ASAP7_75t_SL g3793 ( 
.A(n_3777),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3759),
.B(n_3735),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3772),
.B(n_3754),
.Y(n_3795)
);

NOR2xp33_ASAP7_75t_L g3796 ( 
.A(n_3770),
.B(n_3764),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_3755),
.B(n_32),
.Y(n_3797)
);

OR2x2_ASAP7_75t_L g3798 ( 
.A(n_3756),
.B(n_33),
.Y(n_3798)
);

OR2x2_ASAP7_75t_L g3799 ( 
.A(n_3763),
.B(n_35),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3776),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3779),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3784),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3768),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3773),
.B(n_1624),
.Y(n_3804)
);

NOR2xp33_ASAP7_75t_L g3805 ( 
.A(n_3758),
.B(n_3775),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3762),
.B(n_35),
.Y(n_3806)
);

OR2x2_ASAP7_75t_L g3807 ( 
.A(n_3786),
.B(n_36),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3782),
.Y(n_3808)
);

AOI22xp5_ASAP7_75t_L g3809 ( 
.A1(n_3773),
.A2(n_3785),
.B1(n_3771),
.B2(n_3780),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3781),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3766),
.B(n_39),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3769),
.B(n_1625),
.Y(n_3812)
);

INVx1_ASAP7_75t_SL g3813 ( 
.A(n_3778),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3761),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3771),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3783),
.B(n_40),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3787),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3757),
.B(n_1628),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3760),
.B(n_1629),
.Y(n_3819)
);

OR2x2_ASAP7_75t_L g3820 ( 
.A(n_3760),
.B(n_40),
.Y(n_3820)
);

NOR2xp33_ASAP7_75t_L g3821 ( 
.A(n_3770),
.B(n_1632),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3765),
.B(n_41),
.Y(n_3822)
);

OR2x2_ASAP7_75t_L g3823 ( 
.A(n_3760),
.B(n_41),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3765),
.Y(n_3824)
);

OR2x2_ASAP7_75t_L g3825 ( 
.A(n_3760),
.B(n_42),
.Y(n_3825)
);

NAND3xp33_ASAP7_75t_SL g3826 ( 
.A(n_3760),
.B(n_1635),
.C(n_1634),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3765),
.Y(n_3827)
);

OR2x2_ASAP7_75t_L g3828 ( 
.A(n_3760),
.B(n_43),
.Y(n_3828)
);

INVx2_ASAP7_75t_SL g3829 ( 
.A(n_3765),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3774),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3774),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3760),
.B(n_1636),
.Y(n_3832)
);

INVx1_ASAP7_75t_SL g3833 ( 
.A(n_3792),
.Y(n_3833)
);

CKINVDCx16_ASAP7_75t_R g3834 ( 
.A(n_3806),
.Y(n_3834)
);

HB1xp67_ASAP7_75t_L g3835 ( 
.A(n_3813),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3810),
.Y(n_3836)
);

HB1xp67_ASAP7_75t_L g3837 ( 
.A(n_3789),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3810),
.Y(n_3838)
);

AOI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3817),
.A2(n_1673),
.B1(n_1345),
.B2(n_1643),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3803),
.B(n_1640),
.Y(n_3840)
);

BUFx3_ASAP7_75t_L g3841 ( 
.A(n_3822),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3802),
.B(n_1645),
.Y(n_3842)
);

INVx2_ASAP7_75t_SL g3843 ( 
.A(n_3788),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3820),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3796),
.B(n_1646),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3829),
.B(n_43),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3823),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3824),
.B(n_45),
.Y(n_3848)
);

HB1xp67_ASAP7_75t_L g3849 ( 
.A(n_3827),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3825),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3793),
.B(n_45),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3828),
.Y(n_3852)
);

INVx2_ASAP7_75t_SL g3853 ( 
.A(n_3811),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3805),
.B(n_46),
.Y(n_3854)
);

INVxp67_ASAP7_75t_SL g3855 ( 
.A(n_3819),
.Y(n_3855)
);

NAND2x1p5_ASAP7_75t_L g3856 ( 
.A(n_3797),
.B(n_47),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3790),
.B(n_48),
.Y(n_3857)
);

OR2x2_ASAP7_75t_L g3858 ( 
.A(n_3808),
.B(n_3832),
.Y(n_3858)
);

OR2x2_ASAP7_75t_L g3859 ( 
.A(n_3799),
.B(n_49),
.Y(n_3859)
);

AND2x4_ASAP7_75t_L g3860 ( 
.A(n_3816),
.B(n_50),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3801),
.B(n_50),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3791),
.Y(n_3862)
);

NOR2x1_ASAP7_75t_L g3863 ( 
.A(n_3826),
.B(n_53),
.Y(n_3863)
);

INVxp67_ASAP7_75t_L g3864 ( 
.A(n_3821),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3800),
.Y(n_3865)
);

INVxp67_ASAP7_75t_SL g3866 ( 
.A(n_3804),
.Y(n_3866)
);

NOR4xp25_ASAP7_75t_L g3867 ( 
.A(n_3795),
.B(n_3815),
.C(n_3831),
.D(n_3830),
.Y(n_3867)
);

NAND4xp75_ASAP7_75t_L g3868 ( 
.A(n_3809),
.B(n_3814),
.C(n_3794),
.D(n_3818),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3798),
.B(n_52),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3812),
.B(n_53),
.Y(n_3870)
);

AND3x1_ASAP7_75t_L g3871 ( 
.A(n_3807),
.B(n_54),
.C(n_55),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3810),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3829),
.B(n_55),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3810),
.Y(n_3874)
);

AND3x2_ASAP7_75t_L g3875 ( 
.A(n_3789),
.B(n_56),
.C(n_57),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3829),
.B(n_56),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3810),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3810),
.Y(n_3878)
);

INVx1_ASAP7_75t_SL g3879 ( 
.A(n_3792),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3829),
.B(n_57),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3829),
.B(n_59),
.Y(n_3881)
);

OR2x2_ASAP7_75t_L g3882 ( 
.A(n_3792),
.B(n_60),
.Y(n_3882)
);

HB1xp67_ASAP7_75t_L g3883 ( 
.A(n_3792),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3829),
.B(n_60),
.Y(n_3884)
);

AND2x4_ASAP7_75t_L g3885 ( 
.A(n_3829),
.B(n_62),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3810),
.Y(n_3886)
);

OR2x2_ASAP7_75t_L g3887 ( 
.A(n_3792),
.B(n_62),
.Y(n_3887)
);

AND2x4_ASAP7_75t_L g3888 ( 
.A(n_3829),
.B(n_63),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3813),
.B(n_1653),
.Y(n_3889)
);

INVx2_ASAP7_75t_SL g3890 ( 
.A(n_3788),
.Y(n_3890)
);

NOR2xp33_ASAP7_75t_L g3891 ( 
.A(n_3826),
.B(n_1656),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3813),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3813),
.Y(n_3893)
);

OR2x6_ASAP7_75t_L g3894 ( 
.A(n_3816),
.B(n_63),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3829),
.B(n_64),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3810),
.Y(n_3896)
);

AND2x2_ASAP7_75t_L g3897 ( 
.A(n_3829),
.B(n_64),
.Y(n_3897)
);

INVx1_ASAP7_75t_SL g3898 ( 
.A(n_3834),
.Y(n_3898)
);

INVx1_ASAP7_75t_SL g3899 ( 
.A(n_3841),
.Y(n_3899)
);

OR2x2_ASAP7_75t_L g3900 ( 
.A(n_3867),
.B(n_3833),
.Y(n_3900)
);

OR2x2_ASAP7_75t_L g3901 ( 
.A(n_3879),
.B(n_65),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3853),
.B(n_1657),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3835),
.B(n_1658),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3883),
.B(n_1659),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3875),
.B(n_3857),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3856),
.B(n_1660),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3843),
.B(n_1662),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3837),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3849),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3882),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3887),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3859),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3855),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3844),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3890),
.B(n_1663),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3894),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_3876),
.B(n_1668),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3848),
.B(n_1669),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3861),
.B(n_1672),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3894),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3847),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3846),
.B(n_1677),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3850),
.B(n_1684),
.Y(n_3923)
);

OR2x2_ASAP7_75t_L g3924 ( 
.A(n_3892),
.B(n_65),
.Y(n_3924)
);

OR2x4_ASAP7_75t_L g3925 ( 
.A(n_3858),
.B(n_67),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3873),
.B(n_1686),
.Y(n_3926)
);

OR2x2_ASAP7_75t_L g3927 ( 
.A(n_3893),
.B(n_3852),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3885),
.B(n_1691),
.Y(n_3928)
);

INVxp67_ASAP7_75t_SL g3929 ( 
.A(n_3863),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3888),
.B(n_1695),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3869),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3880),
.B(n_3881),
.Y(n_3932)
);

NAND3xp33_ASAP7_75t_L g3933 ( 
.A(n_3839),
.B(n_1698),
.C(n_1697),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3851),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3884),
.B(n_3897),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3895),
.B(n_1700),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3866),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3854),
.B(n_1706),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3842),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3864),
.B(n_1708),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3836),
.B(n_3838),
.Y(n_3941)
);

OR2x2_ASAP7_75t_L g3942 ( 
.A(n_3889),
.B(n_67),
.Y(n_3942)
);

INVx1_ASAP7_75t_SL g3943 ( 
.A(n_3860),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3871),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3870),
.B(n_1710),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3872),
.B(n_1716),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3840),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_L g3948 ( 
.A1(n_3845),
.A2(n_1673),
.B1(n_1727),
.B2(n_1724),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3874),
.B(n_1730),
.Y(n_3949)
);

INVxp67_ASAP7_75t_L g3950 ( 
.A(n_3891),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3877),
.B(n_1732),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3878),
.B(n_1735),
.Y(n_3952)
);

INVxp67_ASAP7_75t_L g3953 ( 
.A(n_3868),
.Y(n_3953)
);

NAND3xp33_ASAP7_75t_L g3954 ( 
.A(n_3886),
.B(n_1738),
.C(n_1736),
.Y(n_3954)
);

HB1xp67_ASAP7_75t_L g3955 ( 
.A(n_3896),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3862),
.B(n_1739),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3865),
.B(n_1741),
.Y(n_3957)
);

INVxp67_ASAP7_75t_L g3958 ( 
.A(n_3868),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3835),
.Y(n_3959)
);

INVx1_ASAP7_75t_SL g3960 ( 
.A(n_3834),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3835),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3835),
.Y(n_3962)
);

NOR3xp33_ASAP7_75t_SL g3963 ( 
.A(n_3834),
.B(n_1748),
.C(n_1744),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3867),
.A2(n_1755),
.B(n_1749),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3835),
.Y(n_3965)
);

BUFx2_ASAP7_75t_L g3966 ( 
.A(n_3841),
.Y(n_3966)
);

NOR2xp33_ASAP7_75t_L g3967 ( 
.A(n_3834),
.B(n_1760),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_L g3968 ( 
.A(n_3834),
.B(n_1762),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3835),
.Y(n_3969)
);

INVx2_ASAP7_75t_SL g3970 ( 
.A(n_3841),
.Y(n_3970)
);

HB1xp67_ASAP7_75t_L g3971 ( 
.A(n_3834),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3835),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3835),
.B(n_1763),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3856),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3834),
.B(n_1769),
.Y(n_3975)
);

INVx1_ASAP7_75t_SL g3976 ( 
.A(n_3834),
.Y(n_3976)
);

INVx2_ASAP7_75t_SL g3977 ( 
.A(n_3841),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3834),
.B(n_68),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3835),
.B(n_68),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3835),
.B(n_69),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3835),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3856),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3834),
.B(n_69),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3835),
.B(n_70),
.Y(n_3984)
);

AOI22xp5_ASAP7_75t_L g3985 ( 
.A1(n_3953),
.A2(n_1308),
.B1(n_1310),
.B2(n_1301),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3898),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3900),
.A2(n_1767),
.B1(n_1320),
.B2(n_1324),
.Y(n_3987)
);

AOI221xp5_ASAP7_75t_L g3988 ( 
.A1(n_3958),
.A2(n_1332),
.B1(n_1334),
.B2(n_1326),
.C(n_1314),
.Y(n_3988)
);

OAI22xp5_ASAP7_75t_L g3989 ( 
.A1(n_3960),
.A2(n_3976),
.B1(n_3971),
.B2(n_3899),
.Y(n_3989)
);

OAI22xp33_ASAP7_75t_L g3990 ( 
.A1(n_3929),
.A2(n_1337),
.B1(n_1348),
.B2(n_1335),
.Y(n_3990)
);

NOR3xp33_ASAP7_75t_L g3991 ( 
.A(n_3913),
.B(n_1355),
.C(n_1351),
.Y(n_3991)
);

INVxp67_ASAP7_75t_L g3992 ( 
.A(n_3966),
.Y(n_3992)
);

AOI31xp33_ASAP7_75t_L g3993 ( 
.A1(n_3959),
.A2(n_3977),
.A3(n_3970),
.B(n_3962),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3979),
.Y(n_3994)
);

OAI211xp5_ASAP7_75t_L g3995 ( 
.A1(n_3959),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_3995)
);

NOR3xp33_ASAP7_75t_SL g3996 ( 
.A(n_3961),
.B(n_71),
.C(n_72),
.Y(n_3996)
);

AOI21xp33_ASAP7_75t_L g3997 ( 
.A1(n_3944),
.A2(n_73),
.B(n_75),
.Y(n_3997)
);

OAI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3964),
.A2(n_73),
.B(n_76),
.Y(n_3998)
);

OAI221xp5_ASAP7_75t_L g3999 ( 
.A1(n_3905),
.A2(n_1386),
.B1(n_1388),
.B2(n_1361),
.C(n_1358),
.Y(n_3999)
);

AOI31xp33_ASAP7_75t_L g4000 ( 
.A1(n_3965),
.A2(n_3972),
.A3(n_3981),
.B(n_3969),
.Y(n_4000)
);

OAI211xp5_ASAP7_75t_L g4001 ( 
.A1(n_3908),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_4001)
);

OAI221xp5_ASAP7_75t_L g4002 ( 
.A1(n_3910),
.A2(n_1394),
.B1(n_1396),
.B2(n_1391),
.C(n_1390),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3967),
.B(n_3968),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_SL g4004 ( 
.A(n_3943),
.B(n_1407),
.Y(n_4004)
);

INVxp67_ASAP7_75t_SL g4005 ( 
.A(n_3975),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3980),
.B(n_77),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3922),
.B(n_78),
.Y(n_4007)
);

INVx1_ASAP7_75t_SL g4008 ( 
.A(n_3932),
.Y(n_4008)
);

AOI22xp5_ASAP7_75t_L g4009 ( 
.A1(n_3911),
.A2(n_1416),
.B1(n_1435),
.B2(n_1408),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3984),
.Y(n_4010)
);

AOI31xp33_ASAP7_75t_L g4011 ( 
.A1(n_3927),
.A2(n_82),
.A3(n_79),
.B(n_81),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3935),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3926),
.B(n_79),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3978),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3983),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3925),
.A2(n_3955),
.B(n_3938),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3901),
.Y(n_4017)
);

AOI221xp5_ASAP7_75t_L g4018 ( 
.A1(n_3937),
.A2(n_1452),
.B1(n_1454),
.B2(n_1444),
.C(n_1443),
.Y(n_4018)
);

NAND4xp25_ASAP7_75t_L g4019 ( 
.A(n_3909),
.B(n_86),
.C(n_84),
.D(n_85),
.Y(n_4019)
);

INVx1_ASAP7_75t_SL g4020 ( 
.A(n_3936),
.Y(n_4020)
);

OAI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3931),
.A2(n_84),
.B(n_87),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3940),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3934),
.B(n_87),
.Y(n_4023)
);

OAI21xp5_ASAP7_75t_SL g4024 ( 
.A1(n_3914),
.A2(n_88),
.B(n_89),
.Y(n_4024)
);

NAND2x1_ASAP7_75t_L g4025 ( 
.A(n_3963),
.B(n_88),
.Y(n_4025)
);

OAI22xp33_ASAP7_75t_L g4026 ( 
.A1(n_3924),
.A2(n_1470),
.B1(n_1482),
.B2(n_1459),
.Y(n_4026)
);

OR2x2_ASAP7_75t_L g4027 ( 
.A(n_3921),
.B(n_89),
.Y(n_4027)
);

XOR2x2_ASAP7_75t_L g4028 ( 
.A(n_3945),
.B(n_91),
.Y(n_4028)
);

AOI22xp5_ASAP7_75t_L g4029 ( 
.A1(n_3939),
.A2(n_3947),
.B1(n_3912),
.B2(n_3974),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3902),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_L g4031 ( 
.A(n_3982),
.B(n_90),
.Y(n_4031)
);

AOI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_3923),
.A2(n_92),
.B(n_94),
.Y(n_4032)
);

OAI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3954),
.A2(n_1489),
.B1(n_1493),
.B2(n_1483),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3941),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3903),
.Y(n_4035)
);

AOI211xp5_ASAP7_75t_L g4036 ( 
.A1(n_3904),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_4036)
);

NOR2xp33_ASAP7_75t_L g4037 ( 
.A(n_3973),
.B(n_99),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3916),
.Y(n_4038)
);

OAI22xp33_ASAP7_75t_L g4039 ( 
.A1(n_3920),
.A2(n_1513),
.B1(n_1526),
.B2(n_1506),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3907),
.B(n_99),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3956),
.Y(n_4041)
);

AOI22xp5_ASAP7_75t_L g4042 ( 
.A1(n_3950),
.A2(n_3918),
.B1(n_3919),
.B2(n_3906),
.Y(n_4042)
);

AOI22xp5_ASAP7_75t_L g4043 ( 
.A1(n_3946),
.A2(n_1540),
.B1(n_1545),
.B2(n_1538),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3942),
.Y(n_4044)
);

INVxp67_ASAP7_75t_L g4045 ( 
.A(n_3917),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3949),
.Y(n_4046)
);

NOR2xp33_ASAP7_75t_L g4047 ( 
.A(n_3915),
.B(n_100),
.Y(n_4047)
);

OAI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3951),
.A2(n_1552),
.B1(n_1553),
.B2(n_1546),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3957),
.B(n_3952),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_3928),
.B(n_100),
.Y(n_4050)
);

OAI22xp33_ASAP7_75t_L g4051 ( 
.A1(n_3933),
.A2(n_1560),
.B1(n_1561),
.B2(n_1558),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3948),
.A2(n_1655),
.B1(n_1702),
.B2(n_1598),
.Y(n_4052)
);

INVxp67_ASAP7_75t_L g4053 ( 
.A(n_3930),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3898),
.B(n_101),
.Y(n_4054)
);

INVx2_ASAP7_75t_SL g4055 ( 
.A(n_3971),
.Y(n_4055)
);

AOI211x1_ASAP7_75t_L g4056 ( 
.A1(n_3959),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3971),
.Y(n_4057)
);

NOR3xp33_ASAP7_75t_SL g4058 ( 
.A(n_3961),
.B(n_103),
.C(n_104),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3971),
.Y(n_4059)
);

O2A1O1Ixp33_ASAP7_75t_SL g4060 ( 
.A1(n_3900),
.A2(n_108),
.B(n_105),
.C(n_107),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3898),
.B(n_110),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3971),
.Y(n_4062)
);

OAI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_3900),
.A2(n_110),
.B(n_111),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3971),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3898),
.B(n_111),
.Y(n_4065)
);

OR2x2_ASAP7_75t_L g4066 ( 
.A(n_3898),
.B(n_112),
.Y(n_4066)
);

INVxp33_ASAP7_75t_L g4067 ( 
.A(n_3971),
.Y(n_4067)
);

AOI22xp5_ASAP7_75t_L g4068 ( 
.A1(n_3953),
.A2(n_1579),
.B1(n_1581),
.B2(n_1570),
.Y(n_4068)
);

OAI22xp33_ASAP7_75t_L g4069 ( 
.A1(n_3900),
.A2(n_1592),
.B1(n_1596),
.B2(n_1589),
.Y(n_4069)
);

INVx1_ASAP7_75t_SL g4070 ( 
.A(n_3898),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3898),
.Y(n_4071)
);

OAI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_3900),
.A2(n_1611),
.B1(n_1616),
.B2(n_1597),
.Y(n_4072)
);

AOI322xp5_ASAP7_75t_L g4073 ( 
.A1(n_3929),
.A2(n_118),
.A3(n_117),
.B1(n_115),
.B2(n_112),
.C1(n_114),
.C2(n_116),
.Y(n_4073)
);

AND2x4_ASAP7_75t_L g4074 ( 
.A(n_3898),
.B(n_118),
.Y(n_4074)
);

AOI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_3953),
.A2(n_1639),
.B1(n_1641),
.B2(n_1633),
.Y(n_4075)
);

AOI222xp33_ASAP7_75t_L g4076 ( 
.A1(n_3953),
.A2(n_1664),
.B1(n_1649),
.B2(n_1666),
.C1(n_1661),
.C2(n_1648),
.Y(n_4076)
);

AOI21xp33_ASAP7_75t_SL g4077 ( 
.A1(n_3900),
.A2(n_119),
.B(n_120),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3971),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3953),
.A2(n_1718),
.B1(n_1680),
.B2(n_1687),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3900),
.A2(n_1764),
.B1(n_1766),
.B2(n_1758),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3898),
.B(n_120),
.Y(n_4081)
);

NOR2x1_ASAP7_75t_L g4082 ( 
.A(n_3900),
.B(n_121),
.Y(n_4082)
);

OAI21xp33_ASAP7_75t_SL g4083 ( 
.A1(n_3900),
.A2(n_121),
.B(n_122),
.Y(n_4083)
);

O2A1O1Ixp33_ASAP7_75t_L g4084 ( 
.A1(n_3900),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_4084)
);

NOR3xp33_ASAP7_75t_L g4085 ( 
.A(n_3953),
.B(n_1694),
.C(n_1679),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3898),
.Y(n_4086)
);

OAI211xp5_ASAP7_75t_SL g4087 ( 
.A1(n_3900),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_4087)
);

AND2x2_ASAP7_75t_L g4088 ( 
.A(n_3898),
.B(n_127),
.Y(n_4088)
);

OR2x2_ASAP7_75t_L g4089 ( 
.A(n_3898),
.B(n_130),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3898),
.B(n_131),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3971),
.Y(n_4091)
);

AOI22xp5_ASAP7_75t_L g4092 ( 
.A1(n_3953),
.A2(n_1709),
.B1(n_1731),
.B2(n_1723),
.Y(n_4092)
);

OAI21xp5_ASAP7_75t_L g4093 ( 
.A1(n_3900),
.A2(n_131),
.B(n_132),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3971),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3971),
.Y(n_4095)
);

AOI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_3964),
.A2(n_132),
.B(n_133),
.Y(n_4096)
);

NAND3xp33_ASAP7_75t_L g4097 ( 
.A(n_3900),
.B(n_1704),
.C(n_134),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3898),
.Y(n_4098)
);

NOR2xp33_ASAP7_75t_L g4099 ( 
.A(n_3898),
.B(n_134),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3971),
.Y(n_4100)
);

OAI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_3900),
.A2(n_135),
.B(n_136),
.Y(n_4101)
);

O2A1O1Ixp33_ASAP7_75t_L g4102 ( 
.A1(n_3900),
.A2(n_139),
.B(n_137),
.C(n_138),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3971),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3898),
.B(n_140),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3898),
.B(n_140),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3971),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3971),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3898),
.B(n_141),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3898),
.B(n_142),
.Y(n_4109)
);

OAI221xp5_ASAP7_75t_L g4110 ( 
.A1(n_3929),
.A2(n_147),
.B1(n_143),
.B2(n_145),
.C(n_149),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3971),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3971),
.Y(n_4112)
);

OAI21xp5_ASAP7_75t_SL g4113 ( 
.A1(n_3900),
.A2(n_150),
.B(n_151),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3971),
.Y(n_4114)
);

NOR2xp33_ASAP7_75t_L g4115 ( 
.A(n_3898),
.B(n_152),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3971),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3971),
.Y(n_4117)
);

OR3x1_ASAP7_75t_L g4118 ( 
.A(n_3959),
.B(n_152),
.C(n_153),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3971),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3898),
.B(n_153),
.Y(n_4120)
);

OAI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_3900),
.A2(n_158),
.B1(n_154),
.B2(n_155),
.Y(n_4121)
);

NOR3xp33_ASAP7_75t_SL g4122 ( 
.A(n_3961),
.B(n_154),
.C(n_155),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3971),
.Y(n_4123)
);

INVxp67_ASAP7_75t_SL g4124 ( 
.A(n_3971),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3971),
.Y(n_4125)
);

OAI322xp33_ASAP7_75t_L g4126 ( 
.A1(n_3900),
.A2(n_165),
.A3(n_163),
.B1(n_161),
.B2(n_158),
.C1(n_160),
.C2(n_162),
.Y(n_4126)
);

AOI311xp33_ASAP7_75t_L g4127 ( 
.A1(n_3961),
.A2(n_166),
.A3(n_160),
.B(n_161),
.C(n_168),
.Y(n_4127)
);

OR2x2_ASAP7_75t_L g4128 ( 
.A(n_3898),
.B(n_166),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_3898),
.Y(n_4129)
);

OAI21xp33_ASAP7_75t_L g4130 ( 
.A1(n_3898),
.A2(n_169),
.B(n_170),
.Y(n_4130)
);

NAND4xp25_ASAP7_75t_L g4131 ( 
.A(n_3898),
.B(n_171),
.C(n_169),
.D(n_170),
.Y(n_4131)
);

AOI211xp5_ASAP7_75t_L g4132 ( 
.A1(n_3900),
.A2(n_175),
.B(n_172),
.C(n_174),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3971),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_3898),
.Y(n_4134)
);

AND2x4_ASAP7_75t_L g4135 ( 
.A(n_4012),
.B(n_4070),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_4124),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_4074),
.B(n_172),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_4028),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4008),
.B(n_174),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3986),
.Y(n_4140)
);

OR2x2_ASAP7_75t_L g4141 ( 
.A(n_4071),
.B(n_175),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4086),
.Y(n_4142)
);

INVx1_ASAP7_75t_SL g4143 ( 
.A(n_4118),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4098),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4129),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_4074),
.B(n_178),
.Y(n_4146)
);

NOR2x1_ASAP7_75t_L g4147 ( 
.A(n_4097),
.B(n_179),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_4088),
.B(n_179),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_4056),
.B(n_180),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4134),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4109),
.B(n_180),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4055),
.B(n_181),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4006),
.Y(n_4153)
);

OR2x2_ASAP7_75t_L g4154 ( 
.A(n_4066),
.B(n_4089),
.Y(n_4154)
);

INVx1_ASAP7_75t_SL g4155 ( 
.A(n_4128),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_4040),
.Y(n_4156)
);

INVx2_ASAP7_75t_SL g4157 ( 
.A(n_4057),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_4067),
.B(n_182),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_3992),
.B(n_185),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4011),
.B(n_186),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_4020),
.B(n_188),
.Y(n_4161)
);

INVx2_ASAP7_75t_SL g4162 ( 
.A(n_4059),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3996),
.B(n_189),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4058),
.B(n_190),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4062),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4064),
.Y(n_4166)
);

INVxp33_ASAP7_75t_L g4167 ( 
.A(n_4082),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4078),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_4122),
.B(n_191),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_SL g4170 ( 
.A(n_3989),
.B(n_2198),
.Y(n_4170)
);

INVx1_ASAP7_75t_SL g4171 ( 
.A(n_4054),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4037),
.B(n_191),
.Y(n_4172)
);

HB1xp67_ASAP7_75t_L g4173 ( 
.A(n_4091),
.Y(n_4173)
);

INVx1_ASAP7_75t_SL g4174 ( 
.A(n_4061),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4094),
.Y(n_4175)
);

OR2x2_ASAP7_75t_L g4176 ( 
.A(n_4034),
.B(n_192),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4095),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4100),
.Y(n_4178)
);

INVx1_ASAP7_75t_SL g4179 ( 
.A(n_4065),
.Y(n_4179)
);

OR2x2_ASAP7_75t_L g4180 ( 
.A(n_4081),
.B(n_194),
.Y(n_4180)
);

INVxp67_ASAP7_75t_L g4181 ( 
.A(n_4099),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4103),
.Y(n_4182)
);

OAI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_4000),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_4183)
);

OR2x2_ASAP7_75t_L g4184 ( 
.A(n_4090),
.B(n_195),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3994),
.B(n_198),
.Y(n_4185)
);

INVx1_ASAP7_75t_SL g4186 ( 
.A(n_4104),
.Y(n_4186)
);

OR2x2_ASAP7_75t_L g4187 ( 
.A(n_4105),
.B(n_198),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4106),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_L g4189 ( 
.A(n_4083),
.B(n_199),
.Y(n_4189)
);

AOI22xp33_ASAP7_75t_L g4190 ( 
.A1(n_4087),
.A2(n_3987),
.B1(n_4080),
.B2(n_4072),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_4107),
.B(n_4111),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4112),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_4114),
.B(n_200),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4116),
.Y(n_4194)
);

OR2x2_ASAP7_75t_L g4195 ( 
.A(n_4108),
.B(n_202),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4117),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4119),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4123),
.Y(n_4198)
);

INVx1_ASAP7_75t_SL g4199 ( 
.A(n_4120),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4010),
.B(n_202),
.Y(n_4200)
);

OR2x2_ASAP7_75t_L g4201 ( 
.A(n_4125),
.B(n_204),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_4133),
.B(n_204),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_4047),
.B(n_4005),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4027),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4044),
.Y(n_4205)
);

NAND2x1p5_ASAP7_75t_L g4206 ( 
.A(n_4025),
.B(n_206),
.Y(n_4206)
);

NOR2xp33_ASAP7_75t_L g4207 ( 
.A(n_4131),
.B(n_205),
.Y(n_4207)
);

NOR2x1_ASAP7_75t_L g4208 ( 
.A(n_4113),
.B(n_206),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4077),
.B(n_207),
.Y(n_4209)
);

INVxp33_ASAP7_75t_L g4210 ( 
.A(n_4115),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4017),
.Y(n_4211)
);

NOR2x1_ASAP7_75t_L g4212 ( 
.A(n_3993),
.B(n_207),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4007),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4013),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4049),
.B(n_4035),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4036),
.B(n_208),
.Y(n_4216)
);

AND2x2_ASAP7_75t_SL g4217 ( 
.A(n_4003),
.B(n_210),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_4063),
.B(n_211),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_4093),
.B(n_212),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4023),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_4024),
.B(n_213),
.Y(n_4221)
);

OR2x2_ASAP7_75t_L g4222 ( 
.A(n_4121),
.B(n_213),
.Y(n_4222)
);

OAI21xp33_ASAP7_75t_L g4223 ( 
.A1(n_4022),
.A2(n_214),
.B(n_215),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_4101),
.B(n_4127),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4041),
.Y(n_4225)
);

OAI31xp33_ASAP7_75t_L g4226 ( 
.A1(n_4069),
.A2(n_4060),
.A3(n_4102),
.B(n_4084),
.Y(n_4226)
);

HB1xp67_ASAP7_75t_L g4227 ( 
.A(n_4046),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_4050),
.Y(n_4228)
);

INVx1_ASAP7_75t_SL g4229 ( 
.A(n_4004),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_4132),
.B(n_214),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4014),
.Y(n_4231)
);

OA21x2_ASAP7_75t_L g4232 ( 
.A1(n_4016),
.A2(n_215),
.B(n_217),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4031),
.B(n_217),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4015),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4032),
.B(n_218),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_4076),
.B(n_219),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_4096),
.B(n_223),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_3995),
.B(n_223),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4038),
.Y(n_4239)
);

NOR2xp33_ASAP7_75t_L g4240 ( 
.A(n_4126),
.B(n_224),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4001),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4042),
.B(n_224),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4029),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4030),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4019),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4110),
.Y(n_4246)
);

OR2x2_ASAP7_75t_L g4247 ( 
.A(n_4021),
.B(n_225),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4045),
.Y(n_4248)
);

OR2x2_ASAP7_75t_L g4249 ( 
.A(n_4053),
.B(n_225),
.Y(n_4249)
);

AND2x4_ASAP7_75t_L g4250 ( 
.A(n_3998),
.B(n_226),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4130),
.B(n_227),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4009),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_3991),
.B(n_228),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4143),
.B(n_4026),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4135),
.B(n_4079),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_4212),
.B(n_3985),
.Y(n_4256)
);

INVxp67_ASAP7_75t_L g4257 ( 
.A(n_4189),
.Y(n_4257)
);

AOI22xp5_ASAP7_75t_L g4258 ( 
.A1(n_4155),
.A2(n_4085),
.B1(n_4068),
.B2(n_4075),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4215),
.Y(n_4259)
);

AOI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_4171),
.A2(n_3999),
.B1(n_3997),
.B2(n_4092),
.Y(n_4260)
);

INVx2_ASAP7_75t_SL g4261 ( 
.A(n_4139),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_4217),
.B(n_4073),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4154),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4206),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4137),
.Y(n_4265)
);

AND2x2_ASAP7_75t_L g4266 ( 
.A(n_4227),
.B(n_4043),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4146),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4148),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4151),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4191),
.B(n_3988),
.Y(n_4270)
);

OR2x2_ASAP7_75t_L g4271 ( 
.A(n_4136),
.B(n_4002),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4173),
.Y(n_4272)
);

NOR2xp67_ASAP7_75t_L g4273 ( 
.A(n_4140),
.B(n_4033),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4153),
.B(n_4048),
.Y(n_4274)
);

INVxp67_ASAP7_75t_L g4275 ( 
.A(n_4208),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4203),
.Y(n_4276)
);

INVx1_ASAP7_75t_SL g4277 ( 
.A(n_4152),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4228),
.B(n_3990),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4224),
.B(n_4051),
.Y(n_4279)
);

INVxp67_ASAP7_75t_L g4280 ( 
.A(n_4232),
.Y(n_4280)
);

OA21x2_ASAP7_75t_L g4281 ( 
.A1(n_4243),
.A2(n_4052),
.B(n_4018),
.Y(n_4281)
);

NAND2x1_ASAP7_75t_L g4282 ( 
.A(n_4142),
.B(n_4039),
.Y(n_4282)
);

OR2x2_ASAP7_75t_L g4283 ( 
.A(n_4144),
.B(n_230),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4156),
.Y(n_4284)
);

NOR3xp33_ASAP7_75t_SL g4285 ( 
.A(n_4145),
.B(n_232),
.C(n_234),
.Y(n_4285)
);

NOR2xp33_ASAP7_75t_L g4286 ( 
.A(n_4210),
.B(n_232),
.Y(n_4286)
);

NOR2xp33_ASAP7_75t_L g4287 ( 
.A(n_4167),
.B(n_235),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4149),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_4193),
.B(n_236),
.Y(n_4289)
);

BUFx2_ASAP7_75t_L g4290 ( 
.A(n_4150),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4158),
.B(n_236),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_4202),
.B(n_237),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4250),
.B(n_238),
.Y(n_4293)
);

OR2x2_ASAP7_75t_L g4294 ( 
.A(n_4201),
.B(n_4157),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4204),
.B(n_239),
.Y(n_4295)
);

NOR2xp33_ASAP7_75t_L g4296 ( 
.A(n_4181),
.B(n_239),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4176),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4160),
.Y(n_4298)
);

NOR2xp33_ASAP7_75t_L g4299 ( 
.A(n_4138),
.B(n_240),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4180),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4218),
.B(n_240),
.Y(n_4301)
);

OR2x2_ASAP7_75t_L g4302 ( 
.A(n_4162),
.B(n_241),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4232),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4184),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4187),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4195),
.Y(n_4306)
);

NOR3xp33_ASAP7_75t_L g4307 ( 
.A(n_4183),
.B(n_241),
.C(n_242),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4161),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_4219),
.B(n_243),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4141),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_4241),
.B(n_243),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4174),
.B(n_244),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_4159),
.B(n_244),
.Y(n_4313)
);

INVxp67_ASAP7_75t_L g4314 ( 
.A(n_4207),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4179),
.B(n_246),
.Y(n_4315)
);

INVxp67_ASAP7_75t_L g4316 ( 
.A(n_4240),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4249),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4163),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4225),
.B(n_246),
.Y(n_4319)
);

NAND2x1_ASAP7_75t_SL g4320 ( 
.A(n_4211),
.B(n_247),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4164),
.Y(n_4321)
);

AND2x2_ASAP7_75t_L g4322 ( 
.A(n_4205),
.B(n_247),
.Y(n_4322)
);

OR2x2_ASAP7_75t_L g4323 ( 
.A(n_4165),
.B(n_248),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4166),
.B(n_248),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4169),
.Y(n_4325)
);

NAND3xp33_ASAP7_75t_L g4326 ( 
.A(n_4239),
.B(n_249),
.C(n_250),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4186),
.B(n_249),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4199),
.B(n_250),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_4226),
.B(n_251),
.Y(n_4329)
);

OAI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_4147),
.A2(n_4175),
.B(n_4168),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4229),
.B(n_251),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4213),
.B(n_252),
.Y(n_4332)
);

AND2x2_ASAP7_75t_L g4333 ( 
.A(n_4177),
.B(n_252),
.Y(n_4333)
);

INVx2_ASAP7_75t_L g4334 ( 
.A(n_4247),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4214),
.B(n_253),
.Y(n_4335)
);

INVxp67_ASAP7_75t_L g4336 ( 
.A(n_4172),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4209),
.Y(n_4337)
);

AND2x2_ASAP7_75t_L g4338 ( 
.A(n_4178),
.B(n_253),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4182),
.B(n_257),
.Y(n_4339)
);

NOR2xp33_ASAP7_75t_L g4340 ( 
.A(n_4223),
.B(n_257),
.Y(n_4340)
);

NOR2xp33_ASAP7_75t_L g4341 ( 
.A(n_4235),
.B(n_258),
.Y(n_4341)
);

INVxp67_ASAP7_75t_L g4342 ( 
.A(n_4233),
.Y(n_4342)
);

XNOR2x1_ASAP7_75t_L g4343 ( 
.A(n_4222),
.B(n_259),
.Y(n_4343)
);

INVx1_ASAP7_75t_SL g4344 ( 
.A(n_4237),
.Y(n_4344)
);

NOR2xp33_ASAP7_75t_L g4345 ( 
.A(n_4248),
.B(n_259),
.Y(n_4345)
);

INVx2_ASAP7_75t_SL g4346 ( 
.A(n_4188),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_4220),
.B(n_260),
.Y(n_4347)
);

NOR2xp33_ASAP7_75t_L g4348 ( 
.A(n_4221),
.B(n_260),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_SL g4349 ( 
.A1(n_4245),
.A2(n_261),
.B(n_262),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4253),
.Y(n_4350)
);

OR2x2_ASAP7_75t_L g4351 ( 
.A(n_4192),
.B(n_261),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4238),
.Y(n_4352)
);

OAI22xp33_ASAP7_75t_L g4353 ( 
.A1(n_4230),
.A2(n_4216),
.B1(n_4236),
.B2(n_4185),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4244),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_4231),
.B(n_262),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4242),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4234),
.Y(n_4357)
);

OAI21xp5_ASAP7_75t_SL g4358 ( 
.A1(n_4194),
.A2(n_263),
.B(n_264),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4200),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4251),
.Y(n_4360)
);

NOR2xp33_ASAP7_75t_L g4361 ( 
.A(n_4196),
.B(n_264),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_4197),
.B(n_265),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4198),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_4190),
.B(n_266),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4246),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4252),
.B(n_267),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4170),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4135),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4135),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4217),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_SL g4371 ( 
.A(n_4135),
.B(n_2198),
.Y(n_4371)
);

OR2x2_ASAP7_75t_L g4372 ( 
.A(n_4135),
.B(n_268),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4135),
.Y(n_4373)
);

AOI21xp33_ASAP7_75t_L g4374 ( 
.A1(n_4167),
.A2(n_268),
.B(n_269),
.Y(n_4374)
);

HB1xp67_ASAP7_75t_L g4375 ( 
.A(n_4212),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4135),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_4143),
.B(n_270),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_4143),
.B(n_270),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4135),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4143),
.B(n_273),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4143),
.B(n_274),
.Y(n_4381)
);

OR2x2_ASAP7_75t_L g4382 ( 
.A(n_4135),
.B(n_275),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4217),
.Y(n_4383)
);

AND2x2_ASAP7_75t_L g4384 ( 
.A(n_4135),
.B(n_277),
.Y(n_4384)
);

NOR2xp33_ASAP7_75t_L g4385 ( 
.A(n_4143),
.B(n_277),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4135),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4135),
.Y(n_4387)
);

INVx2_ASAP7_75t_SL g4388 ( 
.A(n_4135),
.Y(n_4388)
);

OAI22xp5_ASAP7_75t_L g4389 ( 
.A1(n_4140),
.A2(n_281),
.B1(n_278),
.B2(n_279),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_4143),
.B(n_278),
.Y(n_4390)
);

XNOR2xp5_ASAP7_75t_L g4391 ( 
.A(n_4217),
.B(n_282),
.Y(n_4391)
);

HB1xp67_ASAP7_75t_L g4392 ( 
.A(n_4212),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4143),
.B(n_283),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4135),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_4135),
.B(n_286),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4135),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4135),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4135),
.Y(n_4398)
);

OR2x2_ASAP7_75t_L g4399 ( 
.A(n_4135),
.B(n_287),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4135),
.Y(n_4400)
);

NAND2x1_ASAP7_75t_SL g4401 ( 
.A(n_4212),
.B(n_288),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4135),
.B(n_288),
.Y(n_4402)
);

OAI211xp5_ASAP7_75t_L g4403 ( 
.A1(n_4290),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4303),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4388),
.B(n_290),
.Y(n_4405)
);

AOI21xp5_ASAP7_75t_L g4406 ( 
.A1(n_4375),
.A2(n_292),
.B(n_293),
.Y(n_4406)
);

HB1xp67_ASAP7_75t_L g4407 ( 
.A(n_4280),
.Y(n_4407)
);

NOR2xp33_ASAP7_75t_L g4408 ( 
.A(n_4392),
.B(n_292),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4401),
.B(n_296),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4320),
.B(n_297),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4391),
.Y(n_4411)
);

NOR2xp67_ASAP7_75t_L g4412 ( 
.A(n_4368),
.B(n_298),
.Y(n_4412)
);

AOI32xp33_ASAP7_75t_L g4413 ( 
.A1(n_4263),
.A2(n_301),
.A3(n_298),
.B1(n_300),
.B2(n_302),
.Y(n_4413)
);

A2O1A1Ixp33_ASAP7_75t_L g4414 ( 
.A1(n_4385),
.A2(n_304),
.B(n_300),
.C(n_303),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4313),
.Y(n_4415)
);

OAI221xp5_ASAP7_75t_L g4416 ( 
.A1(n_4330),
.A2(n_306),
.B1(n_303),
.B2(n_305),
.C(n_307),
.Y(n_4416)
);

NAND4xp25_ASAP7_75t_L g4417 ( 
.A(n_4369),
.B(n_309),
.C(n_307),
.D(n_308),
.Y(n_4417)
);

NAND4xp25_ASAP7_75t_L g4418 ( 
.A(n_4373),
.B(n_311),
.C(n_308),
.D(n_309),
.Y(n_4418)
);

NOR3xp33_ASAP7_75t_L g4419 ( 
.A(n_4275),
.B(n_312),
.C(n_313),
.Y(n_4419)
);

NOR3xp33_ASAP7_75t_L g4420 ( 
.A(n_4329),
.B(n_312),
.C(n_313),
.Y(n_4420)
);

AND2x2_ASAP7_75t_L g4421 ( 
.A(n_4402),
.B(n_314),
.Y(n_4421)
);

BUFx2_ASAP7_75t_L g4422 ( 
.A(n_4376),
.Y(n_4422)
);

NOR3xp33_ASAP7_75t_L g4423 ( 
.A(n_4377),
.B(n_4380),
.C(n_4378),
.Y(n_4423)
);

OAI221xp5_ASAP7_75t_L g4424 ( 
.A1(n_4316),
.A2(n_4277),
.B1(n_4264),
.B2(n_4257),
.C(n_4298),
.Y(n_4424)
);

NAND3xp33_ASAP7_75t_SL g4425 ( 
.A(n_4370),
.B(n_315),
.C(n_316),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_4383),
.B(n_316),
.Y(n_4426)
);

NAND3xp33_ASAP7_75t_L g4427 ( 
.A(n_4379),
.B(n_318),
.C(n_319),
.Y(n_4427)
);

NOR2xp33_ASAP7_75t_L g4428 ( 
.A(n_4261),
.B(n_319),
.Y(n_4428)
);

NOR3xp33_ASAP7_75t_SL g4429 ( 
.A(n_4386),
.B(n_320),
.C(n_321),
.Y(n_4429)
);

NAND4xp75_ASAP7_75t_L g4430 ( 
.A(n_4273),
.B(n_327),
.C(n_322),
.D(n_323),
.Y(n_4430)
);

NAND3xp33_ASAP7_75t_L g4431 ( 
.A(n_4387),
.B(n_322),
.C(n_323),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4394),
.Y(n_4432)
);

NOR2xp33_ASAP7_75t_L g4433 ( 
.A(n_4396),
.B(n_4397),
.Y(n_4433)
);

AOI211xp5_ASAP7_75t_L g4434 ( 
.A1(n_4272),
.A2(n_330),
.B(n_327),
.C(n_329),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4398),
.Y(n_4435)
);

INVx1_ASAP7_75t_SL g4436 ( 
.A(n_4384),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_4395),
.B(n_329),
.Y(n_4437)
);

NOR3x1_ASAP7_75t_L g4438 ( 
.A(n_4358),
.B(n_330),
.C(n_331),
.Y(n_4438)
);

AOI22xp33_ASAP7_75t_L g4439 ( 
.A1(n_4288),
.A2(n_2255),
.B1(n_2268),
.B2(n_2228),
.Y(n_4439)
);

NOR3x1_ASAP7_75t_SL g4440 ( 
.A(n_4400),
.B(n_331),
.C(n_332),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4259),
.B(n_333),
.Y(n_4441)
);

NAND4xp25_ASAP7_75t_L g4442 ( 
.A(n_4276),
.B(n_339),
.C(n_335),
.D(n_337),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4291),
.B(n_337),
.Y(n_4443)
);

AOI21xp5_ASAP7_75t_L g4444 ( 
.A1(n_4282),
.A2(n_339),
.B(n_340),
.Y(n_4444)
);

NOR2xp33_ASAP7_75t_SL g4445 ( 
.A(n_4294),
.B(n_340),
.Y(n_4445)
);

NOR3xp33_ASAP7_75t_L g4446 ( 
.A(n_4381),
.B(n_341),
.C(n_343),
.Y(n_4446)
);

AOI21xp5_ASAP7_75t_L g4447 ( 
.A1(n_4390),
.A2(n_341),
.B(n_343),
.Y(n_4447)
);

NAND2xp33_ASAP7_75t_L g4448 ( 
.A(n_4372),
.B(n_344),
.Y(n_4448)
);

AOI211xp5_ASAP7_75t_L g4449 ( 
.A1(n_4311),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4285),
.B(n_345),
.Y(n_4450)
);

NAND4xp75_ASAP7_75t_L g4451 ( 
.A(n_4256),
.B(n_350),
.C(n_347),
.D(n_348),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4262),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4289),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_SL g4454 ( 
.A(n_4346),
.B(n_2228),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_4268),
.B(n_347),
.Y(n_4455)
);

NOR3x1_ASAP7_75t_L g4456 ( 
.A(n_4349),
.B(n_350),
.C(n_351),
.Y(n_4456)
);

AOI221xp5_ASAP7_75t_L g4457 ( 
.A1(n_4318),
.A2(n_4321),
.B1(n_4325),
.B2(n_4353),
.C(n_4352),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4269),
.B(n_351),
.Y(n_4458)
);

INVxp67_ASAP7_75t_L g4459 ( 
.A(n_4382),
.Y(n_4459)
);

AND3x1_ASAP7_75t_L g4460 ( 
.A(n_4255),
.B(n_352),
.C(n_353),
.Y(n_4460)
);

CKINVDCx5p33_ASAP7_75t_R g4461 ( 
.A(n_4344),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4292),
.Y(n_4462)
);

AOI321xp33_ASAP7_75t_L g4463 ( 
.A1(n_4365),
.A2(n_355),
.A3(n_357),
.B1(n_352),
.B2(n_353),
.C(n_356),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4319),
.Y(n_4464)
);

NAND3xp33_ASAP7_75t_L g4465 ( 
.A(n_4287),
.B(n_4299),
.C(n_4361),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4322),
.Y(n_4466)
);

NOR2xp33_ASAP7_75t_L g4467 ( 
.A(n_4399),
.B(n_355),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4302),
.Y(n_4468)
);

OR2x2_ASAP7_75t_L g4469 ( 
.A(n_4284),
.B(n_356),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4266),
.B(n_358),
.Y(n_4470)
);

NOR2xp33_ASAP7_75t_L g4471 ( 
.A(n_4297),
.B(n_358),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4270),
.B(n_359),
.Y(n_4472)
);

NAND4xp25_ASAP7_75t_L g4473 ( 
.A(n_4279),
.B(n_362),
.C(n_360),
.D(n_361),
.Y(n_4473)
);

NAND3xp33_ASAP7_75t_L g4474 ( 
.A(n_4260),
.B(n_362),
.C(n_363),
.Y(n_4474)
);

NAND3xp33_ASAP7_75t_L g4475 ( 
.A(n_4307),
.B(n_364),
.C(n_365),
.Y(n_4475)
);

XNOR2xp5_ASAP7_75t_L g4476 ( 
.A(n_4343),
.B(n_364),
.Y(n_4476)
);

OAI21xp33_ASAP7_75t_L g4477 ( 
.A1(n_4254),
.A2(n_365),
.B(n_366),
.Y(n_4477)
);

NOR2x1_ASAP7_75t_L g4478 ( 
.A(n_4354),
.B(n_367),
.Y(n_4478)
);

NOR4xp25_ASAP7_75t_L g4479 ( 
.A(n_4317),
.B(n_369),
.C(n_367),
.D(n_368),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4283),
.Y(n_4480)
);

NOR3xp33_ASAP7_75t_L g4481 ( 
.A(n_4393),
.B(n_370),
.C(n_371),
.Y(n_4481)
);

AND2x2_ASAP7_75t_L g4482 ( 
.A(n_4357),
.B(n_370),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_SL g4483 ( 
.A(n_4324),
.B(n_2255),
.Y(n_4483)
);

OAI21xp5_ASAP7_75t_L g4484 ( 
.A1(n_4326),
.A2(n_371),
.B(n_372),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4323),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4333),
.Y(n_4486)
);

AND2x4_ASAP7_75t_L g4487 ( 
.A(n_4338),
.B(n_372),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_4339),
.B(n_373),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4362),
.B(n_376),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_4351),
.Y(n_4490)
);

AOI322xp5_ASAP7_75t_L g4491 ( 
.A1(n_4407),
.A2(n_4337),
.A3(n_4360),
.B1(n_4308),
.B2(n_4356),
.C1(n_4305),
.C2(n_4304),
.Y(n_4491)
);

AOI21xp33_ASAP7_75t_SL g4492 ( 
.A1(n_4461),
.A2(n_4404),
.B(n_4408),
.Y(n_4492)
);

AOI21xp5_ASAP7_75t_L g4493 ( 
.A1(n_4422),
.A2(n_4355),
.B(n_4295),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_4433),
.A2(n_4274),
.B(n_4278),
.Y(n_4494)
);

AOI22xp5_ASAP7_75t_L g4495 ( 
.A1(n_4452),
.A2(n_4359),
.B1(n_4341),
.B2(n_4348),
.Y(n_4495)
);

OAI211xp5_ASAP7_75t_L g4496 ( 
.A1(n_4432),
.A2(n_4363),
.B(n_4258),
.C(n_4271),
.Y(n_4496)
);

AOI211xp5_ASAP7_75t_L g4497 ( 
.A1(n_4424),
.A2(n_4314),
.B(n_4374),
.C(n_4267),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4440),
.Y(n_4498)
);

AOI221xp5_ASAP7_75t_L g4499 ( 
.A1(n_4457),
.A2(n_4265),
.B1(n_4336),
.B2(n_4342),
.C(n_4306),
.Y(n_4499)
);

AOI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4468),
.A2(n_4345),
.B1(n_4310),
.B2(n_4334),
.Y(n_4500)
);

NOR2x1_ASAP7_75t_L g4501 ( 
.A(n_4405),
.B(n_4389),
.Y(n_4501)
);

AND2x4_ASAP7_75t_L g4502 ( 
.A(n_4435),
.B(n_4300),
.Y(n_4502)
);

INVx2_ASAP7_75t_SL g4503 ( 
.A(n_4441),
.Y(n_4503)
);

OAI211xp5_ASAP7_75t_SL g4504 ( 
.A1(n_4436),
.A2(n_4350),
.B(n_4367),
.C(n_4347),
.Y(n_4504)
);

AOI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_4423),
.A2(n_4340),
.B1(n_4309),
.B2(n_4301),
.Y(n_4505)
);

O2A1O1Ixp33_ASAP7_75t_L g4506 ( 
.A1(n_4448),
.A2(n_4364),
.B(n_4335),
.C(n_4332),
.Y(n_4506)
);

AOI322xp5_ASAP7_75t_L g4507 ( 
.A1(n_4478),
.A2(n_4312),
.A3(n_4327),
.B1(n_4328),
.B2(n_4315),
.C1(n_4286),
.C2(n_4331),
.Y(n_4507)
);

AOI221x1_ASAP7_75t_L g4508 ( 
.A1(n_4420),
.A2(n_4296),
.B1(n_4366),
.B2(n_4293),
.C(n_4371),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4487),
.B(n_4281),
.Y(n_4509)
);

AOI221xp5_ASAP7_75t_L g4510 ( 
.A1(n_4479),
.A2(n_4281),
.B1(n_380),
.B2(n_377),
.C(n_378),
.Y(n_4510)
);

OAI21xp33_ASAP7_75t_L g4511 ( 
.A1(n_4428),
.A2(n_4445),
.B(n_4459),
.Y(n_4511)
);

OAI221xp5_ASAP7_75t_SL g4512 ( 
.A1(n_4411),
.A2(n_381),
.B1(n_377),
.B2(n_380),
.C(n_382),
.Y(n_4512)
);

NOR3xp33_ASAP7_75t_L g4513 ( 
.A(n_4425),
.B(n_383),
.C(n_384),
.Y(n_4513)
);

NOR2xp33_ASAP7_75t_L g4514 ( 
.A(n_4473),
.B(n_4403),
.Y(n_4514)
);

NAND5xp2_ASAP7_75t_L g4515 ( 
.A(n_4464),
.B(n_385),
.C(n_383),
.D(n_384),
.E(n_386),
.Y(n_4515)
);

NOR3x1_ASAP7_75t_L g4516 ( 
.A(n_4416),
.B(n_387),
.C(n_388),
.Y(n_4516)
);

OAI22xp5_ASAP7_75t_L g4517 ( 
.A1(n_4434),
.A2(n_396),
.B1(n_390),
.B2(n_393),
.Y(n_4517)
);

INVxp67_ASAP7_75t_L g4518 ( 
.A(n_4460),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4476),
.Y(n_4519)
);

INVx3_ASAP7_75t_SL g4520 ( 
.A(n_4469),
.Y(n_4520)
);

INVxp67_ASAP7_75t_L g4521 ( 
.A(n_4412),
.Y(n_4521)
);

AND4x2_ASAP7_75t_L g4522 ( 
.A(n_4444),
.B(n_397),
.C(n_390),
.D(n_396),
.Y(n_4522)
);

AOI22xp5_ASAP7_75t_L g4523 ( 
.A1(n_4466),
.A2(n_4486),
.B1(n_4415),
.B2(n_4462),
.Y(n_4523)
);

AOI221xp5_ASAP7_75t_L g4524 ( 
.A1(n_4453),
.A2(n_400),
.B1(n_397),
.B2(n_398),
.C(n_401),
.Y(n_4524)
);

AOI221xp5_ASAP7_75t_L g4525 ( 
.A1(n_4465),
.A2(n_406),
.B1(n_403),
.B2(n_404),
.C(n_407),
.Y(n_4525)
);

OAI211xp5_ASAP7_75t_SL g4526 ( 
.A1(n_4480),
.A2(n_407),
.B(n_404),
.C(n_406),
.Y(n_4526)
);

AOI211xp5_ASAP7_75t_L g4527 ( 
.A1(n_4484),
.A2(n_412),
.B(n_408),
.C(n_410),
.Y(n_4527)
);

OAI221xp5_ASAP7_75t_L g4528 ( 
.A1(n_4455),
.A2(n_413),
.B1(n_408),
.B2(n_410),
.C(n_414),
.Y(n_4528)
);

AOI221xp5_ASAP7_75t_L g4529 ( 
.A1(n_4485),
.A2(n_416),
.B1(n_413),
.B2(n_415),
.C(n_419),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4487),
.B(n_419),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4470),
.Y(n_4531)
);

AOI21xp33_ASAP7_75t_L g4532 ( 
.A1(n_4490),
.A2(n_420),
.B(n_422),
.Y(n_4532)
);

NOR2xp33_ASAP7_75t_R g4533 ( 
.A(n_4421),
.B(n_420),
.Y(n_4533)
);

AOI221xp5_ASAP7_75t_L g4534 ( 
.A1(n_4426),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.C(n_426),
.Y(n_4534)
);

AOI222xp33_ASAP7_75t_L g4535 ( 
.A1(n_4472),
.A2(n_429),
.B1(n_431),
.B2(n_424),
.C1(n_427),
.C2(n_430),
.Y(n_4535)
);

AOI21xp5_ASAP7_75t_L g4536 ( 
.A1(n_4406),
.A2(n_429),
.B(n_430),
.Y(n_4536)
);

XOR2x2_ASAP7_75t_L g4537 ( 
.A(n_4430),
.B(n_433),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4489),
.Y(n_4538)
);

AOI22xp33_ASAP7_75t_SL g4539 ( 
.A1(n_4471),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_4539)
);

OAI21xp33_ASAP7_75t_L g4540 ( 
.A1(n_4458),
.A2(n_434),
.B(n_435),
.Y(n_4540)
);

OAI222xp33_ASAP7_75t_L g4541 ( 
.A1(n_4409),
.A2(n_438),
.B1(n_440),
.B2(n_436),
.C1(n_437),
.C2(n_439),
.Y(n_4541)
);

OAI221xp5_ASAP7_75t_L g4542 ( 
.A1(n_4477),
.A2(n_441),
.B1(n_436),
.B2(n_439),
.C(n_444),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4429),
.B(n_445),
.Y(n_4543)
);

NOR2xp33_ASAP7_75t_R g4544 ( 
.A(n_4437),
.B(n_446),
.Y(n_4544)
);

AOI211xp5_ASAP7_75t_L g4545 ( 
.A1(n_4474),
.A2(n_449),
.B(n_446),
.C(n_447),
.Y(n_4545)
);

OAI22xp5_ASAP7_75t_L g4546 ( 
.A1(n_4427),
.A2(n_450),
.B1(n_447),
.B2(n_449),
.Y(n_4546)
);

AOI211xp5_ASAP7_75t_SL g4547 ( 
.A1(n_4467),
.A2(n_453),
.B(n_450),
.C(n_452),
.Y(n_4547)
);

AOI32xp33_ASAP7_75t_L g4548 ( 
.A1(n_4482),
.A2(n_454),
.A3(n_452),
.B1(n_453),
.B2(n_456),
.Y(n_4548)
);

AOI222xp33_ASAP7_75t_L g4549 ( 
.A1(n_4498),
.A2(n_4510),
.B1(n_4518),
.B2(n_4521),
.C1(n_4509),
.C2(n_4520),
.Y(n_4549)
);

AOI22xp5_ASAP7_75t_L g4550 ( 
.A1(n_4514),
.A2(n_4446),
.B1(n_4481),
.B2(n_4410),
.Y(n_4550)
);

AOI322xp5_ASAP7_75t_L g4551 ( 
.A1(n_4501),
.A2(n_4450),
.A3(n_4419),
.B1(n_4443),
.B2(n_4488),
.C1(n_4439),
.C2(n_4414),
.Y(n_4551)
);

NAND3xp33_ASAP7_75t_SL g4552 ( 
.A(n_4497),
.B(n_4449),
.C(n_4447),
.Y(n_4552)
);

OAI21xp33_ASAP7_75t_L g4553 ( 
.A1(n_4496),
.A2(n_4418),
.B(n_4417),
.Y(n_4553)
);

OAI221xp5_ASAP7_75t_L g4554 ( 
.A1(n_4511),
.A2(n_4513),
.B1(n_4523),
.B2(n_4492),
.C(n_4493),
.Y(n_4554)
);

AOI221xp5_ASAP7_75t_SL g4555 ( 
.A1(n_4499),
.A2(n_4454),
.B1(n_4442),
.B2(n_4483),
.C(n_4438),
.Y(n_4555)
);

OAI21xp5_ASAP7_75t_L g4556 ( 
.A1(n_4494),
.A2(n_4431),
.B(n_4475),
.Y(n_4556)
);

AOI22xp5_ASAP7_75t_L g4557 ( 
.A1(n_4503),
.A2(n_4451),
.B1(n_4456),
.B2(n_4463),
.Y(n_4557)
);

AO221x1_ASAP7_75t_L g4558 ( 
.A1(n_4517),
.A2(n_4413),
.B1(n_460),
.B2(n_457),
.C(n_458),
.Y(n_4558)
);

AOI321xp33_ASAP7_75t_L g4559 ( 
.A1(n_4519),
.A2(n_4502),
.A3(n_4531),
.B1(n_4538),
.B2(n_4500),
.C(n_4495),
.Y(n_4559)
);

OAI22xp5_ASAP7_75t_L g4560 ( 
.A1(n_4502),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4491),
.B(n_462),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4522),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4516),
.B(n_4539),
.Y(n_4563)
);

HB1xp67_ASAP7_75t_L g4564 ( 
.A(n_4533),
.Y(n_4564)
);

OAI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4536),
.A2(n_463),
.B(n_464),
.Y(n_4565)
);

NOR3xp33_ASAP7_75t_L g4566 ( 
.A(n_4504),
.B(n_464),
.C(n_465),
.Y(n_4566)
);

AOI221xp5_ASAP7_75t_L g4567 ( 
.A1(n_4506),
.A2(n_468),
.B1(n_465),
.B2(n_467),
.C(n_469),
.Y(n_4567)
);

OAI221xp5_ASAP7_75t_L g4568 ( 
.A1(n_4527),
.A2(n_470),
.B1(n_467),
.B2(n_468),
.C(n_471),
.Y(n_4568)
);

OAI21xp33_ASAP7_75t_L g4569 ( 
.A1(n_4507),
.A2(n_470),
.B(n_472),
.Y(n_4569)
);

AOI221xp5_ASAP7_75t_L g4570 ( 
.A1(n_4540),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.C(n_475),
.Y(n_4570)
);

AOI221xp5_ASAP7_75t_L g4571 ( 
.A1(n_4546),
.A2(n_479),
.B1(n_475),
.B2(n_478),
.C(n_481),
.Y(n_4571)
);

OAI22xp5_ASAP7_75t_L g4572 ( 
.A1(n_4528),
.A2(n_482),
.B1(n_479),
.B2(n_481),
.Y(n_4572)
);

OA22x2_ASAP7_75t_L g4573 ( 
.A1(n_4505),
.A2(n_4508),
.B1(n_4543),
.B2(n_4530),
.Y(n_4573)
);

NAND3xp33_ASAP7_75t_SL g4574 ( 
.A(n_4544),
.B(n_483),
.C(n_487),
.Y(n_4574)
);

OAI211xp5_ASAP7_75t_L g4575 ( 
.A1(n_4525),
.A2(n_491),
.B(n_489),
.C(n_490),
.Y(n_4575)
);

OAI221xp5_ASAP7_75t_R g4576 ( 
.A1(n_4537),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.C(n_495),
.Y(n_4576)
);

AOI221xp5_ASAP7_75t_L g4577 ( 
.A1(n_4542),
.A2(n_496),
.B1(n_492),
.B2(n_493),
.C(n_497),
.Y(n_4577)
);

AO21x1_ASAP7_75t_L g4578 ( 
.A1(n_4545),
.A2(n_496),
.B(n_497),
.Y(n_4578)
);

AOI22xp33_ASAP7_75t_L g4579 ( 
.A1(n_4526),
.A2(n_2281),
.B1(n_2283),
.B2(n_2268),
.Y(n_4579)
);

HB1xp67_ASAP7_75t_L g4580 ( 
.A(n_4547),
.Y(n_4580)
);

AOI211x1_ASAP7_75t_SL g4581 ( 
.A1(n_4532),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_4581)
);

NOR2x1_ASAP7_75t_L g4582 ( 
.A(n_4541),
.B(n_500),
.Y(n_4582)
);

NOR2x1_ASAP7_75t_L g4583 ( 
.A(n_4515),
.B(n_4512),
.Y(n_4583)
);

INVx1_ASAP7_75t_SL g4584 ( 
.A(n_4580),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4564),
.Y(n_4585)
);

NOR4xp25_ASAP7_75t_L g4586 ( 
.A(n_4554),
.B(n_4548),
.C(n_4534),
.D(n_4524),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4562),
.Y(n_4587)
);

AOI22xp33_ASAP7_75t_L g4588 ( 
.A1(n_4573),
.A2(n_4535),
.B1(n_4529),
.B2(n_2283),
.Y(n_4588)
);

OAI31xp33_ASAP7_75t_L g4589 ( 
.A1(n_4575),
.A2(n_506),
.A3(n_501),
.B(n_505),
.Y(n_4589)
);

AOI221xp5_ASAP7_75t_L g4590 ( 
.A1(n_4553),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.C(n_508),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4582),
.Y(n_4591)
);

AND2x4_ASAP7_75t_L g4592 ( 
.A(n_4583),
.B(n_507),
.Y(n_4592)
);

AOI22xp5_ASAP7_75t_L g4593 ( 
.A1(n_4549),
.A2(n_2287),
.B1(n_2296),
.B2(n_2281),
.Y(n_4593)
);

NOR4xp75_ASAP7_75t_L g4594 ( 
.A(n_4556),
.B(n_510),
.C(n_508),
.D(n_509),
.Y(n_4594)
);

AOI21xp5_ASAP7_75t_L g4595 ( 
.A1(n_4560),
.A2(n_509),
.B(n_510),
.Y(n_4595)
);

NOR2xp33_ASAP7_75t_L g4596 ( 
.A(n_4574),
.B(n_4557),
.Y(n_4596)
);

NOR3xp33_ASAP7_75t_L g4597 ( 
.A(n_4561),
.B(n_511),
.C(n_512),
.Y(n_4597)
);

AOI22xp5_ASAP7_75t_L g4598 ( 
.A1(n_4550),
.A2(n_4552),
.B1(n_4563),
.B2(n_4566),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4581),
.B(n_511),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4578),
.Y(n_4600)
);

O2A1O1Ixp33_ASAP7_75t_L g4601 ( 
.A1(n_4569),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4600),
.B(n_4558),
.Y(n_4602)
);

NOR2xp67_ASAP7_75t_L g4603 ( 
.A(n_4585),
.B(n_4568),
.Y(n_4603)
);

BUFx2_ASAP7_75t_L g4604 ( 
.A(n_4591),
.Y(n_4604)
);

AND2x4_ASAP7_75t_L g4605 ( 
.A(n_4584),
.B(n_4565),
.Y(n_4605)
);

OAI221xp5_ASAP7_75t_SL g4606 ( 
.A1(n_4598),
.A2(n_4559),
.B1(n_4551),
.B2(n_4555),
.C(n_4577),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4592),
.B(n_4570),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4594),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4586),
.B(n_4567),
.Y(n_4609)
);

OAI22xp5_ASAP7_75t_L g4610 ( 
.A1(n_4587),
.A2(n_4572),
.B1(n_4571),
.B2(n_4579),
.Y(n_4610)
);

AND2x4_ASAP7_75t_SL g4611 ( 
.A(n_4596),
.B(n_4576),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4599),
.Y(n_4612)
);

OR2x2_ASAP7_75t_L g4613 ( 
.A(n_4589),
.B(n_513),
.Y(n_4613)
);

HB1xp67_ASAP7_75t_L g4614 ( 
.A(n_4604),
.Y(n_4614)
);

HB1xp67_ASAP7_75t_L g4615 ( 
.A(n_4608),
.Y(n_4615)
);

CKINVDCx14_ASAP7_75t_R g4616 ( 
.A(n_4609),
.Y(n_4616)
);

NAND4xp25_ASAP7_75t_L g4617 ( 
.A(n_4606),
.B(n_4597),
.C(n_4601),
.D(n_4588),
.Y(n_4617)
);

BUFx6f_ASAP7_75t_L g4618 ( 
.A(n_4605),
.Y(n_4618)
);

HB1xp67_ASAP7_75t_L g4619 ( 
.A(n_4602),
.Y(n_4619)
);

CKINVDCx5p33_ASAP7_75t_R g4620 ( 
.A(n_4611),
.Y(n_4620)
);

CKINVDCx5p33_ASAP7_75t_R g4621 ( 
.A(n_4612),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4613),
.Y(n_4622)
);

AOI22xp33_ASAP7_75t_L g4623 ( 
.A1(n_4616),
.A2(n_4607),
.B1(n_4603),
.B2(n_4610),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4618),
.Y(n_4624)
);

OAI22xp5_ASAP7_75t_SL g4625 ( 
.A1(n_4620),
.A2(n_4593),
.B1(n_4590),
.B2(n_4595),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4614),
.B(n_516),
.Y(n_4626)
);

OAI22xp5_ASAP7_75t_SL g4627 ( 
.A1(n_4623),
.A2(n_4621),
.B1(n_4619),
.B2(n_4618),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4624),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4626),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4627),
.Y(n_4630)
);

HB1xp67_ASAP7_75t_L g4631 ( 
.A(n_4630),
.Y(n_4631)
);

XOR2xp5_ASAP7_75t_L g4632 ( 
.A(n_4631),
.B(n_4615),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4632),
.Y(n_4633)
);

AOI22xp33_ASAP7_75t_L g4634 ( 
.A1(n_4633),
.A2(n_4628),
.B1(n_4622),
.B2(n_4629),
.Y(n_4634)
);

AOI22xp5_ASAP7_75t_L g4635 ( 
.A1(n_4634),
.A2(n_4617),
.B1(n_4625),
.B2(n_522),
.Y(n_4635)
);

AOI21xp33_ASAP7_75t_SL g4636 ( 
.A1(n_4635),
.A2(n_517),
.B(n_518),
.Y(n_4636)
);

NAND3xp33_ASAP7_75t_SL g4637 ( 
.A(n_4636),
.B(n_522),
.C(n_523),
.Y(n_4637)
);

AOI211xp5_ASAP7_75t_L g4638 ( 
.A1(n_4637),
.A2(n_2298),
.B(n_2297),
.C(n_525),
.Y(n_4638)
);


endmodule