module real_jpeg_25199_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_40),
.B1(n_68),
.B2(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_1),
.A2(n_40),
.B1(n_55),
.B2(n_63),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_1),
.A2(n_23),
.B1(n_28),
.B2(n_40),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_23),
.B1(n_28),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_3),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_68),
.B1(n_70),
.B2(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_36),
.B1(n_41),
.B2(n_97),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_3),
.A2(n_55),
.B1(n_63),
.B2(n_97),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_5),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_23),
.B1(n_28),
.B2(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_5),
.A2(n_68),
.B1(n_70),
.B2(n_83),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_55),
.B1(n_63),
.B2(n_83),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_7),
.A2(n_124),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_7),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_7),
.A2(n_23),
.B1(n_28),
.B2(n_173),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_7),
.A2(n_68),
.B1(n_70),
.B2(n_173),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_7),
.A2(n_55),
.B1(n_63),
.B2(n_173),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_23),
.B1(n_28),
.B2(n_67),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_8),
.A2(n_42),
.B1(n_67),
.B2(n_122),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_8),
.A2(n_55),
.B1(n_63),
.B2(n_67),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_11),
.A2(n_32),
.B1(n_42),
.B2(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_11),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_11),
.A2(n_23),
.B1(n_28),
.B2(n_87),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_68),
.B1(n_70),
.B2(n_87),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_11),
.A2(n_55),
.B1(n_63),
.B2(n_87),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_12),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_12),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_12),
.A2(n_23),
.B1(n_28),
.B2(n_121),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_12),
.A2(n_68),
.B1(n_70),
.B2(n_121),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_12),
.A2(n_55),
.B1(n_63),
.B2(n_121),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_13),
.B(n_36),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_13),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_13),
.B(n_22),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_68),
.C(n_93),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_13),
.A2(n_23),
.B1(n_28),
.B2(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_13),
.B(n_139),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_13),
.A2(n_68),
.B1(n_70),
.B2(n_225),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_13),
.B(n_55),
.C(n_73),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_13),
.A2(n_54),
.B(n_285),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_15),
.A2(n_35),
.B1(n_55),
.B2(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_15),
.A2(n_35),
.B1(n_68),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_15),
.A2(n_23),
.B1(n_28),
.B2(n_35),
.Y(n_161)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_16),
.B(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_16),
.Y(n_299)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_44),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_34),
.Y(n_21)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_29),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_22),
.A2(n_29),
.B1(n_120),
.B2(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_22),
.A2(n_29),
.B1(n_39),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_22)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_23),
.A2(n_28),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_23),
.B(n_27),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_23),
.B(n_251),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g195 ( 
.A1(n_26),
.A2(n_28),
.A3(n_122),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_29),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_29),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_29),
.A2(n_127),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_31),
.Y(n_124)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_33),
.A2(n_82),
.B(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_33),
.B(n_86),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_33),
.A2(n_82),
.B1(n_125),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_33),
.A2(n_125),
.B1(n_147),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_33),
.A2(n_84),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_38),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_38),
.B(n_358),
.Y(n_359)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_357),
.B(n_359),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_345),
.B(n_356),
.Y(n_47)
);

OAI31xp33_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_149),
.A3(n_163),
.B(n_342),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_128),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_50),
.B(n_128),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_88),
.C(n_104),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_51),
.A2(n_88),
.B1(n_89),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_51),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_78),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_52),
.A2(n_53),
.B(n_80),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_53),
.A2(n_64),
.B1(n_65),
.B2(n_79),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_59),
.B(n_62),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_62),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_54),
.A2(n_109),
.B1(n_110),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_54),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_54),
.A2(n_201),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_54),
.B(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_54),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_63),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_56),
.Y(n_202)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_61),
.B(n_225),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_63),
.B(n_310),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_71),
.B1(n_77),
.B2(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_70),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_68),
.B(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_71),
.A2(n_77),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_71),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_71),
.A2(n_77),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_75),
.A2(n_100),
.B1(n_115),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_75),
.A2(n_184),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_75),
.A2(n_221),
.B(n_258),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_75),
.B(n_225),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_77),
.B(n_222),
.Y(n_273)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_103),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_91),
.A2(n_92),
.B1(n_141),
.B2(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_91),
.A2(n_191),
.B(n_193),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_91),
.A2(n_193),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_92),
.A2(n_117),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_92),
.A2(n_177),
.B(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_100),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_100),
.A2(n_273),
.B(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_102),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_104),
.A2(n_105),
.B1(n_337),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.C(n_118),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_106),
.A2(n_107),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_108),
.A2(n_112),
.B1(n_113),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_116),
.B(n_118),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_125),
.B(n_126),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_122),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_131),
.C(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_146),
.B2(n_148),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_143),
.C(n_146),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_138),
.A2(n_139),
.B1(n_192),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_138),
.A2(n_139),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_178),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_143),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_143),
.B(n_156),
.C(n_160),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_146),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_148),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_146),
.B(n_152),
.C(n_155),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_150),
.A2(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_162),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_151),
.B(n_162),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_157),
.Y(n_352)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_161),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_335),
.B(n_341),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_210),
.B(n_334),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_203),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_166),
.B(n_203),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_185),
.C(n_187),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_167),
.A2(n_168),
.B1(n_185),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_175),
.C(n_179),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_183),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_185),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_187),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_194),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_190),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_194),
.B(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_198),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_199),
.A2(n_296),
.B1(n_298),
.B2(n_300),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_202),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_205),
.B(n_206),
.C(n_209),
.Y(n_340)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_243),
.B(n_328),
.C(n_333),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_237),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_227),
.C(n_228),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_213),
.A2(n_214),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_219),
.C(n_223),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_227),
.B(n_228),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_233),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_322),
.B(n_327),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_274),
.B(n_321),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_263),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_248),
.B(n_263),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.C(n_260),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_256),
.A2(n_260),
.B1(n_261),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_270),
.C(n_271),
.Y(n_326)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_315),
.B(n_320),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_293),
.B(n_314),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_287),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_287),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_319)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_284),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_291),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_303),
.B(n_313),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_301),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_301),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_299),
.B(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_308),
.B(n_312),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_340),
.Y(n_341)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_347),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_351),
.B1(n_353),
.B2(n_354),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_349),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_351),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_353),
.C(n_355),
.Y(n_358)
);


endmodule