module fake_jpeg_977_n_314 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_48),
.Y(n_133)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_52),
.Y(n_100)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_72),
.Y(n_98)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_57),
.B(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_17),
.B(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_21),
.B(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_37),
.Y(n_104)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_18),
.B(n_7),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_76),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_67),
.Y(n_130)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_18),
.B(n_7),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_11),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_88),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_79),
.B(n_82),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_31),
.B1(n_28),
.B2(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_25),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_84),
.Y(n_112)
);

CKINVDCx9p33_ASAP7_75t_R g84 ( 
.A(n_30),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_89),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_33),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_38),
.B1(n_34),
.B2(n_45),
.Y(n_94)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_94),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_34),
.B1(n_43),
.B2(n_37),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_95),
.A2(n_114),
.B1(n_118),
.B2(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_104),
.B(n_99),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_67),
.A2(n_33),
.B1(n_27),
.B2(n_40),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_111),
.A2(n_120),
.B1(n_132),
.B2(n_140),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_31),
.B1(n_28),
.B2(n_40),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_5),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_122),
.B(n_139),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_129),
.B1(n_131),
.B2(n_108),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_75),
.A2(n_6),
.B1(n_13),
.B2(n_14),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_78),
.A2(n_13),
.B1(n_15),
.B2(n_1),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_61),
.A2(n_1),
.B1(n_15),
.B2(n_91),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_88),
.B1(n_70),
.B2(n_51),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_79),
.B(n_85),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_64),
.B1(n_71),
.B2(n_63),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_57),
.A2(n_58),
.B1(n_66),
.B2(n_42),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_138),
.B1(n_127),
.B2(n_125),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_144),
.B(n_152),
.Y(n_198)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_112),
.B1(n_108),
.B2(n_117),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_146),
.A2(n_148),
.B1(n_147),
.B2(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_96),
.B(n_136),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_152),
.B(n_157),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_165),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_100),
.A2(n_129),
.B(n_123),
.C(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_156),
.B(n_167),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_161),
.Y(n_192)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_105),
.B1(n_109),
.B2(n_150),
.Y(n_185)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_134),
.B1(n_93),
.B2(n_97),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_180),
.B1(n_105),
.B2(n_109),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_121),
.B(n_116),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_97),
.B(n_116),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_125),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_110),
.B(n_128),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_177),
.Y(n_201)
);

OA22x2_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_107),
.B1(n_93),
.B2(n_127),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_176),
.A3(n_105),
.B1(n_152),
.B2(n_171),
.Y(n_195)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_99),
.C(n_107),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_161),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_206),
.B1(n_207),
.B2(n_176),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_172),
.B1(n_174),
.B2(n_180),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_203),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_192),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_151),
.B1(n_162),
.B2(n_154),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_161),
.B1(n_145),
.B2(n_179),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_158),
.B1(n_161),
.B2(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_166),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_196),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_213),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_204),
.B1(n_185),
.B2(n_197),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_153),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_224),
.C(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_178),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_220),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_160),
.C(n_163),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_205),
.B(n_175),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_143),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_143),
.C(n_149),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_159),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_231),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_199),
.B(n_200),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_197),
.B(n_198),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_203),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_246),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_214),
.B1(n_217),
.B2(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_241),
.B(n_249),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_188),
.C(n_194),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_230),
.C(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_195),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_226),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_212),
.B(n_191),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_254),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_253),
.A2(n_234),
.B1(n_236),
.B2(n_238),
.Y(n_268)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_219),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_265),
.Y(n_269)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_243),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_260),
.C(n_267),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_245),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_235),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_209),
.C(n_224),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_211),
.B1(n_216),
.B2(n_221),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_248),
.B1(n_242),
.B2(n_243),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_220),
.B1(n_223),
.B2(n_222),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_242),
.B1(n_235),
.B2(n_239),
.Y(n_279)
);

OAI322xp33_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_199),
.A3(n_200),
.B1(n_181),
.B2(n_187),
.C1(n_202),
.C2(n_193),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_244),
.C(n_238),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_202),
.C(n_181),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_279),
.B1(n_263),
.B2(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_274),
.C(n_265),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_278),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_255),
.B(n_247),
.CI(n_240),
.CON(n_274),
.SN(n_274)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_275),
.A2(n_253),
.B1(n_261),
.B2(n_252),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_249),
.C(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_257),
.C(n_260),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_279),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_262),
.B1(n_255),
.B2(n_239),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_258),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_287),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_262),
.B(n_264),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_286),
.A2(n_278),
.B(n_289),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_271),
.C(n_272),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_259),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_271),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_292),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.C(n_302),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_284),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_296),
.B(n_301),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_281),
.B(n_283),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_294),
.C(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_281),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_305),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_309),
.B(n_275),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_311),
.C(n_270),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_270),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_273),
.Y(n_314)
);


endmodule