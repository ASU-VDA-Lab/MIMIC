module fake_jpeg_17854_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_40),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_30),
.B(n_29),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_28),
.B(n_24),
.C(n_26),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_45),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_55),
.B1(n_58),
.B2(n_54),
.Y(n_69)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_27),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_61),
.B1(n_56),
.B2(n_52),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_81),
.B1(n_84),
.B2(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_16),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_24),
.B(n_26),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_76),
.B(n_50),
.Y(n_88)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_40),
.B1(n_28),
.B2(n_27),
.Y(n_73)
);

AOI22x1_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_74),
.B1(n_22),
.B2(n_25),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_27),
.B1(n_2),
.B2(n_1),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_31),
.B(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_38),
.B1(n_25),
.B2(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_89),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_45),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_97),
.Y(n_120)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_69),
.B1(n_106),
.B2(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_104),
.B1(n_84),
.B2(n_103),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_35),
.CI(n_47),
.CON(n_108),
.SN(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_117),
.B1(n_127),
.B2(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_67),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_73),
.B1(n_68),
.B2(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_64),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_129),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_76),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_80),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_90),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_112),
.B1(n_110),
.B2(n_121),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_88),
.B(n_85),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_138),
.B(n_142),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_148),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_108),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_131),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_152),
.Y(n_168)
);

AO21x2_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_102),
.B(n_94),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_153),
.B1(n_111),
.B2(n_116),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_105),
.B1(n_90),
.B2(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_115),
.C(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_99),
.B1(n_79),
.B2(n_81),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_79),
.B1(n_81),
.B2(n_53),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_113),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_31),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_82),
.B1(n_53),
.B2(n_17),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_145),
.B(n_139),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_157),
.B1(n_161),
.B2(n_164),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_111),
.B1(n_116),
.B2(n_130),
.Y(n_157)
);

XOR2x2_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_82),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_147),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_126),
.B1(n_82),
.B2(n_125),
.Y(n_164)
);

AOI22x1_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_17),
.B1(n_37),
.B2(n_39),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_171),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_126),
.B1(n_125),
.B2(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_72),
.B1(n_109),
.B2(n_125),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_39),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_152),
.C(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_57),
.B1(n_107),
.B2(n_41),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_107),
.B1(n_31),
.B2(n_41),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_173),
.B1(n_140),
.B2(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_146),
.B1(n_134),
.B2(n_136),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_1),
.B(n_2),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_1),
.B(n_2),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_192),
.C(n_160),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_142),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_187),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_144),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_134),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_183),
.B(n_186),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_189),
.B1(n_191),
.B2(n_162),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_133),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_182),
.Y(n_202)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_133),
.B1(n_154),
.B2(n_2),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_191),
.B1(n_178),
.B2(n_184),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_3),
.C(n_4),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_196),
.B1(n_201),
.B2(n_203),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_156),
.B1(n_158),
.B2(n_175),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_160),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_181),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.C(n_197),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_187),
.C(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_164),
.B1(n_171),
.B2(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_174),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_190),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_188),
.B(n_186),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_198),
.B(n_204),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_6),
.B(n_7),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_194),
.C(n_199),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_3),
.C(n_4),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_3),
.C(n_6),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_224),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_193),
.C(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_209),
.B(n_217),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_8),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_212),
.A2(n_6),
.B(n_7),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_228),
.A2(n_220),
.B(n_219),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_15),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_9),
.C(n_10),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_222),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_224),
.Y(n_237)
);

OAI31xp33_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_230),
.A3(n_233),
.B(n_228),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_241),
.B(n_9),
.Y(n_243)
);

AOI21x1_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_233),
.B(n_218),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_244),
.B(n_10),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_245),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_239),
.C(n_13),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_239),
.B(n_13),
.Y(n_248)
);


endmodule