module fake_ariane_251_n_783 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_783);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_783;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_58),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_49),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_0),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_133),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_21),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_73),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_63),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_66),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_15),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_31),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_85),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_34),
.Y(n_167)
);

BUFx4f_ASAP7_75t_SL g168 ( 
.A(n_44),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_86),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_2),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_39),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_25),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_30),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_111),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_71),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_35),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_54),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_60),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_81),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_43),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_20),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_78),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_55),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_46),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_41),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_11),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_29),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_50),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_33),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_13),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_88),
.B(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

CKINVDCx6p67_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

BUFx8_ASAP7_75t_SL g210 ( 
.A(n_175),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_1),
.Y(n_212)
);

OAI22x1_ASAP7_75t_SL g213 ( 
.A1(n_147),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_3),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_4),
.Y(n_223)
);

BUFx8_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

OA22x2_ASAP7_75t_SL g229 ( 
.A1(n_175),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

OAI22x1_ASAP7_75t_SL g231 ( 
.A1(n_181),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_151),
.B(n_8),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_185),
.A2(n_196),
.B(n_168),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_210),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_210),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_205),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_206),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_241),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_222),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_227),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_R g260 ( 
.A(n_239),
.B(n_196),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_145),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_R g263 ( 
.A(n_232),
.B(n_148),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_230),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_230),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_181),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_230),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_224),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_SL g270 ( 
.A(n_220),
.B(n_169),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_204),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_204),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_224),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_215),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_150),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_203),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_191),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_203),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_205),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_239),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_238),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_238),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_235),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_212),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_205),
.B(n_153),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_220),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_237),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_237),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_223),
.B(n_240),
.C(n_242),
.Y(n_295)
);

BUFx6f_ASAP7_75t_SL g296 ( 
.A(n_274),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_235),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_235),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_223),
.B(n_240),
.C(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_237),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_235),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_240),
.B1(n_223),
.B2(n_213),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_267),
.C(n_250),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_274),
.B(n_233),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_218),
.C(n_229),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_236),
.B(n_228),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_271),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_251),
.B(n_215),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_257),
.B(n_209),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_255),
.B(n_219),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_219),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_219),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_SL g317 ( 
.A(n_244),
.B(n_231),
.C(n_214),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_269),
.B(n_209),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_209),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_228),
.C(n_202),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_L g325 ( 
.A(n_260),
.B(n_154),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_245),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_275),
.B(n_202),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_279),
.B(n_155),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_201),
.C(n_221),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_272),
.B(n_157),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_262),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_264),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_265),
.B(n_219),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_256),
.B(n_221),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_247),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_256),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_247),
.B(n_160),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_246),
.B(n_164),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_246),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_286),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_271),
.B(n_221),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_253),
.B(n_221),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_286),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_287),
.B(n_165),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_287),
.B(n_171),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_311),
.B(n_226),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_307),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_226),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_301),
.B(n_226),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_293),
.B(n_226),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_R g364 ( 
.A(n_296),
.B(n_173),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

OR2x6_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_200),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_319),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_306),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_174),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_352),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_346),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_293),
.B(n_200),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_177),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_312),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_8),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_294),
.B(n_180),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_183),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_294),
.A2(n_207),
.B(n_194),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_348),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_309),
.A2(n_190),
.B1(n_188),
.B2(n_186),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_336),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_295),
.B(n_208),
.Y(n_390)
);

AND2x6_ASAP7_75t_SL g391 ( 
.A(n_351),
.B(n_9),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_347),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_300),
.B(n_208),
.Y(n_396)
);

BUFx12f_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_299),
.B(n_207),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_330),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_345),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_310),
.B(n_298),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_296),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_305),
.A2(n_211),
.B1(n_208),
.B2(n_207),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_344),
.B(n_207),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_208),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_308),
.A2(n_211),
.B1(n_10),
.B2(n_11),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_310),
.A2(n_211),
.B(n_10),
.C(n_12),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_339),
.B(n_9),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_328),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_313),
.B(n_211),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_333),
.B(n_357),
.Y(n_422)
);

AND3x2_ASAP7_75t_SL g423 ( 
.A(n_317),
.B(n_12),
.C(n_13),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_321),
.Y(n_424)
);

NOR2x1p5_ASAP7_75t_L g425 ( 
.A(n_341),
.B(n_14),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_342),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_349),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

AO21x1_ASAP7_75t_L g429 ( 
.A1(n_402),
.A2(n_320),
.B(n_304),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_360),
.A2(n_343),
.B(n_340),
.C(n_337),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_350),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_325),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_369),
.B(n_326),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_374),
.A2(n_321),
.B(n_326),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

AOI221xp5_ASAP7_75t_L g437 ( 
.A1(n_415),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_17),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

NOR2x1_ASAP7_75t_R g439 ( 
.A(n_403),
.B(n_17),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_368),
.A2(n_375),
.B(n_380),
.C(n_413),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_L g441 ( 
.A(n_381),
.B(n_326),
.C(n_19),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_397),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_376),
.A2(n_326),
.B1(n_22),
.B2(n_23),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_326),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_392),
.B(n_18),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_378),
.B(n_24),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_374),
.A2(n_26),
.B(n_27),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_395),
.B(n_28),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_32),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_392),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_369),
.B(n_36),
.Y(n_455)
);

AO21x1_ASAP7_75t_L g456 ( 
.A1(n_402),
.A2(n_143),
.B(n_38),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_406),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_361),
.A2(n_37),
.B(n_40),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_361),
.A2(n_42),
.B(n_45),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_383),
.B(n_47),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_408),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_384),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_53),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

O2A1O1Ixp33_ASAP7_75t_SL g466 ( 
.A1(n_409),
.A2(n_371),
.B(n_411),
.C(n_390),
.Y(n_466)
);

O2A1O1Ixp33_ASAP7_75t_L g467 ( 
.A1(n_362),
.A2(n_56),
.B(n_57),
.C(n_59),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_362),
.A2(n_61),
.B(n_62),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_388),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_389),
.B(n_64),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_379),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_363),
.A2(n_72),
.B(n_74),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

O2A1O1Ixp5_ASAP7_75t_L g474 ( 
.A1(n_382),
.A2(n_77),
.B(n_79),
.C(n_80),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_415),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_385),
.B(n_82),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_364),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_400),
.B(n_84),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_418),
.B(n_87),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_399),
.B(n_139),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

BUFx2_ASAP7_75t_SL g485 ( 
.A(n_443),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_435),
.A2(n_450),
.B(n_479),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_432),
.B(n_431),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_429),
.A2(n_390),
.B(n_396),
.Y(n_488)
);

BUFx8_ASAP7_75t_L g489 ( 
.A(n_475),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_438),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

AOI22x1_ASAP7_75t_L g493 ( 
.A1(n_451),
.A2(n_425),
.B1(n_377),
.B2(n_422),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_396),
.B(n_421),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_457),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_434),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_450),
.A2(n_363),
.B(n_421),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_470),
.A2(n_424),
.B(n_398),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_447),
.Y(n_501)
);

AO21x2_ASAP7_75t_L g502 ( 
.A1(n_470),
.A2(n_417),
.B(n_414),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_449),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_479),
.A2(n_420),
.B(n_412),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_440),
.A2(n_366),
.B(n_407),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_442),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

CKINVDCx8_ASAP7_75t_R g508 ( 
.A(n_464),
.Y(n_508)
);

AO21x2_ASAP7_75t_L g509 ( 
.A1(n_466),
.A2(n_379),
.B(n_366),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_447),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_472),
.A2(n_459),
.B(n_458),
.Y(n_511)
);

INVx8_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_448),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_482),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_482),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_465),
.B(n_410),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_468),
.A2(n_366),
.B(n_90),
.Y(n_519)
);

INVx3_ASAP7_75t_SL g520 ( 
.A(n_427),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_441),
.A2(n_423),
.B(n_91),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_469),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_446),
.B(n_391),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_433),
.B(n_89),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_463),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_456),
.A2(n_92),
.B(n_93),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_477),
.A2(n_94),
.B(n_95),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_484),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_476),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_480),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_460),
.B(n_96),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_455),
.B(n_97),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_494),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_512),
.A2(n_437),
.B1(n_462),
.B2(n_481),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_512),
.A2(n_437),
.B1(n_462),
.B2(n_483),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

BUFx4f_ASAP7_75t_L g539 ( 
.A(n_512),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_519),
.A2(n_452),
.B(n_467),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_487),
.B(n_430),
.C(n_471),
.Y(n_541)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_494),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g545 ( 
.A1(n_508),
.A2(n_444),
.B1(n_445),
.B2(n_453),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_496),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_499),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_492),
.Y(n_548)
);

AO21x1_ASAP7_75t_SL g549 ( 
.A1(n_528),
.A2(n_522),
.B(n_524),
.Y(n_549)
);

BUFx8_ASAP7_75t_SL g550 ( 
.A(n_523),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_529),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_508),
.A2(n_445),
.B1(n_478),
.B2(n_439),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_512),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_498),
.A2(n_103),
.B(n_105),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_492),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_523),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_497),
.B(n_106),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_519),
.A2(n_107),
.B(n_108),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_516),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_506),
.Y(n_561)
);

AO21x2_ASAP7_75t_L g562 ( 
.A1(n_502),
.A2(n_109),
.B(n_110),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_489),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_506),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

INVxp33_ASAP7_75t_L g566 ( 
.A(n_516),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_523),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_523),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_530),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_489),
.Y(n_570)
);

AOI21x1_ASAP7_75t_L g571 ( 
.A1(n_498),
.A2(n_123),
.B(n_124),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_520),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_514),
.B(n_126),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_520),
.Y(n_575)
);

AOI21x1_ASAP7_75t_L g576 ( 
.A1(n_495),
.A2(n_127),
.B(n_128),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_536),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_544),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_SL g579 ( 
.A(n_535),
.B(n_533),
.C(n_525),
.Y(n_579)
);

NOR2x1_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_517),
.Y(n_580)
);

AO31x2_ASAP7_75t_L g581 ( 
.A1(n_538),
.A2(n_526),
.A3(n_513),
.B(n_502),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_541),
.A2(n_521),
.B1(n_493),
.B2(n_530),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_503),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_SL g585 ( 
.A(n_570),
.B(n_521),
.C(n_485),
.Y(n_585)
);

BUFx3_ASAP7_75t_R g586 ( 
.A(n_563),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_570),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_557),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_573),
.B(n_507),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_573),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_537),
.A2(n_533),
.B(n_532),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_572),
.B(n_507),
.Y(n_592)
);

OA21x2_ASAP7_75t_L g593 ( 
.A1(n_540),
.A2(n_486),
.B(n_500),
.Y(n_593)
);

CKINVDCx8_ASAP7_75t_R g594 ( 
.A(n_575),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_550),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_SL g596 ( 
.A(n_552),
.B(n_521),
.C(n_530),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_550),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_539),
.B(n_517),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_546),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_547),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_SL g601 ( 
.A(n_567),
.B(n_511),
.C(n_527),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_566),
.B(n_501),
.Y(n_602)
);

AO31x2_ASAP7_75t_L g603 ( 
.A1(n_543),
.A2(n_526),
.A3(n_502),
.B(n_486),
.Y(n_603)
);

AO31x2_ASAP7_75t_L g604 ( 
.A1(n_543),
.A2(n_488),
.A3(n_509),
.B(n_504),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_551),
.Y(n_605)
);

AND2x4_ASAP7_75t_SL g606 ( 
.A(n_574),
.B(n_510),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_566),
.B(n_531),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_534),
.B(n_501),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_556),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_545),
.A2(n_532),
.B(n_509),
.C(n_525),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g611 ( 
.A(n_534),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_562),
.A2(n_532),
.B1(n_509),
.B2(n_505),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_510),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_558),
.B(n_510),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_SL g615 ( 
.A1(n_555),
.A2(n_515),
.B(n_514),
.C(n_518),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_561),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_565),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_574),
.B(n_518),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_548),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_548),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_549),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_555),
.Y(n_623)
);

AO32x2_ASAP7_75t_L g624 ( 
.A1(n_562),
.A2(n_488),
.A3(n_505),
.B1(n_504),
.B2(n_495),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_539),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_555),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_564),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_542),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_581),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_488),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_599),
.B(n_562),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_581),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_619),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_603),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_584),
.B(n_568),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_611),
.B(n_554),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_603),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_603),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_609),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_585),
.B(n_518),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_616),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_578),
.B(n_514),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_620),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_602),
.B(n_600),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_593),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_605),
.B(n_554),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_617),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_622),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_627),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_614),
.B(n_515),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_624),
.B(n_626),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_607),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_604),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_608),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_604),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_580),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_579),
.A2(n_518),
.B1(n_569),
.B2(n_553),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_621),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_628),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_624),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_624),
.B(n_554),
.Y(n_662)
);

INVx3_ASAP7_75t_SL g663 ( 
.A(n_595),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_596),
.B(n_559),
.Y(n_665)
);

OAI211xp5_ASAP7_75t_L g666 ( 
.A1(n_591),
.A2(n_571),
.B(n_576),
.C(n_527),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_589),
.B(n_515),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_652),
.B(n_612),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_652),
.B(n_583),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_630),
.B(n_601),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_660),
.B(n_653),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_630),
.B(n_588),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_657),
.B(n_610),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_613),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_655),
.B(n_644),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_633),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_648),
.B(n_594),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_665),
.B(n_590),
.C(n_623),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_650),
.B(n_613),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_636),
.B(n_618),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_633),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_635),
.A2(n_618),
.B1(n_592),
.B2(n_606),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_659),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_639),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_646),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_641),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_631),
.B(n_559),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_631),
.B(n_540),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_641),
.B(n_625),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_661),
.B(n_597),
.Y(n_691)
);

AOI221xp5_ASAP7_75t_L g692 ( 
.A1(n_661),
.A2(n_587),
.B1(n_586),
.B2(n_615),
.C(n_598),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_651),
.B(n_542),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_659),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_646),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_676),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_672),
.B(n_663),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_685),
.B(n_662),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_687),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_670),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_683),
.B(n_643),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_672),
.B(n_663),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_694),
.B(n_691),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_691),
.B(n_643),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_671),
.B(n_664),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_670),
.B(n_662),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_675),
.B(n_664),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_684),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_676),
.Y(n_709)
);

NAND4xp75_ASAP7_75t_SL g710 ( 
.A(n_697),
.B(n_665),
.C(n_669),
.D(n_688),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_700),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_699),
.B(n_669),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_705),
.B(n_683),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_706),
.A2(n_668),
.B1(n_673),
.B2(n_678),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_702),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_708),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_700),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_706),
.B(n_707),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_711),
.B(n_703),
.Y(n_719)
);

OAI21xp33_ASAP7_75t_L g720 ( 
.A1(n_714),
.A2(n_698),
.B(n_668),
.Y(n_720)
);

XOR2x2_ASAP7_75t_L g721 ( 
.A(n_714),
.B(n_678),
.Y(n_721)
);

OAI21xp33_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_712),
.B(n_713),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_L g723 ( 
.A(n_716),
.B(n_683),
.C(n_692),
.Y(n_723)
);

INVxp33_ASAP7_75t_L g724 ( 
.A(n_721),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_719),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_723),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_722),
.B(n_715),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_720),
.B(n_718),
.Y(n_728)
);

NAND4xp25_ASAP7_75t_SL g729 ( 
.A(n_723),
.B(n_710),
.C(n_698),
.D(n_677),
.Y(n_729)
);

AOI211xp5_ASAP7_75t_L g730 ( 
.A1(n_724),
.A2(n_666),
.B(n_690),
.C(n_688),
.Y(n_730)
);

NAND4xp25_ASAP7_75t_SL g731 ( 
.A(n_726),
.B(n_682),
.C(n_704),
.D(n_658),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_727),
.B(n_701),
.Y(n_732)
);

OA22x2_ASAP7_75t_L g733 ( 
.A1(n_732),
.A2(n_725),
.B1(n_724),
.B2(n_727),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_730),
.B(n_728),
.Y(n_734)
);

AOI221xp5_ASAP7_75t_L g735 ( 
.A1(n_734),
.A2(n_731),
.B1(n_729),
.B2(n_684),
.C(n_686),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_733),
.B(n_701),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_733),
.A2(n_642),
.B(n_690),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_735),
.A2(n_690),
.B1(n_686),
.B2(n_679),
.Y(n_738)
);

NOR2x1_ASAP7_75t_L g739 ( 
.A(n_736),
.B(n_640),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_737),
.B(n_645),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_736),
.B(n_679),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_736),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_736),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_742),
.B(n_667),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_741),
.Y(n_745)
);

XNOR2x1_ASAP7_75t_L g746 ( 
.A(n_743),
.B(n_680),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_738),
.B(n_645),
.Y(n_747)
);

NAND4xp75_ASAP7_75t_L g748 ( 
.A(n_739),
.B(n_740),
.C(n_693),
.D(n_689),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_742),
.B(n_674),
.Y(n_749)
);

CKINVDCx14_ASAP7_75t_R g750 ( 
.A(n_745),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_744),
.Y(n_751)
);

AND2x2_ASAP7_75t_SL g752 ( 
.A(n_749),
.B(n_674),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_746),
.B(n_515),
.C(n_645),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_748),
.B(n_747),
.Y(n_754)
);

XNOR2x1_ASAP7_75t_L g755 ( 
.A(n_746),
.B(n_680),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_751),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_750),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_754),
.B(n_515),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_755),
.Y(n_759)
);

NAND3xp33_ASAP7_75t_SL g760 ( 
.A(n_753),
.B(n_689),
.C(n_709),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_752),
.B(n_674),
.Y(n_761)
);

XOR2xp5_ASAP7_75t_L g762 ( 
.A(n_750),
.B(n_680),
.Y(n_762)
);

AOI22x1_ASAP7_75t_L g763 ( 
.A1(n_751),
.A2(n_709),
.B1(n_696),
.B2(n_681),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_754),
.A2(n_681),
.B1(n_542),
.B2(n_634),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_759),
.A2(n_649),
.B1(n_647),
.B2(n_634),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_757),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_762),
.A2(n_637),
.B1(n_638),
.B2(n_495),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_756),
.B(n_130),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_758),
.A2(n_637),
.B1(n_638),
.B2(n_649),
.Y(n_769)
);

OAI31xp33_ASAP7_75t_L g770 ( 
.A1(n_761),
.A2(n_632),
.A3(n_629),
.B(n_656),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_764),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_763),
.A2(n_656),
.B1(n_654),
.B2(n_632),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_768),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_766),
.Y(n_774)
);

XNOR2xp5_ASAP7_75t_L g775 ( 
.A(n_771),
.B(n_760),
.Y(n_775)
);

AOI21xp33_ASAP7_75t_SL g776 ( 
.A1(n_767),
.A2(n_131),
.B(n_132),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_769),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_774),
.B(n_765),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_773),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_778),
.A2(n_775),
.B(n_776),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_SL g781 ( 
.A1(n_780),
.A2(n_779),
.B1(n_777),
.B2(n_772),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_781),
.B(n_770),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_782),
.A2(n_500),
.B1(n_647),
.B2(n_511),
.Y(n_783)
);


endmodule