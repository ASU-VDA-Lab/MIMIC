module fake_netlist_6_1366_n_726 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_726);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_726;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_41),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_4),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_19),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_49),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_4),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_0),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_58),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_18),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_28),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_94),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_64),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_54),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_50),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_11),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_19),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_59),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_24),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_61),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_68),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_53),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_79),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_26),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_82),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_29),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_46),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_124),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

BUFx8_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_22),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_1),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_2),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_3),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_5),
.Y(n_219)
);

CKINVDCx8_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_145),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_23),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_7),
.B(n_8),
.Y(n_224)
);

AOI22x1_ASAP7_75t_L g225 ( 
.A1(n_146),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_144),
.B(n_10),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_156),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_147),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_165),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

BUFx8_ASAP7_75t_SL g236 ( 
.A(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_166),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_187),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_148),
.C(n_194),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_220),
.B(n_153),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_169),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_155),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_174),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_179),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_180),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_183),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

CKINVDCx8_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_212),
.A2(n_195),
.B1(n_193),
.B2(n_192),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_204),
.B(n_158),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_186),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_204),
.B(n_159),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_236),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_227),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_209),
.B(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_191),
.B1(n_188),
.B2(n_190),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_214),
.B(n_167),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_222),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_224),
.B(n_201),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_218),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_219),
.B1(n_225),
.B2(n_237),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_218),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_200),
.B(n_197),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_232),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_252),
.B(n_222),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_247),
.B(n_218),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_211),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_277),
.B(n_211),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_242),
.B(n_252),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_218),
.Y(n_306)
);

NAND2x1p5_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_224),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_211),
.Y(n_308)
);

AND2x6_ASAP7_75t_SL g309 ( 
.A(n_238),
.B(n_199),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_196),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_222),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_210),
.Y(n_313)
);

BUFx6f_ASAP7_75t_SL g314 ( 
.A(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_230),
.B1(n_229),
.B2(n_214),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_263),
.B(n_232),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_196),
.Y(n_319)
);

AO221x1_ASAP7_75t_L g320 ( 
.A1(n_248),
.A2(n_230),
.B1(n_211),
.B2(n_229),
.C(n_216),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_252),
.B(n_198),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_243),
.B(n_168),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_258),
.A2(n_217),
.B(n_201),
.C(n_202),
.Y(n_323)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_234),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_245),
.B(n_205),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_259),
.A2(n_221),
.B1(n_171),
.B2(n_170),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_260),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_261),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_260),
.B(n_267),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_261),
.B(n_229),
.C(n_182),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_254),
.B(n_236),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_267),
.B(n_223),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_268),
.B(n_185),
.C(n_198),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_253),
.B(n_198),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_249),
.B(n_202),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_285),
.A2(n_253),
.B(n_280),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_293),
.A2(n_280),
.B(n_282),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_296),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_250),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_326),
.A2(n_268),
.B1(n_215),
.B2(n_223),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_287),
.A2(n_248),
.B(n_256),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_217),
.B1(n_215),
.B2(n_250),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_311),
.Y(n_349)
);

AOI21x1_ASAP7_75t_L g350 ( 
.A1(n_289),
.A2(n_81),
.B(n_142),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_302),
.A2(n_80),
.B1(n_139),
.B2(n_138),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_289),
.A2(n_75),
.B(n_137),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_25),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_290),
.B(n_13),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_27),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_30),
.Y(n_356)
);

AO22x1_ASAP7_75t_L g357 ( 
.A1(n_333),
.A2(n_321),
.B1(n_318),
.B2(n_330),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_313),
.A2(n_83),
.B1(n_136),
.B2(n_135),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_324),
.A2(n_76),
.B(n_132),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_323),
.A2(n_74),
.B(n_131),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_291),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_14),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_295),
.B(n_31),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g365 ( 
.A(n_322),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_309),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_R g368 ( 
.A(n_314),
.B(n_32),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_286),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_33),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_324),
.A2(n_86),
.B(n_129),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_15),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_324),
.A2(n_73),
.B(n_128),
.Y(n_373)
);

O2A1O1Ixp5_ASAP7_75t_L g374 ( 
.A1(n_299),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_16),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_286),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_312),
.A2(n_88),
.B(n_126),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_310),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_288),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_300),
.B(n_303),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_334),
.A2(n_90),
.B(n_125),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_334),
.A2(n_72),
.B(n_122),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_319),
.A2(n_71),
.B(n_121),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_292),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_294),
.A2(n_69),
.B1(n_120),
.B2(n_34),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_294),
.A2(n_67),
.B1(n_119),
.B2(n_35),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_305),
.A2(n_304),
.B(n_306),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_307),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_306),
.A2(n_91),
.B(n_118),
.Y(n_390)
);

NOR2x1_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_65),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_335),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_315),
.A2(n_62),
.B1(n_116),
.B2(n_36),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_336),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_301),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_317),
.B(n_92),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_339),
.A2(n_60),
.B(n_115),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_343),
.B(n_317),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_320),
.Y(n_399)
);

OAI22x1_ASAP7_75t_L g400 ( 
.A1(n_372),
.A2(n_314),
.B1(n_21),
.B2(n_20),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_363),
.B1(n_366),
.B2(n_381),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_317),
.Y(n_402)
);

AO31x2_ASAP7_75t_L g403 ( 
.A1(n_363),
.A2(n_317),
.A3(n_21),
.B(n_297),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_297),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

AO22x2_ASAP7_75t_L g406 ( 
.A1(n_375),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_40),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_344),
.A2(n_340),
.B(n_369),
.Y(n_409)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_361),
.A2(n_42),
.B(n_43),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_369),
.A2(n_44),
.B(n_45),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_392),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_348),
.B(n_388),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

OAI21xp33_ASAP7_75t_L g415 ( 
.A1(n_379),
.A2(n_47),
.B(n_48),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_347),
.A2(n_51),
.B(n_52),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_353),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_93),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_362),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_95),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_97),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_98),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_365),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_350),
.Y(n_425)
);

NAND2x1_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_99),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_100),
.Y(n_427)
);

AO31x2_ASAP7_75t_L g428 ( 
.A1(n_356),
.A2(n_364),
.A3(n_396),
.B(n_377),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_359),
.B(n_101),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_104),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_105),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_385),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_345),
.B(n_106),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_357),
.B(n_109),
.Y(n_434)
);

AOI21x1_ASAP7_75t_L g435 ( 
.A1(n_342),
.A2(n_111),
.B(n_113),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_368),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_351),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_393),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_360),
.A2(n_373),
.B(n_371),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_374),
.A2(n_397),
.B(n_384),
.Y(n_442)
);

O2A1O1Ixp5_ASAP7_75t_L g443 ( 
.A1(n_374),
.A2(n_382),
.B(n_383),
.C(n_352),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_386),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_390),
.A2(n_387),
.B(n_358),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_369),
.A2(n_376),
.B(n_344),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

AO21x2_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_442),
.B(n_413),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_447),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_436),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_421),
.B(n_412),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_L g453 ( 
.A1(n_401),
.A2(n_415),
.B(n_427),
.C(n_446),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_420),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_404),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_399),
.B(n_415),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_406),
.A2(n_440),
.B1(n_444),
.B2(n_439),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_405),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g460 ( 
.A(n_405),
.B(n_421),
.Y(n_460)
);

CKINVDCx6p67_ASAP7_75t_R g461 ( 
.A(n_424),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_409),
.A2(n_443),
.B(n_419),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_410),
.B(n_398),
.Y(n_463)
);

NOR2x1_ASAP7_75t_SL g464 ( 
.A(n_417),
.B(n_437),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

BUFx4f_ASAP7_75t_SL g466 ( 
.A(n_424),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_423),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_405),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_422),
.A2(n_431),
.B(n_441),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_406),
.B(n_430),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_433),
.A2(n_411),
.B(n_407),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_434),
.B1(n_417),
.B2(n_400),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_418),
.B(n_417),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_403),
.B(n_416),
.Y(n_475)
);

AOI22x1_ASAP7_75t_L g476 ( 
.A1(n_425),
.A2(n_428),
.B1(n_403),
.B2(n_416),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_429),
.A2(n_425),
.B1(n_435),
.B2(n_403),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_428),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

AOI222xp33_ASAP7_75t_SL g480 ( 
.A1(n_414),
.A2(n_172),
.B1(n_200),
.B2(n_149),
.C1(n_189),
.C2(n_178),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_438),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_412),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_421),
.B(n_447),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_440),
.A2(n_401),
.B1(n_447),
.B2(n_275),
.Y(n_486)
);

OAI21x1_ASAP7_75t_SL g487 ( 
.A1(n_410),
.A2(n_407),
.B(n_411),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_447),
.B(n_412),
.Y(n_488)
);

O2A1O1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_415),
.A2(n_379),
.B(n_354),
.C(n_275),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_SL g491 ( 
.A1(n_458),
.A2(n_471),
.B1(n_480),
.B2(n_448),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_462),
.A2(n_477),
.B(n_453),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_478),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_450),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_479),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_459),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_448),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_476),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_457),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_467),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_474),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_472),
.B(n_475),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_483),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_451),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_454),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_459),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_471),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_460),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_484),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_462),
.A2(n_472),
.B(n_477),
.Y(n_514)
);

NAND2x1_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_487),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_463),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_456),
.A2(n_458),
.B(n_489),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_471),
.A2(n_449),
.B1(n_473),
.B2(n_474),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_456),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_465),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_464),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_459),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_469),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_496),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_496),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_525),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_493),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_481),
.Y(n_532)
);

AOI221x1_ASAP7_75t_SL g533 ( 
.A1(n_490),
.A2(n_480),
.B1(n_494),
.B2(n_512),
.C(n_517),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_497),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_502),
.B(n_459),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_461),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_524),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_502),
.B(n_468),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_503),
.B(n_468),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_497),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_526),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_470),
.Y(n_543)
);

NOR2x1_ASAP7_75t_SL g544 ( 
.A(n_504),
.B(n_469),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_490),
.B(n_466),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_526),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_526),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_494),
.B(n_521),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_521),
.B(n_507),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_525),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_524),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_504),
.B(n_510),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_495),
.B(n_491),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_518),
.B(n_495),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_500),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_491),
.B(n_522),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_507),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_498),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_522),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_520),
.B(n_498),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_504),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_504),
.B(n_510),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_500),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_504),
.B(n_523),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_504),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_518),
.B(n_505),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_522),
.B(n_513),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_512),
.B(n_513),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_505),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_517),
.B(n_511),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_504),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_551),
.B(n_492),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_555),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_492),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_508),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_568),
.B(n_492),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_568),
.B(n_492),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_501),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_553),
.B(n_514),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_549),
.B(n_508),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_566),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_519),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_538),
.B(n_519),
.Y(n_586)
);

NAND2x1p5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_566),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_555),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_560),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_553),
.B(n_557),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_539),
.B(n_523),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_556),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_570),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_539),
.B(n_542),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_532),
.B(n_509),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_572),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_557),
.B(n_514),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_545),
.B(n_529),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_535),
.B(n_514),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_528),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_565),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_533),
.B(n_509),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_535),
.B(n_514),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_536),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_527),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_537),
.B(n_514),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_537),
.B(n_516),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_529),
.Y(n_610)
);

NOR2x1_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_536),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_598),
.B(n_564),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_596),
.B(n_528),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_578),
.B(n_571),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_575),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_605),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_595),
.B(n_564),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_575),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_599),
.B(n_554),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_580),
.B(n_563),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_580),
.B(n_563),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_588),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_588),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_599),
.B(n_554),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_604),
.B(n_571),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_583),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_592),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_604),
.B(n_597),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_580),
.B(n_566),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_592),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_601),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_594),
.B(n_548),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_597),
.B(n_574),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_574),
.B(n_541),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_576),
.B(n_541),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_601),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_607),
.B(n_543),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_602),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_602),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_600),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_578),
.B(n_546),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_576),
.B(n_547),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_614),
.B(n_579),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_633),
.B(n_581),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_629),
.B(n_580),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_619),
.B(n_581),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_619),
.B(n_605),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_622),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_616),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_614),
.B(n_579),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_615),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_624),
.B(n_606),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_622),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_623),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_628),
.B(n_608),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_628),
.B(n_608),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_611),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_615),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_627),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_643),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_648),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_657),
.A2(n_589),
.B(n_617),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_653),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_647),
.A2(n_562),
.B1(n_591),
.B2(n_603),
.Y(n_664)
);

OAI221xp5_ASAP7_75t_L g665 ( 
.A1(n_649),
.A2(n_613),
.B1(n_640),
.B2(n_632),
.C(n_637),
.Y(n_665)
);

OAI211xp5_ASAP7_75t_SL g666 ( 
.A1(n_647),
.A2(n_612),
.B(n_586),
.C(n_584),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_644),
.B(n_633),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_654),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_650),
.B(n_625),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_652),
.B(n_646),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_658),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_661),
.Y(n_672)
);

AOI22x1_ASAP7_75t_L g673 ( 
.A1(n_662),
.A2(n_645),
.B1(n_621),
.B2(n_620),
.Y(n_673)
);

OAI322xp33_ASAP7_75t_L g674 ( 
.A1(n_664),
.A2(n_652),
.A3(n_658),
.B1(n_646),
.B2(n_656),
.C1(n_655),
.C2(n_577),
.Y(n_674)
);

AOI211x1_ASAP7_75t_L g675 ( 
.A1(n_665),
.A2(n_590),
.B(n_624),
.C(n_625),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_663),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_670),
.B(n_651),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_671),
.B(n_659),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_667),
.B(n_645),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_SL g680 ( 
.A(n_678),
.B(n_660),
.C(n_668),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_673),
.B(n_666),
.C(n_618),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_674),
.B(n_679),
.Y(n_682)
);

NAND2xp67_ASAP7_75t_SL g683 ( 
.A(n_675),
.B(n_570),
.Y(n_683)
);

OAI211xp5_ASAP7_75t_L g684 ( 
.A1(n_672),
.A2(n_660),
.B(n_590),
.C(n_529),
.Y(n_684)
);

NOR4xp75_ASAP7_75t_L g685 ( 
.A(n_678),
.B(n_626),
.C(n_582),
.D(n_583),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_SL g686 ( 
.A1(n_682),
.A2(n_629),
.B(n_620),
.Y(n_686)
);

NAND4xp25_ASAP7_75t_L g687 ( 
.A(n_681),
.B(n_550),
.C(n_677),
.D(n_676),
.Y(n_687)
);

NAND5xp2_ASAP7_75t_L g688 ( 
.A(n_684),
.B(n_587),
.C(n_543),
.D(n_561),
.E(n_593),
.Y(n_688)
);

NOR3x1_ASAP7_75t_L g689 ( 
.A(n_680),
.B(n_669),
.C(n_585),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_683),
.B(n_629),
.Y(n_690)
);

NAND4xp25_ASAP7_75t_L g691 ( 
.A(n_689),
.B(n_550),
.C(n_621),
.D(n_620),
.Y(n_691)
);

NAND5xp2_ASAP7_75t_L g692 ( 
.A(n_686),
.B(n_587),
.C(n_685),
.D(n_630),
.E(n_585),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_687),
.B(n_550),
.C(n_610),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_693),
.B(n_690),
.Y(n_694)
);

AND3x2_ASAP7_75t_L g695 ( 
.A(n_692),
.B(n_688),
.C(n_559),
.Y(n_695)
);

NAND4xp75_ASAP7_75t_L g696 ( 
.A(n_691),
.B(n_499),
.C(n_639),
.D(n_638),
.Y(n_696)
);

NAND4xp75_ASAP7_75t_L g697 ( 
.A(n_691),
.B(n_499),
.C(n_639),
.D(n_638),
.Y(n_697)
);

XNOR2x1_ASAP7_75t_L g698 ( 
.A(n_695),
.B(n_621),
.Y(n_698)
);

XNOR2xp5_ASAP7_75t_L g699 ( 
.A(n_694),
.B(n_587),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_610),
.B1(n_626),
.B2(n_583),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_697),
.Y(n_701)
);

NAND4xp75_ASAP7_75t_L g702 ( 
.A(n_694),
.B(n_499),
.C(n_636),
.D(n_631),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_698),
.A2(n_626),
.B1(n_636),
.B2(n_623),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_R g704 ( 
.A1(n_699),
.A2(n_573),
.B1(n_552),
.B2(n_564),
.C(n_631),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_702),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_701),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_700),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_701),
.B(n_627),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_706),
.A2(n_566),
.B1(n_564),
.B2(n_552),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_708),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_707),
.A2(n_641),
.B1(n_573),
.B2(n_552),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_705),
.A2(n_515),
.B(n_573),
.Y(n_712)
);

XNOR2xp5_ASAP7_75t_L g713 ( 
.A(n_703),
.B(n_515),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_710),
.Y(n_714)
);

OAI22x1_ASAP7_75t_L g715 ( 
.A1(n_709),
.A2(n_704),
.B1(n_606),
.B2(n_569),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_712),
.A2(n_509),
.B1(n_501),
.B2(n_569),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_713),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_711),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_717),
.A2(n_642),
.B1(n_634),
.B2(n_635),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_718),
.A2(n_642),
.B1(n_634),
.B2(n_635),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_714),
.A2(n_609),
.B1(n_540),
.B2(n_531),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_SL g722 ( 
.A1(n_720),
.A2(n_716),
.B1(n_715),
.B2(n_719),
.Y(n_722)
);

AOI222xp33_ASAP7_75t_L g723 ( 
.A1(n_721),
.A2(n_716),
.B1(n_544),
.B2(n_501),
.C1(n_540),
.C2(n_534),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_723),
.B(n_531),
.C(n_534),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_724),
.B(n_722),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_SL g726 ( 
.A1(n_725),
.A2(n_544),
.B1(n_530),
.B2(n_609),
.Y(n_726)
);


endmodule