module fake_jpeg_4330_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_26),
.B1(n_22),
.B2(n_31),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_35),
.A2(n_26),
.B1(n_22),
.B2(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_8),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_18),
.Y(n_85)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_22),
.B1(n_31),
.B2(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_20),
.B1(n_38),
.B2(n_25),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_27),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_28),
.B(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_66),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_61),
.Y(n_75)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_26),
.B1(n_31),
.B2(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_77),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_34),
.B1(n_40),
.B2(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_71),
.B1(n_20),
.B2(n_45),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_34),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_19),
.B(n_23),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_28),
.B(n_30),
.C(n_25),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_20),
.B1(n_30),
.B2(n_34),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_20),
.B1(n_30),
.B2(n_38),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_90),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_33),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_34),
.C(n_38),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_23),
.C(n_18),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_52),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_63),
.B1(n_62),
.B2(n_57),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_66),
.B1(n_58),
.B2(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_106),
.B1(n_118),
.B2(n_70),
.Y(n_125)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_70),
.B(n_19),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_77),
.B(n_25),
.Y(n_144)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_60),
.B1(n_47),
.B2(n_56),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_78),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_81),
.B1(n_94),
.B2(n_80),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_40),
.C(n_37),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_122),
.C(n_70),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_137),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_76),
.B1(n_70),
.B2(n_88),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_105),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_136),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_143),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_74),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_139),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_90),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_148),
.B(n_152),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_95),
.B1(n_87),
.B2(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_141),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_80),
.C(n_91),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_97),
.B(n_112),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_111),
.B(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_129),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_72),
.C(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_65),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_75),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_96),
.A2(n_83),
.B1(n_72),
.B2(n_75),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_151),
.B1(n_119),
.B2(n_108),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_83),
.B1(n_75),
.B2(n_93),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_32),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_166),
.B(n_153),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_111),
.B(n_103),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_166),
.B(n_183),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_159),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_114),
.C(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_165),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_114),
.B1(n_104),
.B2(n_37),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_129),
.B1(n_141),
.B2(n_131),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_133),
.C(n_146),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_101),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_138),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_98),
.B1(n_101),
.B2(n_108),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_182),
.B1(n_24),
.B2(n_21),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_130),
.B1(n_124),
.B2(n_119),
.Y(n_203)
);

AO22x1_ASAP7_75t_SL g182 ( 
.A1(n_125),
.A2(n_52),
.B1(n_17),
.B2(n_21),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_128),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_200),
.C(n_40),
.Y(n_230)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_179),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_201),
.Y(n_215)
);

OAI22x1_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_144),
.B1(n_132),
.B2(n_135),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_135),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_173),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_153),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_126),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_155),
.CI(n_159),
.CON(n_223),
.SN(n_223)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_152),
.B1(n_93),
.B2(n_52),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_33),
.B1(n_32),
.B2(n_43),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_40),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_178),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_167),
.A2(n_33),
.B1(n_32),
.B2(n_43),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_226),
.B1(n_206),
.B2(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_163),
.B(n_170),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_221),
.B(n_234),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_163),
.B1(n_171),
.B2(n_182),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_196),
.B1(n_197),
.B2(n_210),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_158),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_232),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_190),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_208),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_191),
.A2(n_160),
.B1(n_162),
.B2(n_164),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_157),
.A3(n_183),
.B1(n_169),
.B2(n_43),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_231),
.C(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_65),
.C(n_49),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_73),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_65),
.C(n_49),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_189),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_246),
.C(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_230),
.C(n_195),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_245),
.C(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_195),
.C(n_201),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_0),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_202),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_185),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_229),
.C(n_211),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_193),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_254),
.B1(n_227),
.B2(n_235),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_204),
.B1(n_196),
.B2(n_24),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_49),
.C(n_73),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_234),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_258),
.B(n_259),
.Y(n_273)
);

FAx1_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_218),
.CI(n_223),
.CON(n_258),
.SN(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_219),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_219),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_261),
.B(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_212),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_212),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_214),
.C(n_223),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_227),
.C(n_228),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_236),
.B(n_242),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_21),
.C(n_17),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_244),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_277),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_280),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_276),
.B(n_0),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_253),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_280),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_251),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_245),
.B1(n_255),
.B2(n_240),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_0),
.Y(n_289)
);

FAx1_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_17),
.CI(n_21),
.CON(n_283),
.SN(n_283)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_264),
.B(n_11),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_264),
.B1(n_17),
.B2(n_24),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_287),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_294),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_291),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_10),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_279),
.B1(n_281),
.B2(n_274),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_286),
.Y(n_304)
);

AOI31xp67_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_7),
.A3(n_15),
.B(n_14),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_302),
.C(n_11),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_7),
.C(n_15),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_13),
.B(n_3),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_16),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_304),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_16),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.C1(n_5),
.C2(n_1),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_16),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_310),
.B1(n_302),
.B2(n_300),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_2),
.Y(n_310)
);

AOI321xp33_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_312),
.A3(n_305),
.B1(n_298),
.B2(n_311),
.C(n_2),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_303),
.C2(n_297),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_315),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_3),
.Y(n_317)
);


endmodule