module real_jpeg_5364_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_0),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_0),
.B(n_52),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_0),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_0),
.B(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_2),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_2),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_2),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_2),
.B(n_26),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_2),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_52),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_3),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_3),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_3),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_3),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_3),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_3),
.B(n_239),
.Y(n_447)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_4),
.Y(n_299)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_6),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_6),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_6),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_6),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_6),
.B(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_7),
.Y(n_229)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_7),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_7),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_7),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_7),
.Y(n_419)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_8),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g421 ( 
.A(n_8),
.Y(n_421)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_10),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_11),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_11),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_11),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_11),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_11),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_11),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_11),
.B(n_361),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_11),
.A2(n_416),
.B(n_421),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_12),
.Y(n_149)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_12),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_13),
.B(n_153),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_13),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_13),
.B(n_270),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_13),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_13),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_13),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_14),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_14),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_14),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_14),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_14),
.B(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_14),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_15),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_15),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_15),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_15),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_15),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_15),
.B(n_330),
.Y(n_446)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_101),
.B(n_117),
.C(n_501),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_33),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_19),
.B(n_92),
.CI(n_93),
.CON(n_91),
.SN(n_91)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_25),
.C(n_28),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_20),
.A2(n_21),
.B1(n_28),
.B2(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_20),
.A2(n_21),
.B1(n_96),
.B2(n_99),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g501 ( 
.A(n_20),
.B(n_43),
.C(n_96),
.Y(n_501)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_21),
.B(n_177),
.C(n_180),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_21),
.B(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g361 ( 
.A(n_23),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_24),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_25),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_25),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_25),
.A2(n_82),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_25),
.B(n_131),
.C(n_135),
.Y(n_159)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_28),
.A2(n_38),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_28),
.B(n_224),
.C(n_230),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_28),
.A2(n_70),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_30),
.Y(n_372)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_32),
.Y(n_130)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_32),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_32),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_91),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_77),
.C(n_78),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_35),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_56),
.C(n_67),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_36),
.B(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_49),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_51),
.C(n_54),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_43),
.C(n_46),
.Y(n_37)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_70),
.C(n_76),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_38),
.A2(n_71),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_38),
.A2(n_71),
.B1(n_402),
.B2(n_406),
.Y(n_401)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_41),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_41),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_41),
.Y(n_338)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_42),
.Y(n_134)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_42),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_42),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_43),
.A2(n_94),
.B1(n_95),
.B2(n_100),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_43),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_100),
.Y(n_163)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_46),
.A2(n_47),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_46),
.B(n_111),
.C(n_118),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_46),
.A2(n_47),
.B1(n_369),
.B2(n_373),
.Y(n_368)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_47),
.B(n_369),
.C(n_374),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_56),
.B(n_67),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.C(n_63),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_57),
.Y(n_139)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_59),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_60),
.A2(n_61),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_61),
.B(n_144),
.C(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_65),
.B(n_283),
.Y(n_415)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_76),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_71),
.B(n_395),
.C(n_406),
.Y(n_441)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_118),
.C(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_72),
.A2(n_76),
.B1(n_120),
.B2(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_77),
.B(n_78),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_90),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_87),
.C(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_91),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_96),
.B(n_188),
.C(n_192),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_96),
.A2(n_99),
.B1(n_152),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_96),
.A2(n_99),
.B1(n_192),
.B2(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_142),
.C(n_152),
.Y(n_141)
);

AO21x1_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_496),
.B(n_500),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_245),
.B(n_493),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_200),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_SL g493 ( 
.A1(n_104),
.A2(n_494),
.B(n_495),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_166),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_105),
.B(n_166),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_157),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_106),
.B(n_158),
.C(n_164),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_137),
.C(n_140),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_107),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_119),
.C(n_124),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_108),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_112),
.A2(n_118),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_112),
.A2(n_118),
.B1(n_224),
.B2(n_225),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_112),
.B(n_225),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_116),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_116),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_119),
.B(n_124),
.Y(n_205)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_129),
.Y(n_264)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_130),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_131),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_131),
.B(n_214),
.Y(n_440)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_136),
.B(n_213),
.C(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_143),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_150),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_150),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_144),
.A2(n_183),
.B1(n_189),
.B2(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_144),
.A2(n_183),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_144),
.B(n_279),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_146),
.A2(n_185),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_146),
.B(n_425),
.C(n_428),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_148),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_156),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_167),
.C(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_158),
.B(n_167),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.CI(n_161),
.CON(n_158),
.SN(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_170),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_187),
.C(n_196),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_181),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_172),
.B(n_176),
.Y(n_464)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_180),
.Y(n_221)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_181),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_196),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_189),
.A2(n_211),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_189),
.B(n_381),
.Y(n_409)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_243),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_201),
.B(n_243),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.C(n_206),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_202),
.B(n_204),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_206),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_222),
.C(n_240),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_207),
.B(n_466),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_220),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_208),
.B(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_212),
.B(n_220),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_215),
.B(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_222),
.B(n_240),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.C(n_235),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_223),
.B(n_449),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_224),
.A2(n_225),
.B1(n_230),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_229),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_230),
.Y(n_458)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_231),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_232),
.A2(n_235),
.B1(n_236),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_232),
.Y(n_450)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI221xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_433),
.B1(n_486),
.B2(n_491),
.C(n_492),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_388),
.B(n_432),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_349),
.B(n_387),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_324),
.B(n_348),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_291),
.B(n_323),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_280),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_251),
.B(n_280),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_265),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_252),
.B(n_266),
.C(n_277),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_258),
.C(n_262),
.Y(n_334)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_277),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_268),
.B(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.C(n_287),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_287),
.B1(n_288),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_317),
.B(n_322),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_307),
.B(n_316),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_304),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_304),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_300),
.Y(n_318)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_312),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_326),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_333),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_334),
.C(n_335),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_331),
.C(n_332),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_340),
.C(n_347),
.Y(n_383)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_343),
.B2(n_347),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_386),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_386),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_366),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_355),
.C(n_366),
.Y(n_389)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_355)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_360),
.B2(n_362),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_357),
.B(n_362),
.C(n_363),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_360),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_379),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_383),
.C(n_385),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_374),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_369),
.Y(n_373)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_379)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_380),
.Y(n_385)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_383),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_389),
.B(n_390),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_412),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_392),
.B(n_393),
.C(n_412),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_407),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_394),
.B(n_408),
.C(n_411),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_401),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_402),
.Y(n_406)
);

INVx6_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_431),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_422),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_414),
.B(n_422),
.C(n_431),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_416),
.B(n_420),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_446),
.C(n_447),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_460),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_428),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NOR3xp33_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_468),
.C(n_472),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_434),
.A2(n_487),
.B(n_490),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_461),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_435),
.B(n_461),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_451),
.C(n_453),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_451),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_444),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_445),
.C(n_448),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_441),
.C(n_442),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_443),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_448),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_447),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_481),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.C(n_459),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_459),
.Y(n_476)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_467),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_465),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_465),
.C(n_467),
.Y(n_471)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_471),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_482),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_473),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_480),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_480),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_477),
.C(n_478),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_478),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_484),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_498),
.Y(n_500)
);


endmodule