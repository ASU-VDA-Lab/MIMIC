module fake_jpeg_2255_n_267 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_44),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_58),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_64),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_3),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_88),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_36),
.C(n_33),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_6),
.C(n_8),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_104),
.B1(n_57),
.B2(n_16),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_29),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_35),
.B1(n_32),
.B2(n_38),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_110),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_35),
.B1(n_24),
.B2(n_38),
.Y(n_93)
);

CKINVDCx9p33_ASAP7_75t_R g94 ( 
.A(n_39),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_94),
.Y(n_120)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_95),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_42),
.B1(n_35),
.B2(n_49),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_20),
.C(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_103),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_20),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_62),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_54),
.B(n_34),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_111),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_44),
.B(n_27),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_55),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_40),
.B(n_26),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_65),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_113),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_128),
.B1(n_74),
.B2(n_69),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_127),
.Y(n_148)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_17),
.B1(n_37),
.B2(n_16),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_95),
.B1(n_77),
.B2(n_69),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_76),
.A2(n_85),
.B(n_75),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_4),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_93),
.A2(n_37),
.B1(n_6),
.B2(n_8),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_5),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_9),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_9),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_136),
.B(n_133),
.Y(n_162)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_141),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_142),
.B1(n_11),
.B2(n_99),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_11),
.B1(n_12),
.B2(n_71),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_79),
.B1(n_78),
.B2(n_71),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_153),
.B1(n_157),
.B2(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_146),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_94),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_155),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_120),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_80),
.B1(n_96),
.B2(n_68),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_86),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_77),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_80),
.B1(n_96),
.B2(n_68),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_135),
.B1(n_117),
.B2(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_83),
.B1(n_90),
.B2(n_102),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_122),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_90),
.B1(n_83),
.B2(n_102),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_165),
.B1(n_143),
.B2(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_74),
.B1(n_89),
.B2(n_99),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_117),
.B1(n_135),
.B2(n_123),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_124),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_126),
.C(n_140),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_99),
.C(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_89),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_89),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_120),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_164),
.B(n_169),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_144),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_188),
.B1(n_147),
.B2(n_157),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_186),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_148),
.A2(n_113),
.B(n_116),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_192),
.B(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_129),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_181),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_176),
.A2(n_166),
.B1(n_155),
.B2(n_165),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_172),
.B1(n_176),
.B2(n_188),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_197),
.B(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_207),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_159),
.C(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_209),
.C(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_146),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_170),
.B(n_163),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_178),
.B(n_185),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_170),
.C(n_160),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_223),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_222),
.B(n_224),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_177),
.B(n_179),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_214),
.A2(n_217),
.B(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_177),
.B(n_187),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_192),
.B1(n_200),
.B2(n_195),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_202),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_174),
.A3(n_190),
.B1(n_186),
.B2(n_173),
.C1(n_181),
.C2(n_180),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_180),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_182),
.B(n_173),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_231),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_212),
.B(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_225),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_241),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_234),
.A2(n_225),
.B(n_217),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_239),
.B(n_244),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_229),
.B(n_213),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_218),
.B(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_223),
.C(n_199),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_228),
.C(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_216),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_248),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_235),
.B(n_224),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_236),
.C(n_241),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_194),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_244),
.B1(n_204),
.B2(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_260),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_201),
.B(n_210),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_210),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_175),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_180),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_253),
.A3(n_255),
.B1(n_201),
.B2(n_254),
.C1(n_191),
.C2(n_183),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_265),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_263),
.Y(n_267)
);


endmodule