module fake_jpeg_3568_n_38 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_0),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_20),
.A2(n_18),
.B(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_13),
.C(n_17),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_15),
.B1(n_17),
.B2(n_3),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_15),
.B(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_0),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_11),
.C(n_1),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_30),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_33),
.B(n_8),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_32),
.C(n_9),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_9),
.CI(n_10),
.CON(n_38),
.SN(n_38)
);


endmodule