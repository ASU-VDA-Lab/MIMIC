module fake_jpeg_26519_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_59),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_1),
.CON(n_59),
.SN(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_49),
.B1(n_43),
.B2(n_51),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_69),
.B1(n_71),
.B2(n_50),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_25),
.B(n_36),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_47),
.B1(n_46),
.B2(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_45),
.B1(n_38),
.B2(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_18),
.B1(n_31),
.B2(n_5),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_86),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_74),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_76),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_66),
.B(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_68),
.C(n_72),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_92),
.B1(n_90),
.B2(n_3),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

AOI321xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_20),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_28),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_32),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_27),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_29),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_13),
.B(n_14),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_16),
.Y(n_102)
);


endmodule