module fake_jpeg_21739_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_20),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_26),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_63),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_75),
.B1(n_53),
.B2(n_57),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_87),
.B1(n_92),
.B2(n_51),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_62),
.B1(n_76),
.B2(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_84),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_77),
.B1(n_55),
.B2(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_52),
.B1(n_69),
.B2(n_71),
.Y(n_102)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_98),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_107),
.Y(n_116)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_105),
.B1(n_108),
.B2(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_52),
.B1(n_48),
.B2(n_74),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_55),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_69),
.B1(n_50),
.B2(n_68),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_59),
.A3(n_66),
.B1(n_61),
.B2(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_0),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_118),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_0),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_123),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_63),
.B(n_2),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_1),
.B(n_2),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_1),
.B(n_3),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_65),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_130),
.B1(n_134),
.B2(n_110),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_135),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_64),
.B1(n_70),
.B2(n_14),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_64),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_11),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_146),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_110),
.C(n_15),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_142),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_136),
.B(n_128),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_148),
.A2(n_149),
.B1(n_138),
.B2(n_147),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_142),
.C(n_139),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_145),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_141),
.B(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_19),
.Y(n_159)
);

OAI321xp33_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_22),
.A3(n_24),
.B1(n_25),
.B2(n_31),
.C(n_37),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_40),
.Y(n_161)
);


endmodule