module fake_netlist_6_4763_n_2983 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_628, n_557, n_349, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2983);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2983;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2981;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_2127;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2904;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2978;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_863;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_2952;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_2968;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_2899;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_540),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_167),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_604),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_340),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_200),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_586),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_269),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_583),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_602),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_508),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_601),
.Y(n_640)
);

INVx4_ASAP7_75t_R g641 ( 
.A(n_511),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_620),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_373),
.Y(n_643)
);

BUFx5_ASAP7_75t_L g644 ( 
.A(n_75),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_441),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_214),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_448),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_603),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_327),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_501),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_77),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_592),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_596),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_376),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_584),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_94),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_384),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_299),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_471),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_495),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_591),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_451),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_541),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_589),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_431),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_78),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_178),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_58),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_239),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_348),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_489),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_504),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_235),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_499),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_599),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_244),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_540),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_193),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_317),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_131),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_473),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_305),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_458),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_34),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_504),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_625),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_502),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_95),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_503),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_605),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_224),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_21),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_217),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_336),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_308),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_99),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_588),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_291),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_361),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_61),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_322),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_250),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_135),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_414),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_611),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_598),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_124),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_210),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_593),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_83),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_564),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_82),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_402),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_509),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_290),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_561),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_531),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_581),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_603),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_481),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_586),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_601),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_393),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_582),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_154),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_265),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_523),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_287),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_287),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_501),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_387),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_597),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_176),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_558),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_48),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_71),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_541),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_407),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_206),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_65),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_292),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_357),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_130),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_425),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_525),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_127),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_402),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_97),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_472),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_226),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_510),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_587),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_274),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_354),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_390),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_465),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_72),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_517),
.Y(n_759)
);

BUFx10_ASAP7_75t_L g760 ( 
.A(n_515),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_390),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_547),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_50),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_372),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_302),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_375),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_144),
.Y(n_767)
);

CKINVDCx16_ASAP7_75t_R g768 ( 
.A(n_598),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_556),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_240),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_16),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_114),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_545),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_58),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_204),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_480),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_240),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_365),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_557),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_232),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_477),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_593),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_479),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_442),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_356),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_475),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_477),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_627),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_605),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_595),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_226),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_383),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_531),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_217),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_361),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_313),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_404),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_520),
.Y(n_798)
);

CKINVDCx16_ASAP7_75t_R g799 ( 
.A(n_594),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_316),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_185),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_15),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_623),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_600),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_164),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_418),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_185),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_398),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_462),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_169),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_111),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_371),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_289),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_587),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_511),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_566),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_101),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_623),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_253),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_458),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_353),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_152),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_242),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_473),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_610),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_433),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_25),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_175),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_620),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_627),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_467),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_187),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_43),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_181),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_315),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_352),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_290),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_65),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_50),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_602),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_98),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_548),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_450),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_60),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_585),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_294),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_151),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_628),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_431),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_125),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_484),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_599),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_289),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_560),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_262),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_117),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_445),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_27),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_10),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_400),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_209),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_606),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_36),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_590),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_422),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_27),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_267),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_207),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_172),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_420),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_418),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_150),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_63),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_192),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_644),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_644),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_768),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_630),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_799),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_644),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_644),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_644),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_802),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_636),
.Y(n_884)
);

BUFx10_ASAP7_75t_L g885 ( 
.A(n_725),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_644),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_644),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_725),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_693),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_658),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_637),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_658),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_633),
.B(n_0),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_638),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_684),
.Y(n_895)
);

INVxp33_ASAP7_75t_L g896 ( 
.A(n_686),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_684),
.Y(n_897)
);

INVx4_ASAP7_75t_R g898 ( 
.A(n_657),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_687),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_725),
.Y(n_900)
);

CKINVDCx14_ASAP7_75t_R g901 ( 
.A(n_718),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_757),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_687),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_784),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_784),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_800),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_800),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_771),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_827),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_825),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_642),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_630),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_825),
.Y(n_913)
);

CKINVDCx14_ASAP7_75t_R g914 ( 
.A(n_760),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_643),
.Y(n_915)
);

CKINVDCx16_ASAP7_75t_R g916 ( 
.A(n_760),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_645),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_725),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_725),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_647),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_679),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_634),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_838),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_838),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_634),
.Y(n_925)
);

INVxp33_ASAP7_75t_SL g926 ( 
.A(n_858),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_682),
.Y(n_927)
);

CKINVDCx16_ASAP7_75t_R g928 ( 
.A(n_760),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_650),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_738),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_738),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_690),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_691),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_738),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_697),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_702),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_706),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_708),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_762),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_738),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_738),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_657),
.B(n_0),
.Y(n_942)
);

BUFx10_ASAP7_75t_L g943 ( 
.A(n_785),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_785),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_650),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_762),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_858),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_710),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_785),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_785),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_785),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_762),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_859),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_810),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_810),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_713),
.Y(n_956)
);

BUFx10_ASAP7_75t_L g957 ( 
.A(n_810),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_676),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_714),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_810),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_716),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_810),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_676),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_719),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_839),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_720),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_839),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_839),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_839),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_839),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_859),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_726),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_733),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_631),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_694),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_632),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_918),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_911),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_918),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_878),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_917),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_877),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_920),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_878),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_912),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_918),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_918),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_912),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_922),
.Y(n_989)
);

INVxp67_ASAP7_75t_SL g990 ( 
.A(n_900),
.Y(n_990)
);

BUFx10_ASAP7_75t_L g991 ( 
.A(n_921),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_919),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_919),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_879),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_919),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_927),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_919),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_922),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_940),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_932),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_876),
.B(n_0),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_941),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_940),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_940),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_925),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_940),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_933),
.B(n_659),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_935),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_936),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_969),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_885),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_937),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_930),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_938),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_925),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_930),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_947),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_972),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_960),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_908),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_909),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_960),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_884),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_929),
.Y(n_1024)
);

NOR2xp67_ASAP7_75t_L g1025 ( 
.A(n_880),
.B(n_1),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_929),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_931),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_939),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_884),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_934),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_891),
.Y(n_1031)
);

INVxp33_ASAP7_75t_SL g1032 ( 
.A(n_891),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_944),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_915),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_949),
.Y(n_1035)
);

INVxp67_ASAP7_75t_SL g1036 ( 
.A(n_882),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_885),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_950),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_895),
.B(n_659),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_951),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_946),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_945),
.Y(n_1042)
);

AND2x6_ASAP7_75t_L g1043 ( 
.A(n_1007),
.B(n_882),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1010),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_990),
.B(n_954),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_1028),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1010),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_977),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_1041),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_1020),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_1011),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_R g1052 ( 
.A1(n_1032),
.A2(n_866),
.B1(n_926),
.B2(n_651),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_999),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_977),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_1021),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_979),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1002),
.B(n_955),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_979),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_1030),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_1011),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1016),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_1037),
.B(n_895),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1016),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1022),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1036),
.B(n_962),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_986),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1022),
.Y(n_1067)
);

INVx6_ASAP7_75t_L g1068 ( 
.A(n_1037),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1017),
.A2(n_948),
.B1(n_956),
.B2(n_915),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_999),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_1030),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_986),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_1039),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_987),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_987),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_992),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_992),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_993),
.B(n_965),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_993),
.B(n_967),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1014),
.A2(n_948),
.B1(n_959),
.B2(n_956),
.Y(n_1080)
);

OA21x2_ASAP7_75t_L g1081 ( 
.A1(n_995),
.A2(n_886),
.B(n_881),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1001),
.B(n_959),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1013),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_995),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1027),
.A2(n_875),
.B(n_887),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1013),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_997),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_997),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_1003),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_978),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_982),
.B(n_971),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1003),
.Y(n_1092)
);

NOR2xp67_ASAP7_75t_L g1093 ( 
.A(n_994),
.B(n_953),
.Y(n_1093)
);

INVx6_ASAP7_75t_L g1094 ( 
.A(n_991),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1004),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1027),
.B(n_1033),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1004),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1006),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1019),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1019),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1006),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1023),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_1033),
.A2(n_875),
.B(n_968),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1035),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1001),
.B(n_1025),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1025),
.B(n_961),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_981),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_980),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1035),
.B(n_970),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1038),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_983),
.B(n_961),
.Y(n_1111)
);

BUFx8_ASAP7_75t_L g1112 ( 
.A(n_1038),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1040),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1040),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_991),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_996),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1029),
.Y(n_1117)
);

AND2x6_ASAP7_75t_L g1118 ( 
.A(n_991),
.B(n_635),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_991),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1031),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1000),
.B(n_964),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1034),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1009),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1012),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1018),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_984),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_985),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_L g1129 ( 
.A(n_988),
.B(n_683),
.Y(n_1129)
);

AND2x6_ASAP7_75t_L g1130 ( 
.A(n_1042),
.B(n_635),
.Y(n_1130)
);

INVx6_ASAP7_75t_L g1131 ( 
.A(n_989),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_SL g1132 ( 
.A1(n_998),
.A2(n_704),
.B1(n_729),
.B2(n_694),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1096),
.Y(n_1133)
);

INVx8_ASAP7_75t_L g1134 ( 
.A(n_1130),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_1050),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1096),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1073),
.B(n_926),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1085),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1061),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1049),
.B(n_914),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_1131),
.B(n_903),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1082),
.A2(n_966),
.B1(n_973),
.B2(n_964),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1082),
.A2(n_973),
.B1(n_966),
.B2(n_901),
.Y(n_1143)
);

AO22x2_ASAP7_75t_L g1144 ( 
.A1(n_1052),
.A2(n_902),
.B1(n_952),
.B2(n_727),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1061),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1063),
.Y(n_1146)
);

OAI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1106),
.A2(n_894),
.B1(n_883),
.B2(n_975),
.Y(n_1147)
);

OAI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1091),
.A2(n_896),
.B1(n_928),
.B2(n_916),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1044),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1091),
.A2(n_942),
.B1(n_893),
.B2(n_804),
.Y(n_1150)
);

XNOR2xp5_ASAP7_75t_L g1151 ( 
.A(n_1050),
.B(n_1005),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1047),
.A2(n_656),
.B1(n_696),
.B2(n_648),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1109),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1051),
.B(n_889),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1063),
.Y(n_1155)
);

XOR2xp5_ASAP7_75t_L g1156 ( 
.A(n_1055),
.B(n_1015),
.Y(n_1156)
);

OAI22xp33_ASAP7_75t_SL g1157 ( 
.A1(n_1106),
.A2(n_866),
.B1(n_727),
.B2(n_728),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1049),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1046),
.B(n_903),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1118),
.A2(n_976),
.B1(n_974),
.B2(n_704),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_SL g1161 ( 
.A1(n_1094),
.A2(n_728),
.B1(n_832),
.B2(n_683),
.Y(n_1161)
);

AOI22x1_ASAP7_75t_L g1162 ( 
.A1(n_1113),
.A2(n_890),
.B1(n_897),
.B2(n_892),
.Y(n_1162)
);

OAI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1046),
.A2(n_817),
.B1(n_819),
.B2(n_721),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1109),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1064),
.Y(n_1165)
);

AO22x2_ASAP7_75t_L g1166 ( 
.A1(n_1052),
.A2(n_832),
.B1(n_820),
.B2(n_826),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1115),
.A2(n_869),
.B1(n_673),
.B2(n_699),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1064),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1109),
.Y(n_1169)
);

AOI22x1_ASAP7_75t_L g1170 ( 
.A1(n_1113),
.A2(n_904),
.B1(n_905),
.B2(n_899),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1115),
.B(n_735),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1108),
.Y(n_1172)
);

AO22x2_ASAP7_75t_L g1173 ( 
.A1(n_1117),
.A2(n_673),
.B1(n_699),
.B2(n_649),
.Y(n_1173)
);

OAI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_1094),
.A2(n_651),
.B1(n_652),
.B2(n_629),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1132),
.A2(n_958),
.B1(n_963),
.B2(n_945),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1053),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1093),
.B(n_906),
.Y(n_1177)
);

OAI22xp33_ASAP7_75t_R g1178 ( 
.A1(n_1127),
.A2(n_639),
.B1(n_646),
.B2(n_640),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1118),
.A2(n_770),
.B1(n_816),
.B2(n_759),
.Y(n_1179)
);

OAI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1094),
.A2(n_652),
.B1(n_655),
.B2(n_629),
.Y(n_1180)
);

OAI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1115),
.A2(n_649),
.B1(n_730),
.B2(n_701),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1124),
.B(n_907),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1067),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1118),
.A2(n_1043),
.B1(n_1105),
.B2(n_1065),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1104),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1121),
.B(n_958),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1118),
.A2(n_824),
.B1(n_830),
.B2(n_816),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1118),
.A2(n_830),
.B1(n_836),
.B2(n_824),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1062),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1053),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1069),
.B(n_963),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1094),
.A2(n_1111),
.B1(n_1123),
.B2(n_1120),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1043),
.A2(n_841),
.B1(n_856),
.B2(n_836),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1110),
.Y(n_1194)
);

OR2x6_ASAP7_75t_L g1195 ( 
.A(n_1131),
.B(n_910),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1067),
.Y(n_1196)
);

OA22x2_ASAP7_75t_L g1197 ( 
.A1(n_1080),
.A2(n_753),
.B1(n_857),
.B2(n_670),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1043),
.A2(n_856),
.B1(n_841),
.B2(n_913),
.Y(n_1198)
);

AO22x2_ASAP7_75t_L g1199 ( 
.A1(n_1111),
.A2(n_850),
.B1(n_701),
.B2(n_779),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1043),
.A2(n_924),
.B1(n_923),
.B2(n_737),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1108),
.B(n_655),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1124),
.A2(n_663),
.B1(n_669),
.B2(n_661),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1131),
.A2(n_1026),
.B1(n_1024),
.B2(n_669),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1131),
.A2(n_670),
.B1(n_753),
.B2(n_661),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1128),
.B(n_730),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1114),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1113),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1124),
.B(n_898),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1085),
.Y(n_1209)
);

OAI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1125),
.A2(n_764),
.B1(n_855),
.B2(n_663),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1055),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1125),
.A2(n_855),
.B1(n_857),
.B2(n_764),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1043),
.A2(n_739),
.B1(n_740),
.B2(n_736),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1083),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1083),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1103),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1128),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1051),
.B(n_653),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1103),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1125),
.B(n_744),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1086),
.Y(n_1221)
);

OA22x2_ASAP7_75t_L g1222 ( 
.A1(n_1126),
.A2(n_861),
.B1(n_863),
.B2(n_860),
.Y(n_1222)
);

OAI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1115),
.A2(n_801),
.B1(n_814),
.B2(n_779),
.Y(n_1223)
);

NAND2xp33_ASAP7_75t_SL g1224 ( 
.A(n_1122),
.B(n_860),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1060),
.B(n_654),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1105),
.B(n_885),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1043),
.A2(n_746),
.B1(n_747),
.B2(n_745),
.Y(n_1227)
);

NAND3x1_ASAP7_75t_L g1228 ( 
.A(n_1130),
.B(n_680),
.C(n_667),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1105),
.A2(n_752),
.B1(n_754),
.B2(n_748),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1086),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_R g1231 ( 
.A1(n_1122),
.A2(n_660),
.B1(n_664),
.B2(n_662),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1060),
.B(n_755),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1099),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1068),
.A2(n_863),
.B1(n_864),
.B2(n_861),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1116),
.B(n_758),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1099),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1116),
.B(n_763),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1100),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1102),
.B(n_765),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1115),
.A2(n_814),
.B1(n_850),
.B2(n_801),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1119),
.B(n_766),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1130),
.B(n_665),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1045),
.A2(n_1057),
.B1(n_1130),
.B2(n_1068),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1130),
.A2(n_772),
.B1(n_773),
.B2(n_769),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1130),
.A2(n_778),
.B1(n_780),
.B2(n_774),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1100),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1068),
.B(n_781),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1128),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1119),
.B(n_782),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1053),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_SL g1251 ( 
.A1(n_1090),
.A2(n_865),
.B1(n_867),
.B2(n_864),
.Y(n_1251)
);

AO22x2_ASAP7_75t_L g1252 ( 
.A1(n_1129),
.A2(n_666),
.B1(n_671),
.B2(n_668),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1068),
.A2(n_788),
.B1(n_789),
.B2(n_783),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1048),
.A2(n_791),
.B1(n_793),
.B2(n_790),
.Y(n_1254)
);

AOI22x1_ASAP7_75t_L g1255 ( 
.A1(n_1092),
.A2(n_867),
.B1(n_870),
.B2(n_865),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1119),
.A2(n_672),
.B1(n_675),
.B2(n_674),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1054),
.A2(n_797),
.B1(n_798),
.B2(n_796),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1056),
.A2(n_805),
.B1(n_806),
.B2(n_803),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1058),
.A2(n_808),
.B1(n_809),
.B2(n_807),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1103),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1066),
.B(n_888),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1072),
.A2(n_812),
.B1(n_813),
.B2(n_811),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1119),
.B(n_815),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1078),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1119),
.A2(n_871),
.B1(n_872),
.B2(n_870),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1128),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1090),
.A2(n_872),
.B1(n_873),
.B2(n_871),
.Y(n_1267)
);

AO22x2_ASAP7_75t_L g1268 ( 
.A1(n_1129),
.A2(n_677),
.B1(n_681),
.B2(n_678),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1079),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1092),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1264),
.B(n_1269),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1159),
.B(n_1137),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1260),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1182),
.B(n_1075),
.Y(n_1274)
);

INVx5_ASAP7_75t_L g1275 ( 
.A(n_1134),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1133),
.A2(n_1077),
.B1(n_1084),
.B2(n_1076),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1192),
.B(n_1107),
.Y(n_1277)
);

XNOR2xp5_ASAP7_75t_L g1278 ( 
.A(n_1151),
.B(n_1107),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1208),
.B(n_873),
.Y(n_1279)
);

OAI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1198),
.A2(n_685),
.B1(n_689),
.B2(n_688),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1158),
.B(n_818),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1221),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1176),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1184),
.B(n_1053),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1236),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1217),
.B(n_1087),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1193),
.B(n_1095),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1149),
.B(n_1097),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1177),
.B(n_1098),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1154),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1136),
.B(n_1059),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1176),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1185),
.B(n_1059),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1243),
.B(n_1070),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1216),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1154),
.Y(n_1296)
);

BUFx8_ASAP7_75t_SL g1297 ( 
.A(n_1211),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1207),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1190),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_SL g1300 ( 
.A(n_1140),
.B(n_1070),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1214),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1194),
.B(n_1059),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1248),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1216),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1206),
.B(n_1071),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1199),
.A2(n_1081),
.B1(n_692),
.B2(n_698),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1138),
.A2(n_700),
.B(n_695),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1215),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1270),
.Y(n_1309)
);

INVx4_ASAP7_75t_L g1310 ( 
.A(n_1134),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1199),
.A2(n_1081),
.B1(n_703),
.B2(n_707),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1235),
.B(n_823),
.Y(n_1312)
);

AND2x6_ASAP7_75t_L g1313 ( 
.A(n_1219),
.B(n_1092),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1190),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1160),
.B(n_1070),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1266),
.B(n_1218),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1186),
.B(n_1071),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1219),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1230),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1205),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1250),
.Y(n_1321)
);

AND2x2_ASAP7_75t_SL g1322 ( 
.A(n_1179),
.B(n_1081),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1233),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1135),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1238),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1200),
.B(n_1070),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1220),
.B(n_1071),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1135),
.Y(n_1328)
);

XNOR2xp5_ASAP7_75t_L g1329 ( 
.A(n_1156),
.B(n_1112),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1231),
.A2(n_1178),
.B1(n_1173),
.B2(n_1197),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1246),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1153),
.B(n_1074),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1138),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1164),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1187),
.B(n_1074),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1201),
.B(n_828),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1141),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1250),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1209),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1188),
.B(n_1074),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1231),
.A2(n_705),
.B1(n_711),
.B2(n_709),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1169),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1139),
.Y(n_1343)
);

OR2x6_ASAP7_75t_L g1344 ( 
.A(n_1172),
.B(n_1112),
.Y(n_1344)
);

OAI21xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1209),
.A2(n_715),
.B(n_712),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1147),
.B(n_1074),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1145),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1141),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1226),
.B(n_1157),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1195),
.B(n_829),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1146),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1155),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1242),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1195),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1178),
.A2(n_717),
.B1(n_723),
.B2(n_722),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1165),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1168),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1183),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1196),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1162),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1218),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1162),
.Y(n_1362)
);

INVx5_ASAP7_75t_L g1363 ( 
.A(n_1242),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1170),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1225),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1225),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1205),
.Y(n_1367)
);

OR2x6_ASAP7_75t_L g1368 ( 
.A(n_1228),
.B(n_1112),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1170),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1173),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1255),
.Y(n_1371)
);

NAND2xp33_ASAP7_75t_L g1372 ( 
.A(n_1241),
.B(n_1249),
.Y(n_1372)
);

AND3x1_ASAP7_75t_L g1373 ( 
.A(n_1191),
.B(n_731),
.C(n_724),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1175),
.B(n_732),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1189),
.B(n_734),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1255),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1261),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1222),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1213),
.B(n_1227),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1203),
.B(n_833),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1247),
.B(n_1088),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1232),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1181),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1263),
.B(n_1088),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1142),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1223),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1171),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1240),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1252),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1150),
.B(n_1088),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1237),
.B(n_834),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1252),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1239),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1268),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1143),
.B(n_835),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1268),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1144),
.B(n_741),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1144),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1166),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1167),
.B(n_1088),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1224),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1166),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1174),
.B(n_1089),
.Y(n_1403)
);

AND2x2_ASAP7_75t_SL g1404 ( 
.A(n_1244),
.B(n_742),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1161),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1254),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1229),
.B(n_842),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1202),
.B(n_1089),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1210),
.B(n_1089),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1256),
.Y(n_1410)
);

BUFx10_ASAP7_75t_L g1411 ( 
.A(n_1265),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1245),
.A2(n_1101),
.B1(n_1089),
.B2(n_845),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1180),
.B(n_1234),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1253),
.B(n_844),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1257),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1212),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1148),
.B(n_1101),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1258),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1163),
.A2(n_743),
.B1(n_750),
.B2(n_749),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1204),
.B(n_751),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1259),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1262),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1152),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1251),
.B(n_1101),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1267),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_SL g1426 ( 
.A(n_1211),
.B(n_849),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1217),
.B(n_756),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1176),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1137),
.B(n_1101),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1134),
.Y(n_1430)
);

INVx5_ASAP7_75t_L g1431 ( 
.A(n_1134),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1221),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1221),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1192),
.B(n_888),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1260),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1158),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1192),
.B(n_888),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1270),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1192),
.B(n_943),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1221),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1134),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1264),
.B(n_851),
.Y(n_1442)
);

AND2x6_ASAP7_75t_L g1443 ( 
.A(n_1260),
.B(n_761),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1260),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1264),
.B(n_852),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1217),
.Y(n_1446)
);

BUFx8_ASAP7_75t_SL g1447 ( 
.A(n_1211),
.Y(n_1447)
);

OAI21xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1149),
.A2(n_775),
.B(n_767),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1134),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1199),
.A2(n_776),
.B1(n_786),
.B2(n_777),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1221),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1260),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1221),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1221),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1221),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1260),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1264),
.B(n_853),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1134),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1176),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1270),
.Y(n_1460)
);

AND2x6_ASAP7_75t_L g1461 ( 
.A(n_1260),
.B(n_787),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1260),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1158),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1159),
.B(n_854),
.Y(n_1464)
);

BUFx4f_ASAP7_75t_L g1465 ( 
.A(n_1141),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1264),
.B(n_792),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1216),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1260),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1264),
.B(n_794),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1260),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1221),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1264),
.B(n_795),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1271),
.A2(n_821),
.B1(n_831),
.B2(n_822),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1297),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1272),
.B(n_943),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1356),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1295),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1464),
.B(n_837),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1295),
.Y(n_1479)
);

INVx8_ASAP7_75t_L g1480 ( 
.A(n_1313),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1297),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1366),
.B(n_840),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1304),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1304),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1366),
.B(n_843),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1358),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1418),
.B(n_943),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1318),
.Y(n_1488)
);

BUFx10_ASAP7_75t_L g1489 ( 
.A(n_1328),
.Y(n_1489)
);

NAND2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1275),
.B(n_1431),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1316),
.B(n_846),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1382),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1316),
.B(n_847),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1467),
.B(n_848),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1320),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1318),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1436),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1334),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1358),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1273),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1282),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1467),
.B(n_862),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1385),
.B(n_1),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1446),
.B(n_868),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1404),
.A2(n_874),
.B1(n_957),
.B2(n_641),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1285),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1432),
.Y(n_1507)
);

INVx6_ASAP7_75t_L g1508 ( 
.A(n_1324),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1273),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1446),
.B(n_34),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1361),
.B(n_35),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1374),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1430),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1336),
.B(n_1442),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1433),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1447),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1440),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1463),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1451),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1430),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1365),
.B(n_35),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1430),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1404),
.A2(n_957),
.B1(n_4),
.B2(n_2),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1429),
.B(n_2),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1342),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1312),
.B(n_957),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1453),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1377),
.B(n_613),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1454),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1435),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1391),
.B(n_613),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1342),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1435),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1455),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1320),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1471),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1429),
.B(n_3),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1430),
.Y(n_1538)
);

INVx5_ASAP7_75t_L g1539 ( 
.A(n_1447),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1290),
.B(n_36),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1279),
.B(n_615),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1352),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1450),
.A2(n_1392),
.B1(n_1389),
.B2(n_1311),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1296),
.B(n_37),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1324),
.Y(n_1545)
);

AND2x2_ASAP7_75t_SL g1546 ( 
.A(n_1465),
.B(n_1373),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1342),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1359),
.Y(n_1548)
);

NAND2x1p5_ASAP7_75t_L g1549 ( 
.A(n_1275),
.B(n_37),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1444),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1444),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1452),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1452),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1456),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1421),
.B(n_616),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1456),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1462),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1450),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1317),
.B(n_4),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1393),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1462),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1468),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1468),
.Y(n_1563)
);

AND2x6_ASAP7_75t_L g1564 ( 
.A(n_1441),
.B(n_5),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1281),
.B(n_618),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1395),
.B(n_618),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1286),
.B(n_38),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1441),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1278),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1470),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1317),
.B(n_5),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1470),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1441),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1421),
.B(n_621),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1367),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1441),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1343),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1301),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1329),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1389),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1308),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1286),
.B(n_38),
.Y(n_1582)
);

AND2x6_ASAP7_75t_L g1583 ( 
.A(n_1458),
.B(n_6),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1343),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1303),
.B(n_39),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1319),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1422),
.B(n_622),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1323),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1357),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1303),
.B(n_39),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1458),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1357),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1347),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1354),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1287),
.B(n_6),
.C(n_7),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1351),
.Y(n_1596)
);

AND2x6_ASAP7_75t_L g1597 ( 
.A(n_1458),
.B(n_7),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1325),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1427),
.B(n_626),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1331),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1333),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1354),
.B(n_40),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1422),
.B(n_626),
.Y(n_1603)
);

INVx8_ASAP7_75t_L g1604 ( 
.A(n_1313),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1298),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1333),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1274),
.B(n_8),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1418),
.B(n_40),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1337),
.B(n_41),
.Y(n_1609)
);

INVx4_ASAP7_75t_L g1610 ( 
.A(n_1458),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1339),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1367),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1427),
.B(n_628),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1339),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1288),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1275),
.B(n_41),
.Y(n_1616)
);

AND2x6_ASAP7_75t_L g1617 ( 
.A(n_1392),
.B(n_8),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1287),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1393),
.B(n_610),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1309),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1438),
.Y(n_1621)
);

INVx6_ASAP7_75t_L g1622 ( 
.A(n_1344),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1460),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1276),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1332),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1342),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1289),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1393),
.B(n_611),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1291),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1353),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1465),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1283),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1419),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1344),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1344),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1401),
.B(n_42),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1401),
.B(n_42),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1375),
.B(n_612),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1445),
.B(n_43),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1378),
.B(n_44),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1375),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1353),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1378),
.B(n_1387),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1407),
.B(n_614),
.Y(n_1644)
);

AO22x2_ASAP7_75t_L g1645 ( 
.A1(n_1399),
.A2(n_1402),
.B1(n_1398),
.B2(n_1396),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1350),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1387),
.B(n_44),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1275),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1283),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1418),
.B(n_45),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1387),
.B(n_45),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1457),
.B(n_616),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1419),
.A2(n_1330),
.B1(n_1394),
.B2(n_1341),
.C(n_1423),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1418),
.B(n_617),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1292),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1410),
.B(n_46),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1348),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1292),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1327),
.B(n_9),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1406),
.B(n_617),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1299),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1387),
.B(n_46),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1353),
.Y(n_1663)
);

AND2x6_ASAP7_75t_L g1664 ( 
.A(n_1353),
.B(n_9),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1299),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1466),
.B(n_10),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1469),
.B(n_11),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1314),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1322),
.Y(n_1669)
);

BUFx10_ASAP7_75t_L g1670 ( 
.A(n_1346),
.Y(n_1670)
);

INVx6_ASAP7_75t_L g1671 ( 
.A(n_1411),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1314),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1321),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1405),
.B(n_47),
.Y(n_1674)
);

BUFx4f_ASAP7_75t_L g1675 ( 
.A(n_1410),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1414),
.B(n_624),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1406),
.B(n_1415),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1322),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1321),
.Y(n_1679)
);

BUFx4f_ASAP7_75t_L g1680 ( 
.A(n_1410),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1330),
.B(n_624),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1652),
.B(n_1654),
.C(n_1574),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1675),
.B(n_1426),
.Y(n_1683)
);

INVx5_ASAP7_75t_L g1684 ( 
.A(n_1480),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1618),
.B(n_1472),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1508),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1627),
.B(n_1335),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1675),
.B(n_1410),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1618),
.B(n_1425),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1646),
.A2(n_1277),
.B1(n_1372),
.B2(n_1380),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1615),
.B(n_1335),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1676),
.A2(n_1416),
.B1(n_1415),
.B2(n_1379),
.Y(n_1692)
);

INVx8_ASAP7_75t_L g1693 ( 
.A(n_1513),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1677),
.B(n_1340),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1481),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1625),
.B(n_1680),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1680),
.B(n_1340),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1606),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1514),
.B(n_1416),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1653),
.B(n_1398),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1555),
.A2(n_1277),
.B1(n_1374),
.B2(n_1349),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1653),
.B(n_1399),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1575),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1503),
.A2(n_1374),
.B1(n_1420),
.B2(n_1397),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1611),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1478),
.B(n_1397),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1624),
.B(n_1629),
.Y(n_1707)
);

AOI22x1_ASAP7_75t_L g1708 ( 
.A1(n_1526),
.A2(n_1376),
.B1(n_1371),
.B2(n_1362),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1614),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1500),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1601),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1509),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1513),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1546),
.B(n_1641),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_SL g1715 ( 
.A(n_1503),
.B(n_1355),
.C(n_1341),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1492),
.B(n_1405),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1566),
.B(n_1370),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_SL g1718 ( 
.A(n_1633),
.B(n_1431),
.Y(n_1718)
);

O2A1O1Ixp5_ASAP7_75t_L g1719 ( 
.A1(n_1559),
.A2(n_1379),
.B(n_1349),
.C(n_1417),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1670),
.B(n_1416),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1498),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1670),
.B(n_1560),
.Y(n_1722)
);

INVxp67_ASAP7_75t_SL g1723 ( 
.A(n_1495),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1560),
.B(n_1280),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1644),
.B(n_1346),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1607),
.B(n_1408),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1643),
.B(n_1497),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1607),
.B(n_1408),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1501),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1506),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1523),
.A2(n_1409),
.B1(n_1413),
.B2(n_1420),
.Y(n_1731)
);

NOR2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1631),
.B(n_1390),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1660),
.B(n_1409),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1523),
.A2(n_1413),
.B1(n_1420),
.B2(n_1411),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1535),
.B(n_1612),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1666),
.B(n_1383),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1508),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1530),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1545),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1513),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1612),
.B(n_1424),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1480),
.A2(n_1381),
.B(n_1384),
.Y(n_1742)
);

AND2x6_ASAP7_75t_SL g1743 ( 
.A(n_1602),
.B(n_1397),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1666),
.B(n_1386),
.Y(n_1744)
);

NOR2x1p5_ASAP7_75t_L g1745 ( 
.A(n_1474),
.B(n_1388),
.Y(n_1745)
);

NOR2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1516),
.B(n_1400),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1507),
.Y(n_1747)
);

O2A1O1Ixp5_ASAP7_75t_L g1748 ( 
.A1(n_1559),
.A2(n_1417),
.B(n_1439),
.C(n_1437),
.Y(n_1748)
);

INVx5_ASAP7_75t_L g1749 ( 
.A(n_1480),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1667),
.B(n_1293),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1533),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1551),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1553),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1543),
.B(n_1306),
.Y(n_1754)
);

AO22x1_ASAP7_75t_L g1755 ( 
.A1(n_1558),
.A2(n_1363),
.B1(n_1371),
.B2(n_1443),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1657),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1667),
.B(n_1302),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1561),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1587),
.A2(n_1603),
.B(n_1505),
.C(n_1528),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1681),
.B(n_1305),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1543),
.B(n_1424),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1531),
.B(n_1306),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_SL g1763 ( 
.A1(n_1512),
.A2(n_1368),
.B1(n_1363),
.B2(n_1431),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1639),
.B(n_1311),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1494),
.B(n_1363),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1569),
.B(n_1403),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1594),
.Y(n_1767)
);

BUFx8_ASAP7_75t_L g1768 ( 
.A(n_1602),
.Y(n_1768)
);

AND2x4_ASAP7_75t_SL g1769 ( 
.A(n_1489),
.B(n_1310),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1494),
.B(n_1363),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1502),
.B(n_1448),
.Y(n_1771)
);

NAND2x1p5_ASAP7_75t_L g1772 ( 
.A(n_1648),
.B(n_1431),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1495),
.B(n_1434),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1640),
.B(n_1355),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1608),
.A2(n_1300),
.B1(n_1437),
.B2(n_1434),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1502),
.B(n_1643),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1671),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1515),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1518),
.B(n_1439),
.Y(n_1779)
);

OAI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1633),
.A2(n_1368),
.B1(n_1310),
.B2(n_1449),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1619),
.B(n_1459),
.Y(n_1781)
);

O2A1O1Ixp5_ASAP7_75t_L g1782 ( 
.A1(n_1571),
.A2(n_1326),
.B(n_1294),
.C(n_1315),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1640),
.B(n_1368),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1669),
.A2(n_1315),
.B1(n_1449),
.B2(n_1360),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1604),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1477),
.B(n_1443),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1517),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1671),
.A2(n_1412),
.B1(n_1284),
.B2(n_1443),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1475),
.A2(n_1284),
.B1(n_1461),
.B2(n_1443),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1519),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1604),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1510),
.B(n_1628),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1650),
.A2(n_1461),
.B1(n_1443),
.B2(n_1307),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1524),
.B(n_1461),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1656),
.A2(n_1461),
.B1(n_1307),
.B2(n_1294),
.Y(n_1795)
);

NAND2x1_ASAP7_75t_L g1796 ( 
.A(n_1538),
.B(n_1313),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1585),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1479),
.B(n_1461),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1524),
.B(n_1338),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1510),
.B(n_1338),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1483),
.B(n_1428),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1635),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1636),
.B(n_1428),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1638),
.B(n_1541),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1527),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1585),
.B(n_1459),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1558),
.A2(n_1345),
.B(n_1326),
.C(n_1364),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1529),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1604),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1565),
.A2(n_1313),
.B1(n_1369),
.B2(n_1360),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1534),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1536),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_SL g1813 ( 
.A1(n_1512),
.A2(n_1313),
.B1(n_48),
.B2(n_49),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1537),
.B(n_11),
.Y(n_1814)
);

INVx5_ASAP7_75t_L g1815 ( 
.A(n_1520),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1484),
.Y(n_1816)
);

A2O1A1Ixp33_ASAP7_75t_L g1817 ( 
.A1(n_1571),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1537),
.B(n_12),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1488),
.B(n_1496),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1674),
.A2(n_49),
.B1(n_51),
.B2(n_47),
.Y(n_1820)
);

INVx8_ASAP7_75t_L g1821 ( 
.A(n_1520),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1563),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1570),
.B(n_13),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1636),
.B(n_1637),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1637),
.B(n_51),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1605),
.Y(n_1826)
);

INVxp33_ASAP7_75t_L g1827 ( 
.A(n_1504),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1550),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1552),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1622),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1659),
.B(n_13),
.Y(n_1831)
);

AO22x1_ASAP7_75t_L g1832 ( 
.A1(n_1664),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1599),
.B(n_609),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1504),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1659),
.B(n_14),
.Y(n_1835)
);

OR2x6_ASAP7_75t_L g1836 ( 
.A(n_1622),
.B(n_52),
.Y(n_1836)
);

NAND2xp33_ASAP7_75t_L g1837 ( 
.A(n_1630),
.B(n_1642),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1554),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1567),
.B(n_52),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1556),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1557),
.B(n_15),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1669),
.B(n_53),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1678),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1539),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1542),
.B(n_17),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1476),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1548),
.B(n_1578),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1595),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1539),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1678),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1487),
.A2(n_54),
.B(n_53),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1590),
.B(n_54),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1590),
.B(n_55),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1595),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1581),
.B(n_20),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1674),
.A2(n_56),
.B1(n_57),
.B2(n_55),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1586),
.B(n_21),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1486),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1499),
.Y(n_1859)
);

NOR3xp33_ASAP7_75t_L g1860 ( 
.A(n_1473),
.B(n_22),
.C(n_23),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1588),
.B(n_22),
.Y(n_1861)
);

INVxp33_ASAP7_75t_L g1862 ( 
.A(n_1491),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1482),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1562),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1613),
.B(n_607),
.Y(n_1865)
);

XNOR2xp5_ASAP7_75t_L g1866 ( 
.A(n_1579),
.B(n_56),
.Y(n_1866)
);

NAND2xp33_ASAP7_75t_L g1867 ( 
.A(n_1630),
.B(n_23),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1490),
.A2(n_59),
.B(n_57),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1572),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_1525),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1567),
.B(n_609),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1490),
.A2(n_60),
.B(n_59),
.Y(n_1872)
);

AND2x6_ASAP7_75t_SL g1873 ( 
.A(n_1609),
.B(n_24),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1598),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1715),
.B(n_1682),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1686),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1874),
.Y(n_1877)
);

AND3x1_ASAP7_75t_SL g1878 ( 
.A(n_1746),
.B(n_1600),
.C(n_1626),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1694),
.B(n_1525),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1710),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1759),
.B(n_1647),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1712),
.Y(n_1882)
);

CKINVDCx16_ASAP7_75t_R g1883 ( 
.A(n_1756),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1738),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_1695),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1697),
.B(n_1647),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1684),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1847),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1721),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1733),
.B(n_1651),
.Y(n_1890)
);

OR2x2_ASAP7_75t_SL g1891 ( 
.A(n_1725),
.B(n_1593),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1726),
.B(n_1482),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1694),
.B(n_1532),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1729),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1860),
.A2(n_1580),
.B1(n_1664),
.B2(n_1617),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1730),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1751),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1752),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1728),
.B(n_1485),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1777),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1747),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1797),
.B(n_1582),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1737),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1723),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1778),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1685),
.B(n_1485),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1787),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1691),
.B(n_1532),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1790),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1802),
.Y(n_1910)
);

A2O1A1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1701),
.A2(n_1651),
.B(n_1662),
.C(n_1473),
.Y(n_1911)
);

BUFx3_ASAP7_75t_L g1912 ( 
.A(n_1768),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1805),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1697),
.B(n_1662),
.Y(n_1914)
);

AO22x1_ASAP7_75t_L g1915 ( 
.A1(n_1843),
.A2(n_1664),
.B1(n_1564),
.B2(n_1597),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1848),
.A2(n_1580),
.B1(n_1664),
.B2(n_1617),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1768),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1808),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1753),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1691),
.B(n_1547),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1693),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1687),
.B(n_1547),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1774),
.B(n_1582),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1731),
.A2(n_1645),
.B1(n_1521),
.B2(n_1511),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1758),
.Y(n_1925)
);

INVx2_ASAP7_75t_SL g1926 ( 
.A(n_1739),
.Y(n_1926)
);

AND2x6_ASAP7_75t_L g1927 ( 
.A(n_1785),
.B(n_1511),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1846),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1811),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1687),
.B(n_1645),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1776),
.Y(n_1931)
);

BUFx4f_ASAP7_75t_L g1932 ( 
.A(n_1693),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1684),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1812),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1690),
.B(n_1630),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1826),
.Y(n_1936)
);

O2A1O1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1817),
.A2(n_1521),
.B(n_1621),
.C(n_1620),
.Y(n_1937)
);

BUFx4f_ASAP7_75t_L g1938 ( 
.A(n_1693),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1828),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1797),
.B(n_1642),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1717),
.B(n_1623),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1829),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1732),
.B(n_1642),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1838),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1858),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1854),
.A2(n_1617),
.B1(n_1583),
.B2(n_1597),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1830),
.B(n_1663),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1840),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1864),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1869),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1767),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1745),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1761),
.B(n_1617),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1736),
.B(n_1649),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1711),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1744),
.B(n_1649),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1821),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1859),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1698),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1794),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1705),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1760),
.B(n_1655),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1792),
.B(n_1663),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1821),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1783),
.B(n_1663),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1709),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1707),
.B(n_1700),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_SL g1968 ( 
.A(n_1718),
.B(n_1539),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1702),
.B(n_1655),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1834),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1816),
.Y(n_1971)
);

OR2x4_ASAP7_75t_L g1972 ( 
.A(n_1766),
.B(n_1520),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1804),
.B(n_1491),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1822),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1750),
.B(n_1577),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1704),
.A2(n_1634),
.B1(n_1493),
.B2(n_1489),
.Y(n_1976)
);

BUFx2_ASAP7_75t_L g1977 ( 
.A(n_1703),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1684),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1819),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1821),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1819),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1696),
.B(n_1584),
.Y(n_1982)
);

BUFx8_ASAP7_75t_SL g1983 ( 
.A(n_1844),
.Y(n_1983)
);

BUFx4f_ASAP7_75t_L g1984 ( 
.A(n_1713),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1801),
.Y(n_1985)
);

INVx5_ASAP7_75t_L g1986 ( 
.A(n_1815),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1757),
.B(n_1589),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1800),
.B(n_1538),
.Y(n_1988)
);

INVx2_ASAP7_75t_SL g1989 ( 
.A(n_1703),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1735),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1684),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1823),
.Y(n_1992)
);

BUFx12f_ASAP7_75t_L g1993 ( 
.A(n_1849),
.Y(n_1993)
);

BUFx8_ASAP7_75t_L g1994 ( 
.A(n_1689),
.Y(n_1994)
);

INVx2_ASAP7_75t_SL g1995 ( 
.A(n_1769),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1801),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1713),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1683),
.A2(n_1493),
.B1(n_1544),
.B2(n_1540),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1706),
.A2(n_1540),
.B1(n_1544),
.B2(n_1564),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1873),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1754),
.B(n_1592),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1754),
.B(n_1665),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1696),
.B(n_1596),
.Y(n_2003)
);

NAND2xp33_ASAP7_75t_SL g2004 ( 
.A(n_1827),
.B(n_1522),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1713),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1823),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1799),
.B(n_1673),
.Y(n_2007)
);

INVx5_ASAP7_75t_L g2008 ( 
.A(n_1815),
.Y(n_2008)
);

NOR2x1p5_ASAP7_75t_L g2009 ( 
.A(n_1764),
.B(n_1610),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1727),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1786),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1749),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1824),
.B(n_1609),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1740),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1786),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1815),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1688),
.B(n_1679),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1798),
.Y(n_2018)
);

AOI221xp5_ASAP7_75t_SL g2019 ( 
.A1(n_1843),
.A2(n_1661),
.B1(n_1668),
.B2(n_1658),
.C(n_1632),
.Y(n_2019)
);

INVx3_ASAP7_75t_SL g2020 ( 
.A(n_1836),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1798),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1841),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1749),
.B(n_1610),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1749),
.B(n_1522),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1841),
.Y(n_2025)
);

AND2x6_ASAP7_75t_L g2026 ( 
.A(n_1785),
.B(n_1522),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1692),
.B(n_1616),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1740),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1845),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1749),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1740),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1813),
.A2(n_1616),
.B1(n_1549),
.B2(n_1672),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1839),
.Y(n_2033)
);

OR2x6_ASAP7_75t_L g2034 ( 
.A(n_1755),
.B(n_1549),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1839),
.Y(n_2035)
);

BUFx8_ASAP7_75t_L g2036 ( 
.A(n_1871),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1741),
.B(n_1568),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1722),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1791),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1743),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1833),
.B(n_1564),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1855),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1719),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1857),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_1850),
.A2(n_1583),
.B1(n_1597),
.B2(n_1564),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1875),
.A2(n_1734),
.B1(n_1867),
.B2(n_1699),
.Y(n_2046)
);

NOR2xp67_ASAP7_75t_L g2047 ( 
.A(n_1995),
.B(n_1779),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1881),
.A2(n_1742),
.B(n_1807),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1972),
.A2(n_1763),
.B1(n_1716),
.B2(n_1714),
.Y(n_2049)
);

AOI21xp33_ASAP7_75t_L g2050 ( 
.A1(n_1875),
.A2(n_1771),
.B(n_1814),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_1883),
.B(n_1862),
.Y(n_2051)
);

O2A1O1Ixp5_ASAP7_75t_L g2052 ( 
.A1(n_1881),
.A2(n_1832),
.B(n_1748),
.C(n_1720),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1967),
.B(n_1818),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1889),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1885),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_1876),
.Y(n_2056)
);

O2A1O1Ixp33_ASAP7_75t_L g2057 ( 
.A1(n_1911),
.A2(n_1724),
.B(n_1853),
.C(n_1850),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1967),
.B(n_1831),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1968),
.B(n_1765),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1968),
.B(n_1770),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1931),
.B(n_1835),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1894),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_R g2063 ( 
.A(n_1932),
.B(n_1837),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1931),
.B(n_1842),
.Y(n_2064)
);

AOI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_2034),
.A2(n_1718),
.B(n_1782),
.Y(n_2065)
);

NOR3xp33_ASAP7_75t_L g2066 ( 
.A(n_2032),
.B(n_1762),
.C(n_1780),
.Y(n_2066)
);

AOI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1886),
.A2(n_1914),
.B1(n_2009),
.B2(n_1890),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1973),
.B(n_1866),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1892),
.B(n_1788),
.Y(n_2069)
);

AOI22x1_ASAP7_75t_L g2070 ( 
.A1(n_2022),
.A2(n_1851),
.B1(n_1872),
.B2(n_1868),
.Y(n_2070)
);

CKINVDCx20_ASAP7_75t_R g2071 ( 
.A(n_1983),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2029),
.B(n_1773),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2034),
.A2(n_1784),
.B(n_1708),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1877),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1880),
.Y(n_2075)
);

INVx2_ASAP7_75t_SL g2076 ( 
.A(n_1910),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1960),
.B(n_1861),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2034),
.A2(n_1784),
.B(n_1775),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1890),
.A2(n_1795),
.B(n_1793),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1899),
.B(n_1789),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1882),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_1886),
.A2(n_1825),
.B1(n_1852),
.B2(n_1820),
.Y(n_2082)
);

O2A1O1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_1935),
.A2(n_1806),
.B(n_1836),
.C(n_1781),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2042),
.B(n_1803),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1896),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1901),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1884),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_2027),
.A2(n_1810),
.B(n_1796),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1906),
.B(n_2044),
.Y(n_2089)
);

AOI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_2027),
.A2(n_1870),
.B(n_1772),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2043),
.A2(n_1772),
.B(n_1791),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1937),
.A2(n_1856),
.B(n_1863),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_L g2093 ( 
.A1(n_1916),
.A2(n_1597),
.B1(n_1583),
.B2(n_1836),
.Y(n_2093)
);

O2A1O1Ixp33_ASAP7_75t_L g2094 ( 
.A1(n_1935),
.A2(n_1865),
.B(n_1809),
.C(n_1583),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1897),
.Y(n_2095)
);

A2O1A1Ixp33_ASAP7_75t_L g2096 ( 
.A1(n_1937),
.A2(n_1809),
.B(n_1573),
.C(n_1576),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1905),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_1914),
.B(n_1568),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_1981),
.A2(n_2008),
.B(n_1986),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1888),
.B(n_1573),
.Y(n_2100)
);

AOI211xp5_ASAP7_75t_L g2101 ( 
.A1(n_1915),
.A2(n_1591),
.B(n_1576),
.C(n_26),
.Y(n_2101)
);

INVxp67_ASAP7_75t_L g2102 ( 
.A(n_1977),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_1916),
.A2(n_1591),
.B1(n_26),
.B2(n_24),
.Y(n_2103)
);

AO21x1_ASAP7_75t_L g2104 ( 
.A1(n_1924),
.A2(n_25),
.B(n_26),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_1979),
.A2(n_1591),
.B(n_62),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1992),
.B(n_61),
.Y(n_2106)
);

AOI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1954),
.A2(n_63),
.B(n_62),
.Y(n_2107)
);

O2A1O1Ixp33_ASAP7_75t_L g2108 ( 
.A1(n_2032),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1990),
.B(n_2013),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1923),
.B(n_64),
.Y(n_2110)
);

INVx4_ASAP7_75t_L g2111 ( 
.A(n_1986),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2006),
.B(n_64),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2025),
.B(n_66),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1990),
.B(n_66),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_2038),
.B(n_67),
.Y(n_2115)
);

AOI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_1952),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2116)
);

NAND3xp33_ASAP7_75t_L g2117 ( 
.A(n_1895),
.B(n_28),
.C(n_29),
.Y(n_2117)
);

NOR2xp67_ASAP7_75t_L g2118 ( 
.A(n_1926),
.B(n_29),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1898),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1954),
.B(n_67),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_1956),
.A2(n_69),
.B(n_68),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1919),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_1956),
.A2(n_69),
.B(n_68),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1975),
.B(n_70),
.Y(n_2124)
);

AOI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_1976),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2125)
);

OAI21xp33_ASAP7_75t_SL g2126 ( 
.A1(n_2045),
.A2(n_71),
.B(n_70),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_1900),
.Y(n_2127)
);

AOI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_1998),
.A2(n_1924),
.B1(n_1999),
.B2(n_2041),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1975),
.B(n_72),
.Y(n_2129)
);

INVxp67_ASAP7_75t_L g2130 ( 
.A(n_1989),
.Y(n_2130)
);

AOI21x1_ASAP7_75t_L g2131 ( 
.A1(n_1969),
.A2(n_30),
.B(n_31),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1907),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_2016),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1925),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_2010),
.B(n_2037),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1909),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_2010),
.B(n_73),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1946),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2138)
);

AOI33xp33_ASAP7_75t_L g2139 ( 
.A1(n_2045),
.A2(n_32),
.A3(n_33),
.B1(n_621),
.B2(n_622),
.B3(n_619),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1987),
.B(n_1941),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1913),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1902),
.B(n_73),
.Y(n_2142)
);

BUFx2_ASAP7_75t_L g2143 ( 
.A(n_1994),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_1904),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1987),
.B(n_74),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1928),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2040),
.A2(n_33),
.B1(n_75),
.B2(n_74),
.Y(n_2147)
);

AOI22x1_ASAP7_75t_L g2148 ( 
.A1(n_2020),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1962),
.A2(n_76),
.B(n_79),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_1970),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1960),
.B(n_79),
.Y(n_2151)
);

O2A1O1Ixp33_ASAP7_75t_L g2152 ( 
.A1(n_1969),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1946),
.A2(n_83),
.B1(n_80),
.B2(n_81),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1902),
.B(n_84),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1953),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_2155)
);

AOI21xp5_ASAP7_75t_L g2156 ( 
.A1(n_1962),
.A2(n_85),
.B(n_86),
.Y(n_2156)
);

A2O1A1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_2037),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_2157)
);

BUFx8_ASAP7_75t_SL g2158 ( 
.A(n_1993),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1879),
.B(n_87),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1918),
.Y(n_2160)
);

NOR2x1_ASAP7_75t_SL g2161 ( 
.A(n_1986),
.B(n_88),
.Y(n_2161)
);

INVx5_ASAP7_75t_L g2162 ( 
.A(n_1986),
.Y(n_2162)
);

CKINVDCx11_ASAP7_75t_R g2163 ( 
.A(n_2071),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_L g2164 ( 
.A1(n_2048),
.A2(n_2002),
.B(n_1953),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2144),
.B(n_1904),
.Y(n_2165)
);

AO21x1_ASAP7_75t_L g2166 ( 
.A1(n_2101),
.A2(n_1930),
.B(n_1929),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2054),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2053),
.B(n_1930),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2067),
.B(n_1994),
.Y(n_2169)
);

OA22x2_ASAP7_75t_L g2170 ( 
.A1(n_2125),
.A2(n_2020),
.B1(n_2000),
.B2(n_1934),
.Y(n_2170)
);

NOR2xp67_ASAP7_75t_L g2171 ( 
.A(n_2072),
.B(n_1951),
.Y(n_2171)
);

OAI21x1_ASAP7_75t_L g2172 ( 
.A1(n_2048),
.A2(n_2002),
.B(n_2001),
.Y(n_2172)
);

OAI21x1_ASAP7_75t_L g2173 ( 
.A1(n_2091),
.A2(n_2001),
.B(n_2011),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_L g2174 ( 
.A1(n_2073),
.A2(n_2018),
.B(n_2015),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_2109),
.B(n_2033),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_L g2176 ( 
.A1(n_2073),
.A2(n_2021),
.B(n_1893),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2058),
.B(n_1985),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2065),
.A2(n_2008),
.B(n_2003),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2052),
.A2(n_2019),
.B(n_1982),
.Y(n_2179)
);

AOI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_2065),
.A2(n_2008),
.B(n_2004),
.Y(n_2180)
);

AOI221x1_ASAP7_75t_L g2181 ( 
.A1(n_2149),
.A2(n_1936),
.B1(n_1944),
.B2(n_1942),
.C(n_1939),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2062),
.Y(n_2182)
);

OAI21x1_ASAP7_75t_L g2183 ( 
.A1(n_2088),
.A2(n_1893),
.B(n_1879),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2110),
.B(n_1965),
.Y(n_2184)
);

NAND2x1_ASAP7_75t_L g2185 ( 
.A(n_2099),
.B(n_2111),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2085),
.Y(n_2186)
);

OAI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2092),
.A2(n_2019),
.B(n_1920),
.Y(n_2187)
);

OA21x2_ASAP7_75t_L g2188 ( 
.A1(n_2096),
.A2(n_1920),
.B(n_1908),
.Y(n_2188)
);

OAI21x1_ASAP7_75t_L g2189 ( 
.A1(n_2088),
.A2(n_1922),
.B(n_1908),
.Y(n_2189)
);

NAND2x1p5_ASAP7_75t_L g2190 ( 
.A(n_2162),
.B(n_2008),
.Y(n_2190)
);

NAND3xp33_ASAP7_75t_SL g2191 ( 
.A(n_2139),
.B(n_2017),
.C(n_1971),
.Y(n_2191)
);

O2A1O1Ixp5_ASAP7_75t_L g2192 ( 
.A1(n_2104),
.A2(n_1922),
.B(n_1933),
.C(n_1887),
.Y(n_2192)
);

OAI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2050),
.A2(n_2007),
.B(n_2017),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2061),
.B(n_1996),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_SL g2195 ( 
.A1(n_2108),
.A2(n_2023),
.B(n_2016),
.Y(n_2195)
);

INVxp67_ASAP7_75t_SL g2196 ( 
.A(n_2077),
.Y(n_2196)
);

OAI21x1_ASAP7_75t_L g2197 ( 
.A1(n_2078),
.A2(n_2090),
.B(n_2079),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_2078),
.A2(n_2090),
.B(n_2079),
.Y(n_2198)
);

OAI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_2057),
.A2(n_2007),
.B(n_1963),
.Y(n_2199)
);

INVx1_ASAP7_75t_SL g2200 ( 
.A(n_2150),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2140),
.B(n_1948),
.Y(n_2201)
);

A2O1A1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_2117),
.A2(n_1943),
.B(n_2035),
.C(n_1963),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2064),
.B(n_2089),
.Y(n_2203)
);

OA21x2_ASAP7_75t_L g2204 ( 
.A1(n_2107),
.A2(n_1950),
.B(n_1949),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_L g2205 ( 
.A1(n_2070),
.A2(n_1933),
.B(n_1887),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2086),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2102),
.B(n_1959),
.Y(n_2207)
);

OAI21x1_ASAP7_75t_L g2208 ( 
.A1(n_2105),
.A2(n_2060),
.B(n_2059),
.Y(n_2208)
);

AOI221x1_ASAP7_75t_L g2209 ( 
.A1(n_2149),
.A2(n_1966),
.B1(n_1955),
.B2(n_1961),
.C(n_1974),
.Y(n_2209)
);

OAI21x1_ASAP7_75t_L g2210 ( 
.A1(n_2105),
.A2(n_1991),
.B(n_1978),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_2074),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2162),
.A2(n_1991),
.B(n_1978),
.Y(n_2212)
);

OAI21xp5_ASAP7_75t_L g2213 ( 
.A1(n_2156),
.A2(n_1988),
.B(n_1943),
.Y(n_2213)
);

INVx4_ASAP7_75t_L g2214 ( 
.A(n_2162),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2097),
.B(n_1891),
.Y(n_2215)
);

OAI21x1_ASAP7_75t_L g2216 ( 
.A1(n_2107),
.A2(n_2030),
.B(n_2012),
.Y(n_2216)
);

OAI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2103),
.A2(n_2033),
.B1(n_1945),
.B2(n_1958),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2135),
.B(n_1965),
.Y(n_2218)
);

OAI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2156),
.A2(n_1988),
.B(n_1927),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2098),
.B(n_2033),
.Y(n_2220)
);

AND2x2_ASAP7_75t_SL g2221 ( 
.A(n_2066),
.B(n_1932),
.Y(n_2221)
);

NAND3x1_ASAP7_75t_L g2222 ( 
.A(n_2147),
.B(n_2039),
.C(n_1878),
.Y(n_2222)
);

AND3x4_ASAP7_75t_L g2223 ( 
.A(n_2118),
.B(n_1917),
.C(n_1912),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2132),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_2136),
.B(n_2039),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2094),
.A2(n_2023),
.B(n_1984),
.Y(n_2226)
);

NOR2xp67_ASAP7_75t_L g2227 ( 
.A(n_2076),
.B(n_1903),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2141),
.B(n_1940),
.Y(n_2228)
);

AOI21xp5_ASAP7_75t_L g2229 ( 
.A1(n_2180),
.A2(n_2178),
.B(n_2197),
.Y(n_2229)
);

OAI21x1_ASAP7_75t_L g2230 ( 
.A1(n_2198),
.A2(n_2131),
.B(n_2123),
.Y(n_2230)
);

AOI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_2187),
.A2(n_2069),
.B(n_2080),
.Y(n_2231)
);

BUFx3_ASAP7_75t_L g2232 ( 
.A(n_2163),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2167),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_SL g2234 ( 
.A(n_2171),
.B(n_2055),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2200),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_L g2236 ( 
.A1(n_2170),
.A2(n_2148),
.B1(n_2153),
.B2(n_2121),
.Y(n_2236)
);

OA21x2_ASAP7_75t_L g2237 ( 
.A1(n_2181),
.A2(n_2123),
.B(n_2121),
.Y(n_2237)
);

A2O1A1Ixp33_ASAP7_75t_L g2238 ( 
.A1(n_2208),
.A2(n_2152),
.B(n_2157),
.C(n_2082),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_2215),
.Y(n_2239)
);

AOI221xp5_ASAP7_75t_SL g2240 ( 
.A1(n_2187),
.A2(n_2138),
.B1(n_2115),
.B2(n_2137),
.C(n_2046),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2196),
.B(n_2160),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2219),
.A2(n_2083),
.B(n_2049),
.Y(n_2242)
);

AO31x2_ASAP7_75t_L g2243 ( 
.A1(n_2209),
.A2(n_2111),
.A3(n_2161),
.B(n_2151),
.Y(n_2243)
);

AO21x2_ASAP7_75t_L g2244 ( 
.A1(n_2179),
.A2(n_2159),
.B(n_2120),
.Y(n_2244)
);

OAI21x1_ASAP7_75t_L g2245 ( 
.A1(n_2205),
.A2(n_2100),
.B(n_2124),
.Y(n_2245)
);

NOR2xp67_ASAP7_75t_L g2246 ( 
.A(n_2214),
.B(n_2130),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2182),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_2200),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_2221),
.B(n_2047),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2206),
.Y(n_2250)
);

O2A1O1Ixp33_ASAP7_75t_L g2251 ( 
.A1(n_2202),
.A2(n_2126),
.B(n_2114),
.C(n_2129),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2170),
.A2(n_2093),
.B1(n_2128),
.B2(n_2116),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2213),
.A2(n_2145),
.B1(n_2112),
.B2(n_2106),
.Y(n_2253)
);

OAI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_2213),
.A2(n_2113),
.B1(n_2084),
.B2(n_2143),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2219),
.A2(n_2155),
.B(n_2051),
.Y(n_2255)
);

AO21x1_ASAP7_75t_L g2256 ( 
.A1(n_2203),
.A2(n_2081),
.B(n_2075),
.Y(n_2256)
);

AO31x2_ASAP7_75t_L g2257 ( 
.A1(n_2214),
.A2(n_2095),
.A3(n_2119),
.B(n_2087),
.Y(n_2257)
);

INVx3_ASAP7_75t_L g2258 ( 
.A(n_2225),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_2165),
.Y(n_2259)
);

AOI22xp33_ASAP7_75t_L g2260 ( 
.A1(n_2166),
.A2(n_1927),
.B1(n_2154),
.B2(n_2142),
.Y(n_2260)
);

INVx2_ASAP7_75t_SL g2261 ( 
.A(n_2220),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2199),
.B(n_2226),
.Y(n_2262)
);

AOI21xp33_ASAP7_75t_L g2263 ( 
.A1(n_2204),
.A2(n_2068),
.B(n_2122),
.Y(n_2263)
);

AO31x2_ASAP7_75t_L g2264 ( 
.A1(n_2212),
.A2(n_2134),
.A3(n_2146),
.B(n_2063),
.Y(n_2264)
);

AOI21xp5_ASAP7_75t_L g2265 ( 
.A1(n_2179),
.A2(n_1938),
.B(n_1984),
.Y(n_2265)
);

AOI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2185),
.A2(n_1938),
.B(n_2024),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_2223),
.Y(n_2267)
);

O2A1O1Ixp33_ASAP7_75t_SL g2268 ( 
.A1(n_2169),
.A2(n_2056),
.B(n_1997),
.C(n_1964),
.Y(n_2268)
);

OAI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_2222),
.A2(n_1927),
.B(n_2133),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_2225),
.Y(n_2270)
);

AOI21xp5_ASAP7_75t_L g2271 ( 
.A1(n_2193),
.A2(n_2024),
.B(n_1940),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2190),
.Y(n_2272)
);

AOI21xp33_ASAP7_75t_L g2273 ( 
.A1(n_2244),
.A2(n_2168),
.B(n_2204),
.Y(n_2273)
);

CKINVDCx16_ASAP7_75t_R g2274 ( 
.A(n_2232),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2239),
.B(n_2224),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2236),
.A2(n_2195),
.B1(n_2168),
.B2(n_2199),
.Y(n_2276)
);

OA21x2_ASAP7_75t_L g2277 ( 
.A1(n_2229),
.A2(n_2216),
.B(n_2164),
.Y(n_2277)
);

OAI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2242),
.A2(n_2217),
.B1(n_2177),
.B2(n_2190),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_SL g2279 ( 
.A1(n_2231),
.A2(n_2217),
.B1(n_2218),
.B2(n_2175),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2257),
.Y(n_2280)
);

OAI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2262),
.A2(n_2192),
.B(n_2193),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2230),
.A2(n_2183),
.B(n_2189),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2259),
.B(n_2186),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2233),
.Y(n_2284)
);

OA21x2_ASAP7_75t_L g2285 ( 
.A1(n_2263),
.A2(n_2176),
.B(n_2172),
.Y(n_2285)
);

OAI21xp5_ASAP7_75t_L g2286 ( 
.A1(n_2238),
.A2(n_2210),
.B(n_2227),
.Y(n_2286)
);

NOR2x1_ASAP7_75t_SL g2287 ( 
.A(n_2244),
.B(n_2272),
.Y(n_2287)
);

OA21x2_ASAP7_75t_L g2288 ( 
.A1(n_2245),
.A2(n_2173),
.B(n_2174),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2246),
.B(n_2165),
.Y(n_2289)
);

AO31x2_ASAP7_75t_L g2290 ( 
.A1(n_2256),
.A2(n_2228),
.A3(n_2201),
.B(n_2194),
.Y(n_2290)
);

CKINVDCx16_ASAP7_75t_R g2291 ( 
.A(n_2234),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2247),
.Y(n_2292)
);

OAI21x1_ASAP7_75t_L g2293 ( 
.A1(n_2269),
.A2(n_2188),
.B(n_2228),
.Y(n_2293)
);

OAI21x1_ASAP7_75t_L g2294 ( 
.A1(n_2237),
.A2(n_2188),
.B(n_2201),
.Y(n_2294)
);

AOI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2237),
.A2(n_2191),
.B(n_2177),
.Y(n_2295)
);

CKINVDCx16_ASAP7_75t_R g2296 ( 
.A(n_2267),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2235),
.B(n_2207),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_2272),
.Y(n_2298)
);

CKINVDCx20_ASAP7_75t_R g2299 ( 
.A(n_2274),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2280),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2284),
.Y(n_2301)
);

OA21x2_ASAP7_75t_L g2302 ( 
.A1(n_2280),
.A2(n_2246),
.B(n_2250),
.Y(n_2302)
);

A2O1A1Ixp33_ASAP7_75t_L g2303 ( 
.A1(n_2281),
.A2(n_2286),
.B(n_2295),
.C(n_2276),
.Y(n_2303)
);

OAI21x1_ASAP7_75t_L g2304 ( 
.A1(n_2294),
.A2(n_2258),
.B(n_2249),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2275),
.B(n_2248),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2284),
.Y(n_2306)
);

OAI21x1_ASAP7_75t_L g2307 ( 
.A1(n_2294),
.A2(n_2258),
.B(n_2241),
.Y(n_2307)
);

AO31x2_ASAP7_75t_L g2308 ( 
.A1(n_2287),
.A2(n_2255),
.A3(n_2265),
.B(n_2271),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2299),
.A2(n_2278),
.B1(n_2279),
.B2(n_2254),
.Y(n_2309)
);

AOI22xp33_ASAP7_75t_L g2310 ( 
.A1(n_2305),
.A2(n_2253),
.B1(n_2252),
.B2(n_2267),
.Y(n_2310)
);

BUFx4f_ASAP7_75t_SL g2311 ( 
.A(n_2301),
.Y(n_2311)
);

INVx2_ASAP7_75t_SL g2312 ( 
.A(n_2301),
.Y(n_2312)
);

OAI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2303),
.A2(n_2252),
.B1(n_2291),
.B2(n_2260),
.Y(n_2313)
);

OAI21xp5_ASAP7_75t_SL g2314 ( 
.A1(n_2308),
.A2(n_2251),
.B(n_2267),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2306),
.A2(n_2291),
.B1(n_2296),
.B2(n_2274),
.Y(n_2315)
);

AOI211xp5_ASAP7_75t_L g2316 ( 
.A1(n_2304),
.A2(n_2273),
.B(n_2268),
.C(n_2240),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_2312),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2311),
.Y(n_2318)
);

OA21x2_ASAP7_75t_L g2319 ( 
.A1(n_2314),
.A2(n_2300),
.B(n_2307),
.Y(n_2319)
);

AND2x4_ASAP7_75t_L g2320 ( 
.A(n_2309),
.B(n_2280),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_2316),
.Y(n_2321)
);

BUFx3_ASAP7_75t_L g2322 ( 
.A(n_2315),
.Y(n_2322)
);

INVx2_ASAP7_75t_SL g2323 ( 
.A(n_2313),
.Y(n_2323)
);

AO21x2_ASAP7_75t_L g2324 ( 
.A1(n_2310),
.A2(n_2287),
.B(n_2300),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2312),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2312),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2318),
.B(n_2308),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2318),
.B(n_2308),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2322),
.B(n_2308),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2318),
.B(n_2308),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2318),
.B(n_2308),
.Y(n_2331)
);

HB1xp67_ASAP7_75t_L g2332 ( 
.A(n_2317),
.Y(n_2332)
);

INVx2_ASAP7_75t_SL g2333 ( 
.A(n_2317),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2318),
.B(n_2296),
.Y(n_2334)
);

OR2x2_ASAP7_75t_L g2335 ( 
.A(n_2322),
.B(n_2297),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2317),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2318),
.B(n_2304),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2332),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2334),
.B(n_2322),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2337),
.B(n_2322),
.Y(n_2340)
);

NOR2x1_ASAP7_75t_SL g2341 ( 
.A(n_2333),
.B(n_2323),
.Y(n_2341)
);

INVx3_ASAP7_75t_L g2342 ( 
.A(n_2333),
.Y(n_2342)
);

INVx2_ASAP7_75t_SL g2343 ( 
.A(n_2336),
.Y(n_2343)
);

OR2x2_ASAP7_75t_L g2344 ( 
.A(n_2335),
.B(n_2323),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2327),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2327),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2339),
.B(n_2321),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2339),
.B(n_2322),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2340),
.B(n_2321),
.Y(n_2349)
);

BUFx2_ASAP7_75t_L g2350 ( 
.A(n_2342),
.Y(n_2350)
);

OR2x2_ASAP7_75t_L g2351 ( 
.A(n_2347),
.B(n_2344),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2350),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2348),
.B(n_2340),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_2349),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2353),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2352),
.B(n_2321),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2354),
.B(n_2321),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2351),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2354),
.B(n_2321),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2353),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2355),
.B(n_2338),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2357),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2360),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2356),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2358),
.B(n_2321),
.Y(n_2365)
);

OR2x2_ASAP7_75t_L g2366 ( 
.A(n_2359),
.B(n_2344),
.Y(n_2366)
);

NOR2xp67_ASAP7_75t_L g2367 ( 
.A(n_2358),
.B(n_2342),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2355),
.B(n_2321),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2355),
.B(n_2321),
.Y(n_2369)
);

NAND2x1_ASAP7_75t_L g2370 ( 
.A(n_2357),
.B(n_2342),
.Y(n_2370)
);

NAND2x1p5_ASAP7_75t_L g2371 ( 
.A(n_2370),
.B(n_2342),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2361),
.B(n_2338),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_2367),
.Y(n_2373)
);

OR2x2_ASAP7_75t_L g2374 ( 
.A(n_2365),
.B(n_2343),
.Y(n_2374)
);

INVxp67_ASAP7_75t_L g2375 ( 
.A(n_2366),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2362),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2363),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2368),
.B(n_2341),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2369),
.B(n_2341),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2364),
.B(n_2343),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2367),
.B(n_2323),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2361),
.B(n_2322),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2367),
.B(n_2323),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2372),
.B(n_2323),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2373),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2383),
.Y(n_2386)
);

INVxp67_ASAP7_75t_SL g2387 ( 
.A(n_2371),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2383),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2382),
.B(n_2337),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2381),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2380),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2374),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2376),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2378),
.B(n_2346),
.Y(n_2394)
);

NOR2x1_ASAP7_75t_L g2395 ( 
.A(n_2376),
.B(n_2346),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2379),
.B(n_2320),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2377),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2375),
.Y(n_2398)
);

NAND2x1p5_ASAP7_75t_L g2399 ( 
.A(n_2384),
.B(n_2127),
.Y(n_2399)
);

INVx2_ASAP7_75t_SL g2400 ( 
.A(n_2384),
.Y(n_2400)
);

INVx1_ASAP7_75t_SL g2401 ( 
.A(n_2389),
.Y(n_2401)
);

O2A1O1Ixp33_ASAP7_75t_SL g2402 ( 
.A1(n_2396),
.A2(n_2329),
.B(n_2345),
.C(n_2326),
.Y(n_2402)
);

OAI32xp33_ASAP7_75t_L g2403 ( 
.A1(n_2394),
.A2(n_2345),
.A3(n_2331),
.B1(n_2330),
.B2(n_2328),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2387),
.B(n_2320),
.Y(n_2404)
);

OAI222xp33_ASAP7_75t_L g2405 ( 
.A1(n_2385),
.A2(n_2330),
.B1(n_2331),
.B2(n_2328),
.C1(n_2325),
.C2(n_2326),
.Y(n_2405)
);

NAND3x2_ASAP7_75t_L g2406 ( 
.A(n_2398),
.B(n_2320),
.C(n_2325),
.Y(n_2406)
);

OAI32xp33_ASAP7_75t_L g2407 ( 
.A1(n_2397),
.A2(n_2326),
.A3(n_2325),
.B1(n_2324),
.B2(n_2300),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2391),
.B(n_2158),
.Y(n_2408)
);

AOI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2392),
.A2(n_2390),
.B1(n_2388),
.B2(n_2386),
.Y(n_2409)
);

INVx1_ASAP7_75t_SL g2410 ( 
.A(n_2395),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_2393),
.B(n_2325),
.Y(n_2411)
);

NAND3xp33_ASAP7_75t_L g2412 ( 
.A(n_2387),
.B(n_2326),
.C(n_2319),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2400),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2404),
.Y(n_2414)
);

A2O1A1Ixp33_ASAP7_75t_L g2415 ( 
.A1(n_2408),
.A2(n_2320),
.B(n_2324),
.C(n_2307),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2401),
.B(n_2320),
.Y(n_2416)
);

OAI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2409),
.A2(n_2320),
.B1(n_2319),
.B2(n_2298),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2402),
.Y(n_2418)
);

OAI31xp33_ASAP7_75t_L g2419 ( 
.A1(n_2410),
.A2(n_2320),
.A3(n_2324),
.B(n_2319),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2399),
.B(n_2320),
.Y(n_2420)
);

OAI22xp5_ASAP7_75t_SL g2421 ( 
.A1(n_2411),
.A2(n_2319),
.B1(n_2324),
.B2(n_1980),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2406),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2403),
.B(n_2324),
.Y(n_2423)
);

OAI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2412),
.A2(n_2319),
.B1(n_2298),
.B2(n_2306),
.Y(n_2424)
);

AOI221xp5_ASAP7_75t_L g2425 ( 
.A1(n_2405),
.A2(n_2324),
.B1(n_2319),
.B2(n_1947),
.C(n_2298),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2407),
.B(n_2298),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2408),
.B(n_2324),
.Y(n_2427)
);

OR4x1_ASAP7_75t_L g2428 ( 
.A(n_2400),
.B(n_2324),
.C(n_1957),
.D(n_2319),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2400),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2400),
.A2(n_2319),
.B1(n_1921),
.B2(n_2036),
.Y(n_2430)
);

AOI332xp33_ASAP7_75t_L g2431 ( 
.A1(n_2409),
.A2(n_2319),
.A3(n_94),
.B1(n_91),
.B2(n_95),
.B3(n_93),
.C1(n_89),
.C2(n_90),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2400),
.B(n_2036),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2400),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2404),
.A2(n_2298),
.B1(n_2289),
.B2(n_2302),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_2432),
.A2(n_2266),
.B(n_1947),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2413),
.B(n_2429),
.Y(n_2436)
);

AOI21xp33_ASAP7_75t_L g2437 ( 
.A1(n_2433),
.A2(n_90),
.B(n_91),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2420),
.B(n_92),
.Y(n_2438)
);

OAI211xp5_ASAP7_75t_SL g2439 ( 
.A1(n_2414),
.A2(n_2422),
.B(n_2416),
.C(n_2418),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2427),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2423),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2426),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2424),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2419),
.B(n_92),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2417),
.Y(n_2445)
);

INVx2_ASAP7_75t_SL g2446 ( 
.A(n_2434),
.Y(n_2446)
);

OAI322xp33_ASAP7_75t_L g2447 ( 
.A1(n_2421),
.A2(n_2430),
.A3(n_2431),
.B1(n_2428),
.B2(n_2415),
.C1(n_2425),
.C2(n_2298),
.Y(n_2447)
);

NOR2x1_ASAP7_75t_L g2448 ( 
.A(n_2430),
.B(n_93),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2413),
.B(n_96),
.Y(n_2449)
);

XNOR2x2_ASAP7_75t_L g2450 ( 
.A(n_2418),
.B(n_96),
.Y(n_2450)
);

AO22x2_ASAP7_75t_L g2451 ( 
.A1(n_2418),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2451)
);

OR2x2_ASAP7_75t_L g2452 ( 
.A(n_2416),
.B(n_2243),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2419),
.B(n_1921),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2419),
.B(n_1921),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2416),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2416),
.Y(n_2456)
);

HB1xp67_ASAP7_75t_L g2457 ( 
.A(n_2416),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2416),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2429),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2416),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2429),
.B(n_2275),
.Y(n_2461)
);

NAND3xp33_ASAP7_75t_L g2462 ( 
.A(n_2413),
.B(n_100),
.C(n_101),
.Y(n_2462)
);

AOI221xp5_ASAP7_75t_L g2463 ( 
.A1(n_2422),
.A2(n_2240),
.B1(n_2289),
.B2(n_103),
.C(n_100),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2416),
.Y(n_2464)
);

INVxp67_ASAP7_75t_SL g2465 ( 
.A(n_2416),
.Y(n_2465)
);

AOI31xp33_ASAP7_75t_L g2466 ( 
.A1(n_2413),
.A2(n_110),
.A3(n_118),
.B(n_102),
.Y(n_2466)
);

NOR3xp33_ASAP7_75t_L g2467 ( 
.A(n_2413),
.B(n_110),
.C(n_102),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2416),
.Y(n_2468)
);

OA21x2_ASAP7_75t_L g2469 ( 
.A1(n_2418),
.A2(n_103),
.B(n_104),
.Y(n_2469)
);

INVxp67_ASAP7_75t_L g2470 ( 
.A(n_2432),
.Y(n_2470)
);

OAI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_2416),
.A2(n_2293),
.B(n_2289),
.Y(n_2471)
);

OAI21xp33_ASAP7_75t_L g2472 ( 
.A1(n_2436),
.A2(n_2014),
.B(n_2005),
.Y(n_2472)
);

OAI21xp33_ASAP7_75t_L g2473 ( 
.A1(n_2459),
.A2(n_2031),
.B(n_2028),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_SL g2474 ( 
.A1(n_2465),
.A2(n_2302),
.B1(n_2289),
.B2(n_2272),
.Y(n_2474)
);

OAI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2462),
.A2(n_2302),
.B1(n_2292),
.B2(n_2261),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2466),
.B(n_105),
.Y(n_2476)
);

OAI21xp33_ASAP7_75t_L g2477 ( 
.A1(n_2461),
.A2(n_2292),
.B(n_2283),
.Y(n_2477)
);

AOI222xp33_ASAP7_75t_L g2478 ( 
.A1(n_2442),
.A2(n_106),
.B1(n_108),
.B2(n_104),
.C1(n_105),
.C2(n_107),
.Y(n_2478)
);

AOI221xp5_ASAP7_75t_L g2479 ( 
.A1(n_2447),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.C(n_109),
.Y(n_2479)
);

OAI22xp33_ASAP7_75t_L g2480 ( 
.A1(n_2449),
.A2(n_2302),
.B1(n_2270),
.B2(n_2194),
.Y(n_2480)
);

NOR4xp25_ASAP7_75t_L g2481 ( 
.A(n_2439),
.B(n_112),
.C(n_109),
.D(n_111),
.Y(n_2481)
);

OAI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2455),
.A2(n_2458),
.B1(n_2460),
.B2(n_2456),
.Y(n_2482)
);

NOR2xp67_ASAP7_75t_L g2483 ( 
.A(n_2457),
.B(n_112),
.Y(n_2483)
);

O2A1O1Ixp33_ASAP7_75t_SL g2484 ( 
.A1(n_2453),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2451),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2464),
.A2(n_2283),
.B1(n_2277),
.B2(n_2293),
.Y(n_2486)
);

AOI221xp5_ASAP7_75t_L g2487 ( 
.A1(n_2451),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.C(n_117),
.Y(n_2487)
);

OAI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_2468),
.A2(n_2270),
.B1(n_2277),
.B2(n_2285),
.Y(n_2488)
);

NAND2xp33_ASAP7_75t_SL g2489 ( 
.A(n_2438),
.B(n_116),
.Y(n_2489)
);

AOI221xp5_ASAP7_75t_L g2490 ( 
.A1(n_2443),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.C(n_121),
.Y(n_2490)
);

OAI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2470),
.A2(n_2282),
.B(n_119),
.Y(n_2491)
);

OA21x2_ASAP7_75t_L g2492 ( 
.A1(n_2441),
.A2(n_120),
.B(n_121),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_2463),
.B(n_2270),
.Y(n_2493)
);

XNOR2xp5_ASAP7_75t_L g2494 ( 
.A(n_2450),
.B(n_122),
.Y(n_2494)
);

OAI221xp5_ASAP7_75t_SL g2495 ( 
.A1(n_2452),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.C(n_125),
.Y(n_2495)
);

AOI21xp5_ASAP7_75t_L g2496 ( 
.A1(n_2454),
.A2(n_123),
.B(n_126),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2469),
.Y(n_2497)
);

AO21x1_ASAP7_75t_L g2498 ( 
.A1(n_2444),
.A2(n_126),
.B(n_127),
.Y(n_2498)
);

AOI221xp5_ASAP7_75t_SL g2499 ( 
.A1(n_2445),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2446),
.A2(n_2277),
.B1(n_2285),
.B2(n_2288),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_2437),
.B(n_128),
.Y(n_2501)
);

AOI211xp5_ASAP7_75t_SL g2502 ( 
.A1(n_2440),
.A2(n_133),
.B(n_129),
.C(n_132),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2448),
.A2(n_132),
.B(n_133),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2467),
.B(n_135),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2469),
.Y(n_2505)
);

O2A1O1Ixp5_ASAP7_75t_L g2506 ( 
.A1(n_2471),
.A2(n_137),
.B(n_134),
.C(n_136),
.Y(n_2506)
);

OAI32xp33_ASAP7_75t_L g2507 ( 
.A1(n_2435),
.A2(n_137),
.A3(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2451),
.Y(n_2508)
);

AOI221xp5_ASAP7_75t_L g2509 ( 
.A1(n_2447),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.C(n_141),
.Y(n_2509)
);

OAI211xp5_ASAP7_75t_SL g2510 ( 
.A1(n_2479),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_2510)
);

AOI221x1_ASAP7_75t_L g2511 ( 
.A1(n_2485),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.C(n_145),
.Y(n_2511)
);

OAI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2476),
.A2(n_2277),
.B1(n_2285),
.B2(n_2288),
.Y(n_2512)
);

AOI221xp5_ASAP7_75t_L g2513 ( 
.A1(n_2481),
.A2(n_145),
.B1(n_147),
.B2(n_143),
.C(n_146),
.Y(n_2513)
);

NOR2xp33_ASAP7_75t_L g2514 ( 
.A(n_2505),
.B(n_142),
.Y(n_2514)
);

NOR3xp33_ASAP7_75t_L g2515 ( 
.A(n_2482),
.B(n_148),
.C(n_147),
.Y(n_2515)
);

AOI221xp5_ASAP7_75t_L g2516 ( 
.A1(n_2484),
.A2(n_149),
.B1(n_151),
.B2(n_148),
.C(n_150),
.Y(n_2516)
);

OAI221xp5_ASAP7_75t_SL g2517 ( 
.A1(n_2509),
.A2(n_152),
.B1(n_146),
.B2(n_149),
.C(n_153),
.Y(n_2517)
);

AOI222xp33_ASAP7_75t_L g2518 ( 
.A1(n_2508),
.A2(n_155),
.B1(n_157),
.B2(n_153),
.C1(n_154),
.C2(n_156),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2501),
.A2(n_2026),
.B1(n_2285),
.B2(n_1927),
.Y(n_2519)
);

INVxp67_ASAP7_75t_L g2520 ( 
.A(n_2483),
.Y(n_2520)
);

AOI221xp5_ASAP7_75t_L g2521 ( 
.A1(n_2507),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.C(n_158),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2502),
.B(n_2290),
.Y(n_2522)
);

NAND3xp33_ASAP7_75t_SL g2523 ( 
.A(n_2503),
.B(n_158),
.C(n_159),
.Y(n_2523)
);

OAI32xp33_ASAP7_75t_L g2524 ( 
.A1(n_2504),
.A2(n_161),
.A3(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2494),
.A2(n_2288),
.B1(n_2211),
.B2(n_2184),
.Y(n_2525)
);

NOR2x1_ASAP7_75t_L g2526 ( 
.A(n_2497),
.B(n_160),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2492),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_R g2528 ( 
.A(n_2489),
.B(n_161),
.Y(n_2528)
);

NOR3xp33_ASAP7_75t_L g2529 ( 
.A(n_2495),
.B(n_162),
.C(n_163),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2492),
.Y(n_2530)
);

NAND4xp25_ASAP7_75t_L g2531 ( 
.A(n_2506),
.B(n_165),
.C(n_163),
.D(n_164),
.Y(n_2531)
);

OR2x2_ASAP7_75t_L g2532 ( 
.A(n_2493),
.B(n_165),
.Y(n_2532)
);

OAI221xp5_ASAP7_75t_L g2533 ( 
.A1(n_2499),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.C(n_169),
.Y(n_2533)
);

O2A1O1Ixp33_ASAP7_75t_SL g2534 ( 
.A1(n_2487),
.A2(n_170),
.B(n_166),
.C(n_168),
.Y(n_2534)
);

AOI211xp5_ASAP7_75t_SL g2535 ( 
.A1(n_2496),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2535)
);

NOR3xp33_ASAP7_75t_L g2536 ( 
.A(n_2490),
.B(n_171),
.C(n_173),
.Y(n_2536)
);

INVxp67_ASAP7_75t_L g2537 ( 
.A(n_2478),
.Y(n_2537)
);

O2A1O1Ixp5_ASAP7_75t_L g2538 ( 
.A1(n_2498),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_2538)
);

OAI31xp33_ASAP7_75t_L g2539 ( 
.A1(n_2475),
.A2(n_177),
.A3(n_174),
.B(n_176),
.Y(n_2539)
);

NAND2x1p5_ASAP7_75t_L g2540 ( 
.A(n_2472),
.B(n_2473),
.Y(n_2540)
);

INVx2_ASAP7_75t_SL g2541 ( 
.A(n_2491),
.Y(n_2541)
);

OAI322xp33_ASAP7_75t_L g2542 ( 
.A1(n_2480),
.A2(n_2500),
.A3(n_2488),
.B1(n_2486),
.B2(n_2474),
.C1(n_2477),
.C2(n_179),
.Y(n_2542)
);

AOI211xp5_ASAP7_75t_L g2543 ( 
.A1(n_2507),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2543)
);

NOR3x1_ASAP7_75t_L g2544 ( 
.A(n_2476),
.B(n_180),
.C(n_181),
.Y(n_2544)
);

AOI211xp5_ASAP7_75t_SL g2545 ( 
.A1(n_2482),
.A2(n_183),
.B(n_180),
.C(n_182),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2505),
.Y(n_2546)
);

O2A1O1Ixp33_ASAP7_75t_L g2547 ( 
.A1(n_2505),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2483),
.B(n_184),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2497),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_2481),
.B(n_186),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_SL g2551 ( 
.A(n_2483),
.B(n_186),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2483),
.B(n_187),
.Y(n_2552)
);

AOI221xp5_ASAP7_75t_L g2553 ( 
.A1(n_2481),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2489),
.A2(n_188),
.B(n_189),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2483),
.B(n_190),
.Y(n_2555)
);

OAI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2476),
.A2(n_2288),
.B1(n_2211),
.B2(n_193),
.Y(n_2556)
);

OAI21xp33_ASAP7_75t_L g2557 ( 
.A1(n_2481),
.A2(n_2282),
.B(n_191),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_L g2558 ( 
.A(n_2476),
.B(n_192),
.Y(n_2558)
);

NOR4xp25_ASAP7_75t_L g2559 ( 
.A(n_2485),
.B(n_196),
.C(n_194),
.D(n_195),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2483),
.B(n_194),
.Y(n_2560)
);

A2O1A1Ixp33_ASAP7_75t_L g2561 ( 
.A1(n_2483),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2505),
.Y(n_2562)
);

OAI21xp5_ASAP7_75t_SL g2563 ( 
.A1(n_2494),
.A2(n_197),
.B(n_198),
.Y(n_2563)
);

O2A1O1Ixp5_ASAP7_75t_L g2564 ( 
.A1(n_2497),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_2564)
);

NAND3xp33_ASAP7_75t_L g2565 ( 
.A(n_2479),
.B(n_199),
.C(n_201),
.Y(n_2565)
);

O2A1O1Ixp5_ASAP7_75t_L g2566 ( 
.A1(n_2497),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_2566)
);

AOI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2489),
.A2(n_202),
.B(n_203),
.Y(n_2567)
);

OAI21xp33_ASAP7_75t_L g2568 ( 
.A1(n_2481),
.A2(n_204),
.B(n_205),
.Y(n_2568)
);

AOI21xp33_ASAP7_75t_SL g2569 ( 
.A1(n_2494),
.A2(n_205),
.B(n_206),
.Y(n_2569)
);

NAND4xp25_ASAP7_75t_SL g2570 ( 
.A(n_2479),
.B(n_209),
.C(n_207),
.D(n_208),
.Y(n_2570)
);

AOI221xp5_ASAP7_75t_L g2571 ( 
.A1(n_2481),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.C(n_212),
.Y(n_2571)
);

NOR3xp33_ASAP7_75t_L g2572 ( 
.A(n_2482),
.B(n_211),
.C(n_212),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2489),
.A2(n_213),
.B(n_214),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2514),
.B(n_213),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2527),
.Y(n_2575)
);

OAI211xp5_ASAP7_75t_SL g2576 ( 
.A1(n_2537),
.A2(n_218),
.B(n_215),
.C(n_216),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2530),
.Y(n_2577)
);

OAI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_2517),
.A2(n_2565),
.B1(n_2533),
.B2(n_2520),
.Y(n_2578)
);

NAND3xp33_ASAP7_75t_L g2579 ( 
.A(n_2545),
.B(n_215),
.C(n_216),
.Y(n_2579)
);

AOI221xp5_ASAP7_75t_L g2580 ( 
.A1(n_2569),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.C(n_221),
.Y(n_2580)
);

OAI21xp33_ASAP7_75t_SL g2581 ( 
.A1(n_2550),
.A2(n_219),
.B(n_220),
.Y(n_2581)
);

OAI21xp33_ASAP7_75t_L g2582 ( 
.A1(n_2568),
.A2(n_221),
.B(n_222),
.Y(n_2582)
);

NAND4xp25_ASAP7_75t_L g2583 ( 
.A(n_2543),
.B(n_224),
.C(n_222),
.D(n_223),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2559),
.B(n_2290),
.Y(n_2584)
);

AND3x1_ASAP7_75t_L g2585 ( 
.A(n_2551),
.B(n_223),
.C(n_225),
.Y(n_2585)
);

OAI21xp5_ASAP7_75t_SL g2586 ( 
.A1(n_2563),
.A2(n_2535),
.B(n_2510),
.Y(n_2586)
);

NAND3xp33_ASAP7_75t_L g2587 ( 
.A(n_2515),
.B(n_225),
.C(n_227),
.Y(n_2587)
);

AOI211xp5_ASAP7_75t_SL g2588 ( 
.A1(n_2558),
.A2(n_229),
.B(n_227),
.C(n_228),
.Y(n_2588)
);

AOI211xp5_ASAP7_75t_SL g2589 ( 
.A1(n_2534),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2589)
);

A2O1A1Ixp33_ASAP7_75t_L g2590 ( 
.A1(n_2538),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_2590)
);

NAND3xp33_ASAP7_75t_L g2591 ( 
.A(n_2572),
.B(n_231),
.C(n_233),
.Y(n_2591)
);

AOI211xp5_ASAP7_75t_L g2592 ( 
.A1(n_2570),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_2592)
);

OAI221xp5_ASAP7_75t_L g2593 ( 
.A1(n_2539),
.A2(n_237),
.B1(n_234),
.B2(n_236),
.C(n_238),
.Y(n_2593)
);

OAI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2554),
.A2(n_2573),
.B(n_2567),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2526),
.Y(n_2595)
);

NOR3xp33_ASAP7_75t_L g2596 ( 
.A(n_2548),
.B(n_236),
.C(n_237),
.Y(n_2596)
);

AOI21xp33_ASAP7_75t_SL g2597 ( 
.A1(n_2547),
.A2(n_238),
.B(n_239),
.Y(n_2597)
);

NAND3xp33_ASAP7_75t_L g2598 ( 
.A(n_2521),
.B(n_241),
.C(n_242),
.Y(n_2598)
);

OAI221xp5_ASAP7_75t_L g2599 ( 
.A1(n_2557),
.A2(n_244),
.B1(n_241),
.B2(n_243),
.C(n_245),
.Y(n_2599)
);

OAI211xp5_ASAP7_75t_SL g2600 ( 
.A1(n_2546),
.A2(n_246),
.B(n_243),
.C(n_245),
.Y(n_2600)
);

O2A1O1Ixp5_ASAP7_75t_SL g2601 ( 
.A1(n_2562),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_2601)
);

NAND4xp25_ASAP7_75t_L g2602 ( 
.A(n_2529),
.B(n_2513),
.C(n_2571),
.D(n_2553),
.Y(n_2602)
);

AOI221x1_ASAP7_75t_L g2603 ( 
.A1(n_2549),
.A2(n_2560),
.B1(n_2555),
.B2(n_2552),
.C(n_2536),
.Y(n_2603)
);

NOR3xp33_ASAP7_75t_L g2604 ( 
.A(n_2523),
.B(n_247),
.C(n_248),
.Y(n_2604)
);

AOI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2561),
.A2(n_249),
.B(n_250),
.Y(n_2605)
);

NOR3xp33_ASAP7_75t_L g2606 ( 
.A(n_2532),
.B(n_249),
.C(n_251),
.Y(n_2606)
);

O2A1O1Ixp33_ASAP7_75t_L g2607 ( 
.A1(n_2564),
.A2(n_2566),
.B(n_2524),
.C(n_2541),
.Y(n_2607)
);

OAI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2519),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_2608)
);

A2O1A1Ixp33_ASAP7_75t_L g2609 ( 
.A1(n_2516),
.A2(n_2531),
.B(n_2556),
.C(n_2522),
.Y(n_2609)
);

OAI211xp5_ASAP7_75t_SL g2610 ( 
.A1(n_2518),
.A2(n_255),
.B(n_252),
.C(n_254),
.Y(n_2610)
);

NAND3xp33_ASAP7_75t_L g2611 ( 
.A(n_2511),
.B(n_254),
.C(n_255),
.Y(n_2611)
);

OAI221xp5_ASAP7_75t_L g2612 ( 
.A1(n_2540),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.C(n_259),
.Y(n_2612)
);

AOI222xp33_ASAP7_75t_L g2613 ( 
.A1(n_2525),
.A2(n_258),
.B1(n_260),
.B2(n_256),
.C1(n_257),
.C2(n_259),
.Y(n_2613)
);

OAI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2540),
.A2(n_260),
.B(n_261),
.Y(n_2614)
);

AOI21xp33_ASAP7_75t_L g2615 ( 
.A1(n_2528),
.A2(n_261),
.B(n_262),
.Y(n_2615)
);

OAI21xp5_ASAP7_75t_L g2616 ( 
.A1(n_2544),
.A2(n_2512),
.B(n_2542),
.Y(n_2616)
);

O2A1O1Ixp33_ASAP7_75t_L g2617 ( 
.A1(n_2527),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_2617)
);

AOI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2550),
.A2(n_263),
.B(n_264),
.Y(n_2618)
);

OAI21xp5_ASAP7_75t_SL g2619 ( 
.A1(n_2563),
.A2(n_266),
.B(n_267),
.Y(n_2619)
);

AOI221xp5_ASAP7_75t_L g2620 ( 
.A1(n_2569),
.A2(n_269),
.B1(n_266),
.B2(n_268),
.C(n_270),
.Y(n_2620)
);

O2A1O1Ixp33_ASAP7_75t_L g2621 ( 
.A1(n_2527),
.A2(n_271),
.B(n_268),
.C(n_270),
.Y(n_2621)
);

O2A1O1Ixp33_ASAP7_75t_L g2622 ( 
.A1(n_2527),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_2622)
);

AOI22xp5_ASAP7_75t_L g2623 ( 
.A1(n_2570),
.A2(n_2026),
.B1(n_1927),
.B2(n_274),
.Y(n_2623)
);

AOI32xp33_ASAP7_75t_L g2624 ( 
.A1(n_2510),
.A2(n_275),
.A3(n_272),
.B1(n_273),
.B2(n_276),
.Y(n_2624)
);

OAI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2539),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.C(n_278),
.Y(n_2625)
);

AOI221xp5_ASAP7_75t_L g2626 ( 
.A1(n_2569),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.C(n_280),
.Y(n_2626)
);

OAI211xp5_ASAP7_75t_SL g2627 ( 
.A1(n_2537),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2627)
);

AOI221xp5_ASAP7_75t_L g2628 ( 
.A1(n_2569),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.C(n_284),
.Y(n_2628)
);

AOI221xp5_ASAP7_75t_SL g2629 ( 
.A1(n_2542),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.C(n_285),
.Y(n_2629)
);

NAND5xp2_ASAP7_75t_L g2630 ( 
.A(n_2539),
.B(n_288),
.C(n_285),
.D(n_286),
.E(n_291),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2527),
.Y(n_2631)
);

OA21x2_ASAP7_75t_L g2632 ( 
.A1(n_2527),
.A2(n_286),
.B(n_288),
.Y(n_2632)
);

OAI311xp33_ASAP7_75t_L g2633 ( 
.A1(n_2557),
.A2(n_294),
.A3(n_292),
.B1(n_293),
.C1(n_295),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2514),
.B(n_293),
.Y(n_2634)
);

NAND4xp25_ASAP7_75t_SL g2635 ( 
.A(n_2513),
.B(n_297),
.C(n_295),
.D(n_296),
.Y(n_2635)
);

AOI221xp5_ASAP7_75t_L g2636 ( 
.A1(n_2569),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.C(n_299),
.Y(n_2636)
);

OAI211xp5_ASAP7_75t_L g2637 ( 
.A1(n_2563),
.A2(n_301),
.B(n_298),
.C(n_300),
.Y(n_2637)
);

OAI211xp5_ASAP7_75t_L g2638 ( 
.A1(n_2563),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_2638)
);

OR3x1_ASAP7_75t_L g2639 ( 
.A(n_2570),
.B(n_303),
.C(n_304),
.Y(n_2639)
);

NAND3xp33_ASAP7_75t_L g2640 ( 
.A(n_2545),
.B(n_303),
.C(n_304),
.Y(n_2640)
);

AOI221xp5_ASAP7_75t_L g2641 ( 
.A1(n_2569),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.C(n_308),
.Y(n_2641)
);

OAI221xp5_ASAP7_75t_L g2642 ( 
.A1(n_2539),
.A2(n_309),
.B1(n_306),
.B2(n_307),
.C(n_310),
.Y(n_2642)
);

OAI211xp5_ASAP7_75t_L g2643 ( 
.A1(n_2563),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_2643)
);

OAI211xp5_ASAP7_75t_L g2644 ( 
.A1(n_2563),
.A2(n_313),
.B(n_311),
.C(n_312),
.Y(n_2644)
);

NAND5xp2_ASAP7_75t_L g2645 ( 
.A(n_2539),
.B(n_315),
.C(n_312),
.D(n_314),
.E(n_316),
.Y(n_2645)
);

OAI221xp5_ASAP7_75t_L g2646 ( 
.A1(n_2539),
.A2(n_318),
.B1(n_314),
.B2(n_317),
.C(n_319),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2527),
.Y(n_2647)
);

AO221x1_ASAP7_75t_L g2648 ( 
.A1(n_2569),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.C(n_321),
.Y(n_2648)
);

NOR2xp67_ASAP7_75t_L g2649 ( 
.A(n_2527),
.B(n_321),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_SL g2650 ( 
.A(n_2559),
.B(n_322),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2576),
.B(n_323),
.Y(n_2651)
);

AOI21xp5_ASAP7_75t_L g2652 ( 
.A1(n_2650),
.A2(n_323),
.B(n_324),
.Y(n_2652)
);

AOI311xp33_ASAP7_75t_L g2653 ( 
.A1(n_2578),
.A2(n_326),
.A3(n_324),
.B(n_325),
.C(n_327),
.Y(n_2653)
);

NOR4xp25_ASAP7_75t_L g2654 ( 
.A(n_2607),
.B(n_328),
.C(n_325),
.D(n_326),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2649),
.B(n_328),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2627),
.B(n_329),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2630),
.B(n_329),
.Y(n_2657)
);

NOR3xp33_ASAP7_75t_L g2658 ( 
.A(n_2615),
.B(n_330),
.C(n_331),
.Y(n_2658)
);

NAND3xp33_ASAP7_75t_L g2659 ( 
.A(n_2606),
.B(n_330),
.C(n_331),
.Y(n_2659)
);

OAI211xp5_ASAP7_75t_SL g2660 ( 
.A1(n_2581),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_2660)
);

NAND4xp25_ASAP7_75t_L g2661 ( 
.A(n_2592),
.B(n_334),
.C(n_332),
.D(n_333),
.Y(n_2661)
);

NAND4xp25_ASAP7_75t_L g2662 ( 
.A(n_2589),
.B(n_337),
.C(n_335),
.D(n_336),
.Y(n_2662)
);

NOR4xp75_ASAP7_75t_L g2663 ( 
.A(n_2616),
.B(n_338),
.C(n_335),
.D(n_337),
.Y(n_2663)
);

AOI222xp33_ASAP7_75t_L g2664 ( 
.A1(n_2575),
.A2(n_340),
.B1(n_342),
.B2(n_338),
.C1(n_339),
.C2(n_341),
.Y(n_2664)
);

NAND4xp75_ASAP7_75t_L g2665 ( 
.A(n_2603),
.B(n_342),
.C(n_339),
.D(n_341),
.Y(n_2665)
);

OAI211xp5_ASAP7_75t_L g2666 ( 
.A1(n_2619),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2588),
.B(n_343),
.Y(n_2667)
);

AOI21xp5_ASAP7_75t_L g2668 ( 
.A1(n_2577),
.A2(n_344),
.B(n_345),
.Y(n_2668)
);

NOR3xp33_ASAP7_75t_L g2669 ( 
.A(n_2647),
.B(n_346),
.C(n_347),
.Y(n_2669)
);

OAI211xp5_ASAP7_75t_SL g2670 ( 
.A1(n_2582),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_2670)
);

NAND3xp33_ASAP7_75t_L g2671 ( 
.A(n_2596),
.B(n_349),
.C(n_350),
.Y(n_2671)
);

AOI221xp5_ASAP7_75t_L g2672 ( 
.A1(n_2597),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.C(n_352),
.Y(n_2672)
);

NOR3xp33_ASAP7_75t_L g2673 ( 
.A(n_2647),
.B(n_2634),
.C(n_2574),
.Y(n_2673)
);

NOR3xp33_ASAP7_75t_L g2674 ( 
.A(n_2631),
.B(n_351),
.C(n_353),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2648),
.B(n_2590),
.Y(n_2675)
);

AOI211xp5_ASAP7_75t_L g2676 ( 
.A1(n_2599),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_2676)
);

AO22x2_ASAP7_75t_L g2677 ( 
.A1(n_2595),
.A2(n_358),
.B1(n_355),
.B2(n_357),
.Y(n_2677)
);

AOI211xp5_ASAP7_75t_L g2678 ( 
.A1(n_2593),
.A2(n_360),
.B(n_358),
.C(n_359),
.Y(n_2678)
);

NAND4xp75_ASAP7_75t_L g2679 ( 
.A(n_2629),
.B(n_362),
.C(n_359),
.D(n_360),
.Y(n_2679)
);

OAI221xp5_ASAP7_75t_L g2680 ( 
.A1(n_2624),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.C(n_365),
.Y(n_2680)
);

O2A1O1Ixp5_ASAP7_75t_SL g2681 ( 
.A1(n_2637),
.A2(n_366),
.B(n_363),
.C(n_364),
.Y(n_2681)
);

NOR4xp25_ASAP7_75t_L g2682 ( 
.A(n_2633),
.B(n_368),
.C(n_366),
.D(n_367),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2580),
.B(n_367),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2620),
.B(n_2626),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2585),
.B(n_368),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2645),
.B(n_369),
.Y(n_2686)
);

NOR3xp33_ASAP7_75t_L g2687 ( 
.A(n_2602),
.B(n_369),
.C(n_370),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2628),
.B(n_370),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2636),
.B(n_371),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2641),
.B(n_372),
.Y(n_2690)
);

NAND4xp75_ASAP7_75t_L g2691 ( 
.A(n_2618),
.B(n_375),
.C(n_373),
.D(n_374),
.Y(n_2691)
);

NOR3xp33_ASAP7_75t_L g2692 ( 
.A(n_2638),
.B(n_2644),
.C(n_2643),
.Y(n_2692)
);

XOR2x2_ASAP7_75t_L g2693 ( 
.A(n_2611),
.B(n_374),
.Y(n_2693)
);

NOR4xp25_ASAP7_75t_L g2694 ( 
.A(n_2609),
.B(n_378),
.C(n_376),
.D(n_377),
.Y(n_2694)
);

INVxp67_ASAP7_75t_L g2695 ( 
.A(n_2632),
.Y(n_2695)
);

NAND3xp33_ASAP7_75t_L g2696 ( 
.A(n_2604),
.B(n_377),
.C(n_378),
.Y(n_2696)
);

NOR4xp25_ASAP7_75t_L g2697 ( 
.A(n_2610),
.B(n_381),
.C(n_379),
.D(n_380),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2594),
.B(n_2290),
.Y(n_2698)
);

NOR3xp33_ASAP7_75t_L g2699 ( 
.A(n_2625),
.B(n_379),
.C(n_380),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2614),
.B(n_381),
.Y(n_2700)
);

OAI221xp5_ASAP7_75t_L g2701 ( 
.A1(n_2642),
.A2(n_2646),
.B1(n_2586),
.B2(n_2623),
.C(n_2583),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2605),
.B(n_382),
.Y(n_2702)
);

AOI221xp5_ASAP7_75t_L g2703 ( 
.A1(n_2635),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.C(n_385),
.Y(n_2703)
);

AND4x1_ASAP7_75t_L g2704 ( 
.A(n_2579),
.B(n_387),
.C(n_385),
.D(n_386),
.Y(n_2704)
);

NAND3xp33_ASAP7_75t_SL g2705 ( 
.A(n_2601),
.B(n_386),
.C(n_388),
.Y(n_2705)
);

OAI211xp5_ASAP7_75t_SL g2706 ( 
.A1(n_2613),
.A2(n_391),
.B(n_388),
.C(n_389),
.Y(n_2706)
);

NOR3xp33_ASAP7_75t_SL g2707 ( 
.A(n_2640),
.B(n_389),
.C(n_391),
.Y(n_2707)
);

NAND3xp33_ASAP7_75t_SL g2708 ( 
.A(n_2617),
.B(n_392),
.C(n_393),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2587),
.B(n_392),
.Y(n_2709)
);

NOR3xp33_ASAP7_75t_L g2710 ( 
.A(n_2591),
.B(n_394),
.C(n_395),
.Y(n_2710)
);

AOI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2621),
.A2(n_394),
.B(n_395),
.Y(n_2711)
);

AND3x1_ASAP7_75t_L g2712 ( 
.A(n_2622),
.B(n_396),
.C(n_397),
.Y(n_2712)
);

AND3x2_ASAP7_75t_L g2713 ( 
.A(n_2584),
.B(n_396),
.C(n_397),
.Y(n_2713)
);

NOR3xp33_ASAP7_75t_L g2714 ( 
.A(n_2598),
.B(n_398),
.C(n_399),
.Y(n_2714)
);

AOI22xp33_ASAP7_75t_L g2715 ( 
.A1(n_2608),
.A2(n_2026),
.B1(n_401),
.B2(n_399),
.Y(n_2715)
);

NOR4xp25_ASAP7_75t_L g2716 ( 
.A(n_2600),
.B(n_403),
.C(n_400),
.D(n_401),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2639),
.Y(n_2717)
);

OAI221xp5_ASAP7_75t_L g2718 ( 
.A1(n_2612),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.C(n_406),
.Y(n_2718)
);

OAI211xp5_ASAP7_75t_L g2719 ( 
.A1(n_2632),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_2719)
);

NOR3xp33_ASAP7_75t_SL g2720 ( 
.A(n_2708),
.B(n_408),
.C(n_409),
.Y(n_2720)
);

INVx2_ASAP7_75t_SL g2721 ( 
.A(n_2713),
.Y(n_2721)
);

NAND3xp33_ASAP7_75t_SL g2722 ( 
.A(n_2654),
.B(n_2694),
.C(n_2658),
.Y(n_2722)
);

NAND3xp33_ASAP7_75t_SL g2723 ( 
.A(n_2652),
.B(n_408),
.C(n_409),
.Y(n_2723)
);

NOR2x1_ASAP7_75t_L g2724 ( 
.A(n_2665),
.B(n_410),
.Y(n_2724)
);

NOR2xp67_ASAP7_75t_L g2725 ( 
.A(n_2705),
.B(n_410),
.Y(n_2725)
);

AOI211xp5_ASAP7_75t_L g2726 ( 
.A1(n_2666),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_2726)
);

NOR2x1p5_ASAP7_75t_L g2727 ( 
.A(n_2679),
.B(n_411),
.Y(n_2727)
);

NOR4xp75_ASAP7_75t_L g2728 ( 
.A(n_2655),
.B(n_414),
.C(n_412),
.D(n_413),
.Y(n_2728)
);

NOR3xp33_ASAP7_75t_L g2729 ( 
.A(n_2695),
.B(n_2717),
.C(n_2673),
.Y(n_2729)
);

OAI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_2696),
.A2(n_415),
.B(n_416),
.Y(n_2730)
);

OAI211xp5_ASAP7_75t_L g2731 ( 
.A1(n_2719),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_2731)
);

OAI211xp5_ASAP7_75t_L g2732 ( 
.A1(n_2672),
.A2(n_420),
.B(n_417),
.C(n_419),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2669),
.B(n_419),
.Y(n_2733)
);

NAND4xp25_ASAP7_75t_L g2734 ( 
.A(n_2657),
.B(n_423),
.C(n_421),
.D(n_422),
.Y(n_2734)
);

NAND4xp75_ASAP7_75t_L g2735 ( 
.A(n_2712),
.B(n_424),
.C(n_421),
.D(n_423),
.Y(n_2735)
);

NAND4xp25_ASAP7_75t_L g2736 ( 
.A(n_2686),
.B(n_426),
.C(n_424),
.D(n_425),
.Y(n_2736)
);

NAND4xp75_ASAP7_75t_L g2737 ( 
.A(n_2667),
.B(n_428),
.C(n_426),
.D(n_427),
.Y(n_2737)
);

OA211x2_ASAP7_75t_L g2738 ( 
.A1(n_2685),
.A2(n_429),
.B(n_427),
.C(n_428),
.Y(n_2738)
);

HB1xp67_ASAP7_75t_L g2739 ( 
.A(n_2663),
.Y(n_2739)
);

NOR3xp33_ASAP7_75t_L g2740 ( 
.A(n_2718),
.B(n_429),
.C(n_430),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2653),
.B(n_2682),
.Y(n_2741)
);

NAND3xp33_ASAP7_75t_L g2742 ( 
.A(n_2687),
.B(n_430),
.C(n_432),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2704),
.Y(n_2743)
);

NAND4xp25_ASAP7_75t_SL g2744 ( 
.A(n_2715),
.B(n_434),
.C(n_432),
.D(n_433),
.Y(n_2744)
);

NOR3xp33_ASAP7_75t_L g2745 ( 
.A(n_2701),
.B(n_434),
.C(n_435),
.Y(n_2745)
);

NOR3xp33_ASAP7_75t_L g2746 ( 
.A(n_2702),
.B(n_2700),
.C(n_2680),
.Y(n_2746)
);

NAND5xp2_ASAP7_75t_L g2747 ( 
.A(n_2692),
.B(n_435),
.C(n_436),
.D(n_437),
.E(n_438),
.Y(n_2747)
);

NOR2x1_ASAP7_75t_L g2748 ( 
.A(n_2662),
.B(n_436),
.Y(n_2748)
);

NOR3x1_ASAP7_75t_L g2749 ( 
.A(n_2691),
.B(n_437),
.C(n_438),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2674),
.B(n_439),
.Y(n_2750)
);

OAI211xp5_ASAP7_75t_SL g2751 ( 
.A1(n_2707),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_2751)
);

NAND4xp25_ASAP7_75t_L g2752 ( 
.A(n_2676),
.B(n_443),
.C(n_440),
.D(n_442),
.Y(n_2752)
);

AOI211xp5_ASAP7_75t_L g2753 ( 
.A1(n_2697),
.A2(n_445),
.B(n_443),
.C(n_444),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_SL g2754 ( 
.A(n_2716),
.B(n_444),
.Y(n_2754)
);

OAI211xp5_ASAP7_75t_SL g2755 ( 
.A1(n_2690),
.A2(n_448),
.B(n_446),
.C(n_447),
.Y(n_2755)
);

AND4x1_ASAP7_75t_L g2756 ( 
.A(n_2678),
.B(n_449),
.C(n_446),
.D(n_447),
.Y(n_2756)
);

OAI211xp5_ASAP7_75t_SL g2757 ( 
.A1(n_2675),
.A2(n_2684),
.B(n_2688),
.C(n_2683),
.Y(n_2757)
);

NAND4xp75_ASAP7_75t_L g2758 ( 
.A(n_2711),
.B(n_451),
.C(n_449),
.D(n_450),
.Y(n_2758)
);

NAND3xp33_ASAP7_75t_L g2759 ( 
.A(n_2703),
.B(n_452),
.C(n_453),
.Y(n_2759)
);

OAI211xp5_ASAP7_75t_L g2760 ( 
.A1(n_2689),
.A2(n_454),
.B(n_452),
.C(n_453),
.Y(n_2760)
);

NOR2x1p5_ASAP7_75t_L g2761 ( 
.A(n_2661),
.B(n_454),
.Y(n_2761)
);

NOR2x1_ASAP7_75t_L g2762 ( 
.A(n_2659),
.B(n_455),
.Y(n_2762)
);

NAND4xp25_ASAP7_75t_L g2763 ( 
.A(n_2651),
.B(n_457),
.C(n_455),
.D(n_456),
.Y(n_2763)
);

NAND4xp75_ASAP7_75t_L g2764 ( 
.A(n_2656),
.B(n_459),
.C(n_456),
.D(n_457),
.Y(n_2764)
);

NOR2x1_ASAP7_75t_L g2765 ( 
.A(n_2671),
.B(n_459),
.Y(n_2765)
);

NAND3xp33_ASAP7_75t_L g2766 ( 
.A(n_2710),
.B(n_460),
.C(n_461),
.Y(n_2766)
);

NAND3xp33_ASAP7_75t_L g2767 ( 
.A(n_2714),
.B(n_460),
.C(n_461),
.Y(n_2767)
);

NOR2x1_ASAP7_75t_L g2768 ( 
.A(n_2660),
.B(n_462),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2668),
.B(n_463),
.Y(n_2769)
);

NAND3xp33_ASAP7_75t_L g2770 ( 
.A(n_2699),
.B(n_463),
.C(n_464),
.Y(n_2770)
);

AOI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2693),
.A2(n_464),
.B(n_465),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2698),
.B(n_2243),
.Y(n_2772)
);

NAND3xp33_ASAP7_75t_L g2773 ( 
.A(n_2681),
.B(n_466),
.C(n_467),
.Y(n_2773)
);

OAI211xp5_ASAP7_75t_SL g2774 ( 
.A1(n_2709),
.A2(n_2664),
.B(n_2706),
.C(n_2670),
.Y(n_2774)
);

NOR2x1_ASAP7_75t_L g2775 ( 
.A(n_2737),
.B(n_2735),
.Y(n_2775)
);

INVxp33_ASAP7_75t_SL g2776 ( 
.A(n_2739),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2724),
.Y(n_2777)
);

INVxp67_ASAP7_75t_SL g2778 ( 
.A(n_2725),
.Y(n_2778)
);

OA22x2_ASAP7_75t_L g2779 ( 
.A1(n_2730),
.A2(n_2677),
.B1(n_469),
.B2(n_466),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_SL g2780 ( 
.A1(n_2721),
.A2(n_2741),
.B1(n_2731),
.B2(n_2732),
.Y(n_2780)
);

NOR2x1_ASAP7_75t_L g2781 ( 
.A(n_2773),
.B(n_2677),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2753),
.B(n_468),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2764),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_2728),
.B(n_2743),
.Y(n_2784)
);

AOI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2729),
.A2(n_2026),
.B1(n_470),
.B2(n_468),
.Y(n_2785)
);

NOR2x1_ASAP7_75t_L g2786 ( 
.A(n_2734),
.B(n_469),
.Y(n_2786)
);

INVxp67_ASAP7_75t_L g2787 ( 
.A(n_2747),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2758),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2738),
.Y(n_2789)
);

OR2x2_ASAP7_75t_L g2790 ( 
.A(n_2736),
.B(n_470),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2756),
.Y(n_2791)
);

INVx2_ASAP7_75t_SL g2792 ( 
.A(n_2727),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2749),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2769),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2751),
.A2(n_474),
.B1(n_471),
.B2(n_472),
.Y(n_2795)
);

OR2x2_ASAP7_75t_L g2796 ( 
.A(n_2763),
.B(n_474),
.Y(n_2796)
);

NOR2x1_ASAP7_75t_L g2797 ( 
.A(n_2722),
.B(n_475),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2768),
.Y(n_2798)
);

NOR2x1_ASAP7_75t_L g2799 ( 
.A(n_2723),
.B(n_476),
.Y(n_2799)
);

INVxp67_ASAP7_75t_L g2800 ( 
.A(n_2748),
.Y(n_2800)
);

AND2x4_ASAP7_75t_L g2801 ( 
.A(n_2762),
.B(n_476),
.Y(n_2801)
);

NOR2x1_ASAP7_75t_SL g2802 ( 
.A(n_2754),
.B(n_2760),
.Y(n_2802)
);

OR2x2_ASAP7_75t_L g2803 ( 
.A(n_2752),
.B(n_478),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2733),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2765),
.B(n_478),
.Y(n_2805)
);

NOR2xp33_ASAP7_75t_L g2806 ( 
.A(n_2742),
.B(n_479),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2761),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2750),
.Y(n_2808)
);

NOR3xp33_ASAP7_75t_L g2809 ( 
.A(n_2757),
.B(n_480),
.C(n_481),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2770),
.Y(n_2810)
);

AND3x4_ASAP7_75t_L g2811 ( 
.A(n_2720),
.B(n_482),
.C(n_483),
.Y(n_2811)
);

XNOR2xp5_ASAP7_75t_L g2812 ( 
.A(n_2726),
.B(n_482),
.Y(n_2812)
);

AOI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2745),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_2813)
);

INVx1_ASAP7_75t_SL g2814 ( 
.A(n_2771),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2759),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2772),
.Y(n_2816)
);

AOI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2744),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_2817)
);

OA22x2_ASAP7_75t_L g2818 ( 
.A1(n_2755),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2766),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2740),
.B(n_2243),
.Y(n_2820)
);

INVx1_ASAP7_75t_SL g2821 ( 
.A(n_2767),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_SL g2822 ( 
.A(n_2746),
.B(n_488),
.Y(n_2822)
);

NOR2x1_ASAP7_75t_L g2823 ( 
.A(n_2774),
.B(n_489),
.Y(n_2823)
);

NOR3xp33_ASAP7_75t_L g2824 ( 
.A(n_2780),
.B(n_490),
.C(n_491),
.Y(n_2824)
);

NOR2x1_ASAP7_75t_L g2825 ( 
.A(n_2797),
.B(n_2781),
.Y(n_2825)
);

AND2x4_ASAP7_75t_SL g2826 ( 
.A(n_2784),
.B(n_2789),
.Y(n_2826)
);

NOR3xp33_ASAP7_75t_L g2827 ( 
.A(n_2798),
.B(n_490),
.C(n_491),
.Y(n_2827)
);

NOR3xp33_ASAP7_75t_L g2828 ( 
.A(n_2777),
.B(n_2778),
.C(n_2800),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2809),
.B(n_492),
.Y(n_2829)
);

NAND3xp33_ASAP7_75t_L g2830 ( 
.A(n_2823),
.B(n_492),
.C(n_493),
.Y(n_2830)
);

AOI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2776),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2817),
.B(n_494),
.Y(n_2832)
);

NOR2x1_ASAP7_75t_L g2833 ( 
.A(n_2801),
.B(n_496),
.Y(n_2833)
);

NAND4xp25_ASAP7_75t_L g2834 ( 
.A(n_2795),
.B(n_496),
.C(n_497),
.D(n_498),
.Y(n_2834)
);

AND2x4_ASAP7_75t_L g2835 ( 
.A(n_2775),
.B(n_497),
.Y(n_2835)
);

O2A1O1Ixp33_ASAP7_75t_L g2836 ( 
.A1(n_2822),
.A2(n_498),
.B(n_499),
.C(n_500),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_L g2837 ( 
.A(n_2788),
.B(n_500),
.C(n_502),
.Y(n_2837)
);

AND2x4_ASAP7_75t_L g2838 ( 
.A(n_2791),
.B(n_503),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2779),
.Y(n_2839)
);

NAND4xp75_ASAP7_75t_L g2840 ( 
.A(n_2799),
.B(n_505),
.C(n_506),
.D(n_507),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2818),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2813),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_2842)
);

NAND2x1p5_ASAP7_75t_L g2843 ( 
.A(n_2783),
.B(n_508),
.Y(n_2843)
);

OR2x2_ASAP7_75t_L g2844 ( 
.A(n_2790),
.B(n_509),
.Y(n_2844)
);

NOR3xp33_ASAP7_75t_L g2845 ( 
.A(n_2792),
.B(n_510),
.C(n_512),
.Y(n_2845)
);

NOR2x1_ASAP7_75t_L g2846 ( 
.A(n_2801),
.B(n_512),
.Y(n_2846)
);

NAND3xp33_ASAP7_75t_SL g2847 ( 
.A(n_2821),
.B(n_513),
.C(n_514),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2796),
.Y(n_2848)
);

NAND4xp75_ASAP7_75t_L g2849 ( 
.A(n_2786),
.B(n_513),
.C(n_514),
.D(n_515),
.Y(n_2849)
);

AND4x1_ASAP7_75t_L g2850 ( 
.A(n_2815),
.B(n_516),
.C(n_517),
.D(n_518),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2803),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2805),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2787),
.B(n_2290),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2793),
.B(n_516),
.Y(n_2854)
);

OAI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2830),
.A2(n_2785),
.B1(n_2811),
.B2(n_2819),
.Y(n_2855)
);

NOR3xp33_ASAP7_75t_L g2856 ( 
.A(n_2825),
.B(n_2807),
.C(n_2814),
.Y(n_2856)
);

AOI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2829),
.A2(n_2782),
.B(n_2802),
.Y(n_2857)
);

NOR3x2_ASAP7_75t_L g2858 ( 
.A(n_2840),
.B(n_2805),
.C(n_2812),
.Y(n_2858)
);

NOR3x1_ASAP7_75t_L g2859 ( 
.A(n_2849),
.B(n_2847),
.C(n_2844),
.Y(n_2859)
);

OAI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2832),
.A2(n_2806),
.B1(n_2810),
.B2(n_2816),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2833),
.Y(n_2861)
);

AOI221xp5_ASAP7_75t_L g2862 ( 
.A1(n_2828),
.A2(n_2808),
.B1(n_2804),
.B2(n_2794),
.C(n_2820),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2846),
.Y(n_2863)
);

NOR2x1p5_ASAP7_75t_L g2864 ( 
.A(n_2834),
.B(n_518),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2852),
.A2(n_519),
.B(n_520),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_2843),
.B(n_519),
.Y(n_2866)
);

NAND2xp33_ASAP7_75t_SL g2867 ( 
.A(n_2835),
.B(n_521),
.Y(n_2867)
);

NAND4xp75_ASAP7_75t_L g2868 ( 
.A(n_2839),
.B(n_521),
.C(n_522),
.D(n_523),
.Y(n_2868)
);

NOR4xp25_ASAP7_75t_L g2869 ( 
.A(n_2841),
.B(n_522),
.C(n_524),
.D(n_525),
.Y(n_2869)
);

AO22x2_ASAP7_75t_L g2870 ( 
.A1(n_2851),
.A2(n_2848),
.B1(n_2824),
.B2(n_2842),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_2850),
.Y(n_2871)
);

CKINVDCx5p33_ASAP7_75t_R g2872 ( 
.A(n_2826),
.Y(n_2872)
);

AOI221xp5_ASAP7_75t_L g2873 ( 
.A1(n_2836),
.A2(n_524),
.B1(n_526),
.B2(n_527),
.C(n_528),
.Y(n_2873)
);

AND2x4_ASAP7_75t_L g2874 ( 
.A(n_2837),
.B(n_526),
.Y(n_2874)
);

OAI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2853),
.A2(n_527),
.B1(n_528),
.B2(n_529),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2845),
.B(n_529),
.Y(n_2876)
);

AND2x4_ASAP7_75t_L g2877 ( 
.A(n_2827),
.B(n_530),
.Y(n_2877)
);

OAI221xp5_ASAP7_75t_L g2878 ( 
.A1(n_2831),
.A2(n_530),
.B1(n_532),
.B2(n_533),
.C(n_534),
.Y(n_2878)
);

OAI21xp33_ASAP7_75t_SL g2879 ( 
.A1(n_2854),
.A2(n_532),
.B(n_533),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_2838),
.Y(n_2880)
);

AOI31xp33_ASAP7_75t_L g2881 ( 
.A1(n_2833),
.A2(n_534),
.A3(n_535),
.B(n_536),
.Y(n_2881)
);

NOR2x1_ASAP7_75t_L g2882 ( 
.A(n_2833),
.B(n_535),
.Y(n_2882)
);

NAND4xp25_ASAP7_75t_L g2883 ( 
.A(n_2828),
.B(n_536),
.C(n_537),
.D(n_538),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2833),
.Y(n_2884)
);

BUFx6f_ASAP7_75t_L g2885 ( 
.A(n_2852),
.Y(n_2885)
);

BUFx12f_ASAP7_75t_L g2886 ( 
.A(n_2826),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_SL g2887 ( 
.A1(n_2826),
.A2(n_537),
.B1(n_538),
.B2(n_539),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2825),
.A2(n_539),
.B(n_542),
.Y(n_2888)
);

O2A1O1Ixp33_ASAP7_75t_L g2889 ( 
.A1(n_2828),
.A2(n_542),
.B(n_543),
.C(n_544),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2824),
.B(n_543),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2833),
.Y(n_2891)
);

NAND3x1_ASAP7_75t_L g2892 ( 
.A(n_2833),
.B(n_544),
.C(n_545),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2866),
.Y(n_2893)
);

NAND4xp25_ASAP7_75t_L g2894 ( 
.A(n_2856),
.B(n_2862),
.C(n_2859),
.D(n_2857),
.Y(n_2894)
);

OR2x2_ASAP7_75t_L g2895 ( 
.A(n_2869),
.B(n_546),
.Y(n_2895)
);

XNOR2xp5_ASAP7_75t_L g2896 ( 
.A(n_2872),
.B(n_546),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_2886),
.B(n_547),
.Y(n_2897)
);

NAND4xp75_ASAP7_75t_L g2898 ( 
.A(n_2882),
.B(n_548),
.C(n_549),
.D(n_550),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2868),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2881),
.B(n_549),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2879),
.B(n_550),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2892),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2864),
.B(n_2871),
.Y(n_2903)
);

NOR3xp33_ASAP7_75t_SL g2904 ( 
.A(n_2867),
.B(n_551),
.C(n_552),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2890),
.Y(n_2905)
);

INVx3_ASAP7_75t_L g2906 ( 
.A(n_2858),
.Y(n_2906)
);

NOR2x1_ASAP7_75t_L g2907 ( 
.A(n_2861),
.B(n_551),
.Y(n_2907)
);

NOR2x1p5_ASAP7_75t_L g2908 ( 
.A(n_2885),
.B(n_552),
.Y(n_2908)
);

NOR2xp67_ASAP7_75t_L g2909 ( 
.A(n_2883),
.B(n_553),
.Y(n_2909)
);

AND2x4_ASAP7_75t_L g2910 ( 
.A(n_2885),
.B(n_553),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2873),
.B(n_554),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2877),
.B(n_2264),
.Y(n_2912)
);

NAND3xp33_ASAP7_75t_SL g2913 ( 
.A(n_2880),
.B(n_554),
.C(n_555),
.Y(n_2913)
);

HB1xp67_ASAP7_75t_L g2914 ( 
.A(n_2863),
.Y(n_2914)
);

NAND4xp75_ASAP7_75t_L g2915 ( 
.A(n_2884),
.B(n_555),
.C(n_556),
.D(n_557),
.Y(n_2915)
);

XNOR2x1_ASAP7_75t_L g2916 ( 
.A(n_2870),
.B(n_558),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2874),
.Y(n_2917)
);

AOI22x1_ASAP7_75t_L g2918 ( 
.A1(n_2914),
.A2(n_2870),
.B1(n_2891),
.B2(n_2888),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2909),
.B(n_2889),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2916),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2915),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2908),
.Y(n_2922)
);

OAI22xp5_ASAP7_75t_SL g2923 ( 
.A1(n_2899),
.A2(n_2855),
.B1(n_2860),
.B2(n_2878),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_SL g2924 ( 
.A(n_2900),
.B(n_2865),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2907),
.Y(n_2925)
);

OAI211xp5_ASAP7_75t_SL g2926 ( 
.A1(n_2906),
.A2(n_2876),
.B(n_2887),
.C(n_2875),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2895),
.Y(n_2927)
);

AOI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2913),
.A2(n_559),
.B1(n_560),
.B2(n_561),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2897),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2898),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2896),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2901),
.Y(n_2932)
);

AOI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2894),
.A2(n_559),
.B1(n_562),
.B2(n_563),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2904),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2910),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2902),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2893),
.Y(n_2937)
);

AOI22xp33_ASAP7_75t_L g2938 ( 
.A1(n_2918),
.A2(n_2917),
.B1(n_2905),
.B2(n_2911),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2935),
.Y(n_2939)
);

AND3x2_ASAP7_75t_L g2940 ( 
.A(n_2925),
.B(n_2903),
.C(n_2912),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2922),
.Y(n_2941)
);

INVx3_ASAP7_75t_L g2942 ( 
.A(n_2921),
.Y(n_2942)
);

AND2x4_ASAP7_75t_L g2943 ( 
.A(n_2930),
.B(n_2937),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2928),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2933),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2936),
.B(n_562),
.Y(n_2946)
);

AO22x2_ASAP7_75t_L g2947 ( 
.A1(n_2934),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_2947)
);

XOR2xp5_ASAP7_75t_L g2948 ( 
.A(n_2923),
.B(n_565),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2927),
.Y(n_2949)
);

AOI22x1_ASAP7_75t_L g2950 ( 
.A1(n_2920),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_2950)
);

BUFx2_ASAP7_75t_SL g2951 ( 
.A(n_2939),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2948),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2950),
.Y(n_2953)
);

INVxp67_ASAP7_75t_SL g2954 ( 
.A(n_2942),
.Y(n_2954)
);

OAI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2943),
.A2(n_2919),
.B(n_2926),
.Y(n_2955)
);

HB1xp67_ASAP7_75t_L g2956 ( 
.A(n_2941),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2947),
.Y(n_2957)
);

OAI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2954),
.A2(n_2938),
.B1(n_2949),
.B2(n_2932),
.Y(n_2958)
);

INVx4_ASAP7_75t_L g2959 ( 
.A(n_2956),
.Y(n_2959)
);

XNOR2x1_ASAP7_75t_L g2960 ( 
.A(n_2955),
.B(n_2940),
.Y(n_2960)
);

OR2x6_ASAP7_75t_L g2961 ( 
.A(n_2951),
.B(n_2931),
.Y(n_2961)
);

AOI22xp5_ASAP7_75t_SL g2962 ( 
.A1(n_2957),
.A2(n_2929),
.B1(n_2945),
.B2(n_2944),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2953),
.B(n_2924),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2952),
.Y(n_2964)
);

OAI21xp33_ASAP7_75t_L g2965 ( 
.A1(n_2960),
.A2(n_2946),
.B(n_568),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2959),
.Y(n_2966)
);

OAI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2958),
.A2(n_567),
.B(n_569),
.Y(n_2967)
);

OAI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2961),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2965),
.B(n_2962),
.Y(n_2969)
);

OAI22x1_ASAP7_75t_SL g2970 ( 
.A1(n_2966),
.A2(n_2964),
.B1(n_2963),
.B2(n_2967),
.Y(n_2970)
);

OA22x2_ASAP7_75t_L g2971 ( 
.A1(n_2968),
.A2(n_570),
.B1(n_571),
.B2(n_572),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2970),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2969),
.Y(n_2973)
);

OR2x2_ASAP7_75t_L g2974 ( 
.A(n_2971),
.B(n_572),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2974),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2972),
.B(n_573),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2975),
.Y(n_2977)
);

OAI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2977),
.A2(n_2973),
.B1(n_2976),
.B2(n_576),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2978),
.Y(n_2979)
);

AOI22xp33_ASAP7_75t_SL g2980 ( 
.A1(n_2979),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.Y(n_2980)
);

AOI221xp5_ASAP7_75t_L g2981 ( 
.A1(n_2980),
.A2(n_574),
.B1(n_575),
.B2(n_577),
.C(n_578),
.Y(n_2981)
);

AOI21xp33_ASAP7_75t_L g2982 ( 
.A1(n_2981),
.A2(n_577),
.B(n_578),
.Y(n_2982)
);

AOI211xp5_ASAP7_75t_L g2983 ( 
.A1(n_2982),
.A2(n_579),
.B(n_580),
.C(n_581),
.Y(n_2983)
);


endmodule