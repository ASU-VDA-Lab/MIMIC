module fake_jpeg_19882_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_57),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_28),
.B1(n_20),
.B2(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_39),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_20),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_22),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_28),
.B1(n_20),
.B2(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_27),
.B1(n_22),
.B2(n_25),
.Y(n_81)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_30),
.B1(n_19),
.B2(n_33),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_41),
.B1(n_34),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_21),
.B1(n_32),
.B2(n_30),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_21),
.B1(n_29),
.B2(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_23),
.B1(n_17),
.B2(n_24),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_17),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_43),
.B1(n_48),
.B2(n_54),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_69),
.A2(n_90),
.B1(n_54),
.B2(n_59),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_26),
.B(n_31),
.C(n_33),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_77),
.B(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_82),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_41),
.B1(n_38),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_81),
.B1(n_63),
.B2(n_89),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_31),
.B(n_24),
.C(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_18),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_27),
.B1(n_9),
.B2(n_10),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_R g95 ( 
.A(n_70),
.B(n_60),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_112),
.B(n_73),
.Y(n_122)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_100),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_109),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_54),
.B1(n_58),
.B2(n_47),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_115),
.B1(n_83),
.B2(n_74),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_83),
.B(n_77),
.Y(n_140)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_117),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_93),
.Y(n_123)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_82),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_123),
.Y(n_162)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_127),
.Y(n_181)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_137),
.B1(n_148),
.B2(n_120),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_69),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_110),
.B(n_114),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_72),
.B1(n_80),
.B2(n_61),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_62),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_69),
.B(n_77),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_83),
.B(n_69),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_91),
.B(n_96),
.Y(n_177)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_137),
.B1(n_122),
.B2(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_70),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_79),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_69),
.B1(n_90),
.B2(n_86),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_84),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_51),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_151),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_107),
.B(n_75),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_153),
.A2(n_175),
.B(n_177),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_125),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_102),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_157),
.B(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_112),
.B1(n_102),
.B2(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_164),
.B1(n_183),
.B2(n_185),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_112),
.B1(n_81),
.B2(n_98),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_120),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_168),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_180),
.B1(n_126),
.B2(n_124),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_113),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_113),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_150),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_51),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_139),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_178),
.Y(n_213)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_96),
.B(n_118),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_125),
.B(n_149),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_88),
.B1(n_99),
.B2(n_97),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_129),
.A2(n_94),
.B1(n_54),
.B2(n_59),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_131),
.B(n_137),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_94),
.B1(n_11),
.B2(n_12),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_135),
.C(n_123),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_196),
.C(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_194),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_122),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_199),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_192),
.B(n_203),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_137),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_208),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_132),
.C(n_146),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_197),
.B(n_175),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_129),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_124),
.C(n_142),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_142),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_214),
.C(n_174),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_142),
.B(n_130),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_182),
.B1(n_176),
.B2(n_154),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_27),
.B1(n_18),
.B2(n_25),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_156),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_171),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_59),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_160),
.A2(n_25),
.B1(n_18),
.B2(n_15),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_152),
.B1(n_180),
.B2(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_219),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_169),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_221),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_181),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_153),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_211),
.A2(n_182),
.B(n_160),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_224),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_204),
.B1(n_191),
.B2(n_188),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_152),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_235),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_164),
.C(n_158),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_230),
.C(n_196),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_179),
.C(n_154),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_238),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_198),
.B1(n_199),
.B2(n_187),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_239),
.A2(n_244),
.B1(n_247),
.B2(n_49),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_190),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_251),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_245),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_194),
.B1(n_187),
.B2(n_193),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_49),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_195),
.B1(n_202),
.B2(n_207),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_205),
.B1(n_175),
.B2(n_200),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_186),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_250),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_201),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_214),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_203),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_258),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_211),
.C(n_159),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_257),
.C(n_229),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_233),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_159),
.C(n_178),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_221),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_217),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_261),
.B(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_265),
.C(n_267),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_222),
.B(n_218),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_266),
.B(n_0),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_257),
.C(n_250),
.Y(n_265)
);

OAI22x1_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_226),
.B1(n_223),
.B2(n_225),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_255),
.C(n_245),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_226),
.B(n_225),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_252),
.B(n_15),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_227),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_49),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_276),
.B(n_281),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_12),
.B(n_11),
.C(n_10),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_278),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_0),
.C(n_1),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_284),
.C(n_288),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_0),
.C(n_1),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_269),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_287),
.Y(n_291)
);

NAND2xp67_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_1),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_2),
.C(n_3),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_268),
.B(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_293),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_284),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_282),
.A2(n_274),
.B1(n_279),
.B2(n_286),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_263),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_299),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_259),
.B(n_260),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_298),
.A2(n_288),
.B(n_283),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_263),
.B1(n_259),
.B2(n_4),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_303),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.C(n_294),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_2),
.C(n_3),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_304)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_306),
.C(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_4),
.C(n_5),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_4),
.B(n_6),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_296),
.C(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_291),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_312),
.C(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_294),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_302),
.B(n_308),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_314),
.Y(n_316)
);

AOI321xp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_315),
.C(n_311),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_7),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_7),
.Y(n_319)
);


endmodule