module fake_jpeg_21822_n_28 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_6),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_6),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_4),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.C(n_1),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.C(n_9),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_11),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_13),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_25),
.B(n_22),
.Y(n_26)
);

AOI322xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_8),
.A3(n_17),
.B1(n_23),
.B2(n_24),
.C1(n_14),
.C2(n_20),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_24),
.Y(n_28)
);


endmodule