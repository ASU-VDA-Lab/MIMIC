module fake_netlist_6_4285_n_739 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_739);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_739;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_6),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_68),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_28),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_84),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_35),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_42),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_40),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_46),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_36),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_11),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_96),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_94),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_66),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_121),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_3),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_103),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_49),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_14),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_48),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_52),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_23),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_72),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_53),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_24),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_142),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_59),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_93),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_97),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_56),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_135),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_51),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_38),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_137),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_45),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_2),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_74),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_150),
.B(n_0),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_20),
.Y(n_204)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_1),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_3),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_21),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_22),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

AOI22x1_ASAP7_75t_SL g220 ( 
.A1(n_173),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_25),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_26),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_5),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_27),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_147),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_7),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_173),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_8),
.B(n_9),
.Y(n_234)
);

BUFx8_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

BUFx8_ASAP7_75t_L g238 ( 
.A(n_147),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_152),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_179),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

CKINVDCx6p67_ASAP7_75t_R g243 ( 
.A(n_156),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_29),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_10),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

CKINVDCx6p67_ASAP7_75t_R g249 ( 
.A(n_243),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

BUFx8_ASAP7_75t_SL g255 ( 
.A(n_242),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_217),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_204),
.B(n_207),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_201),
.B(n_161),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_200),
.C(n_195),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_154),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

AND3x2_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_10),
.C(n_11),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_205),
.B(n_157),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_204),
.B(n_159),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_162),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_210),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_233),
.B(n_12),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_208),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_216),
.B(n_165),
.Y(n_278)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_230),
.B(n_194),
.C(n_193),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_228),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_190),
.B1(n_189),
.B2(n_188),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_216),
.B(n_166),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_212),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_216),
.B(n_221),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_240),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_241),
.B1(n_220),
.B2(n_211),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_221),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_241),
.C(n_203),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_221),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_209),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_222),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_222),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_222),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_284),
.B(n_227),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_244),
.A2(n_227),
.B1(n_234),
.B2(n_219),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_268),
.A2(n_227),
.B1(n_174),
.B2(n_169),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

BUFx6f_ASAP7_75t_SL g312 ( 
.A(n_275),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_281),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_245),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g315 ( 
.A1(n_260),
.A2(n_209),
.B1(n_167),
.B2(n_184),
.C(n_171),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_232),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_232),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_235),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_257),
.B(n_235),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_247),
.B(n_172),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_253),
.Y(n_327)
);

BUFx6f_ASAP7_75t_SL g328 ( 
.A(n_244),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_248),
.A2(n_234),
.B(n_186),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_229),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_266),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g332 ( 
.A(n_252),
.B(n_183),
.C(n_238),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_246),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_229),
.Y(n_335)
);

BUFx8_ASAP7_75t_L g336 ( 
.A(n_249),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_254),
.A2(n_265),
.B1(n_288),
.B2(n_235),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_231),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_282),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_283),
.B(n_231),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_255),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_231),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_246),
.B(n_238),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_297),
.B(n_238),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_255),
.Y(n_346)
);

O2A1O1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_298),
.A2(n_290),
.B(n_258),
.C(n_251),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_212),
.B1(n_258),
.B2(n_251),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_290),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_305),
.A2(n_212),
.B(n_250),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_250),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_307),
.A2(n_303),
.B(n_309),
.C(n_308),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_13),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_212),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_13),
.C(n_14),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_291),
.B(n_30),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_296),
.B(n_31),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_319),
.A2(n_89),
.B(n_145),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_88),
.B1(n_144),
.B2(n_143),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_318),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_SL g365 ( 
.A(n_299),
.B(n_15),
.C(n_16),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_321),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_300),
.B(n_18),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_32),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_317),
.A2(n_19),
.B(n_33),
.C(n_34),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_37),
.B(n_39),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_310),
.A2(n_326),
.B(n_343),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_335),
.A2(n_50),
.B(n_54),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_328),
.A2(n_55),
.B1(n_58),
.B2(n_60),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_338),
.A2(n_61),
.B(n_62),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_340),
.A2(n_63),
.B(n_64),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_324),
.B(n_65),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_342),
.A2(n_339),
.B(n_325),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

CKINVDCx8_ASAP7_75t_R g386 ( 
.A(n_320),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_292),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_311),
.A2(n_75),
.B(n_76),
.Y(n_389)
);

O2A1O1Ixp5_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_77),
.B(n_78),
.C(n_80),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_341),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_333),
.A2(n_81),
.B(n_82),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_294),
.B(n_85),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_86),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_333),
.A2(n_87),
.B(n_90),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_337),
.A2(n_91),
.B(n_92),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_337),
.A2(n_294),
.B(n_328),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_294),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_294),
.B(n_95),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_312),
.A2(n_98),
.B(n_99),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_298),
.B(n_100),
.Y(n_401)
);

OR2x6_ASAP7_75t_L g402 ( 
.A(n_327),
.B(n_101),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_352),
.B(n_102),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_349),
.A2(n_104),
.B(n_105),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_108),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_398),
.A2(n_109),
.B(n_110),
.Y(n_406)
);

OAI22x1_ASAP7_75t_L g407 ( 
.A1(n_388),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g409 ( 
.A(n_371),
.B(n_117),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_384),
.A2(n_139),
.B(n_122),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_401),
.A2(n_118),
.B(n_123),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_369),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_350),
.A2(n_124),
.B(n_126),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_351),
.B(n_127),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

OAI21x1_ASAP7_75t_SL g417 ( 
.A1(n_397),
.A2(n_128),
.B(n_129),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_355),
.A2(n_130),
.B(n_131),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_368),
.A2(n_357),
.B(n_399),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_360),
.B(n_132),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_376),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_357),
.A2(n_133),
.B(n_136),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_375),
.A2(n_138),
.B(n_347),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_360),
.B(n_383),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_393),
.A2(n_348),
.B(n_359),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_363),
.A2(n_374),
.B(n_362),
.Y(n_430)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_396),
.A2(n_400),
.B(n_381),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_373),
.A2(n_377),
.B(n_380),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_370),
.A2(n_378),
.B(n_390),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_354),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_358),
.B(n_356),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_389),
.A2(n_392),
.B(n_395),
.Y(n_438)
);

NAND2x1p5_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_388),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_366),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_345),
.A2(n_365),
.B(n_385),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_346),
.A2(n_402),
.B(n_386),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_391),
.A2(n_289),
.B(n_298),
.Y(n_444)
);

AOI21xp33_ASAP7_75t_L g445 ( 
.A1(n_387),
.A2(n_305),
.B(n_306),
.Y(n_445)
);

AO21x2_ASAP7_75t_L g446 ( 
.A1(n_352),
.A2(n_350),
.B(n_401),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_352),
.B(n_297),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_351),
.B(n_297),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_356),
.A2(n_289),
.B1(n_302),
.B2(n_298),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_351),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_352),
.B(n_297),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_352),
.A2(n_289),
.B(n_298),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_352),
.A2(n_289),
.B(n_298),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_352),
.A2(n_309),
.B(n_398),
.Y(n_455)
);

AO21x2_ASAP7_75t_L g456 ( 
.A1(n_427),
.A2(n_454),
.B(n_453),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_422),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_436),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_439),
.A2(n_447),
.B(n_452),
.C(n_437),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_420),
.A2(n_431),
.B(n_434),
.Y(n_461)
);

OAI21x1_ASAP7_75t_SL g462 ( 
.A1(n_417),
.A2(n_421),
.B(n_406),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_410),
.A2(n_429),
.B(n_438),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_450),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_426),
.Y(n_465)
);

BUFx2_ASAP7_75t_SL g466 ( 
.A(n_451),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_409),
.Y(n_469)
);

AO21x2_ASAP7_75t_L g470 ( 
.A1(n_455),
.A2(n_403),
.B(n_435),
.Y(n_470)
);

OA21x2_ASAP7_75t_L g471 ( 
.A1(n_406),
.A2(n_430),
.B(n_449),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_L g472 ( 
.A(n_413),
.B(n_423),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_449),
.A2(n_440),
.B(n_405),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_414),
.A2(n_404),
.B(n_419),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_416),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_436),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_411),
.A2(n_425),
.B(n_444),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_439),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_428),
.A2(n_446),
.B(n_415),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_445),
.B(n_416),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_423),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_445),
.A2(n_418),
.B(n_424),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_432),
.Y(n_484)
);

INVx8_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_413),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_441),
.A2(n_446),
.B(n_407),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_228),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_408),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_408),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_427),
.A2(n_454),
.B(n_453),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_409),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_439),
.A2(n_356),
.B1(n_437),
.B2(n_312),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_448),
.B(n_242),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g497 ( 
.A1(n_409),
.A2(n_312),
.B1(n_439),
.B2(n_238),
.Y(n_497)
);

AO21x2_ASAP7_75t_L g498 ( 
.A1(n_427),
.A2(n_454),
.B(n_453),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_468),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_476),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_476),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_470),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_459),
.B(n_495),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_458),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_460),
.A2(n_479),
.B(n_482),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

CKINVDCx6p67_ASAP7_75t_R g510 ( 
.A(n_483),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_478),
.B(n_464),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_478),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_464),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_483),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_472),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_457),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_457),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

CKINVDCx12_ASAP7_75t_R g522 ( 
.A(n_496),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_466),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_475),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_493),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_469),
.A2(n_493),
.B1(n_497),
.B2(n_471),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_465),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_484),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_475),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_488),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_488),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_475),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_473),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_484),
.B(n_471),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_475),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_473),
.B(n_471),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_535),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_535),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_502),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_519),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_513),
.B(n_484),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_525),
.B(n_469),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_512),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_501),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_531),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_531),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_513),
.B(n_473),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_511),
.B(n_517),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_505),
.B(n_480),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_514),
.B(n_517),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_526),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_536),
.B(n_480),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_519),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_520),
.B(n_481),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_526),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_536),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_533),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_527),
.A2(n_462),
.B1(n_498),
.B2(n_456),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_502),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_516),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_536),
.B(n_456),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_528),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_512),
.B(n_485),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_528),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_529),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_500),
.B(n_481),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_500),
.B(n_506),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_508),
.A2(n_529),
.B1(n_456),
.B2(n_498),
.Y(n_575)
);

NOR2x1_ASAP7_75t_L g576 ( 
.A(n_518),
.B(n_492),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_509),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_523),
.B(n_485),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_529),
.B(n_481),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_574),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_538),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_545),
.A2(n_477),
.B(n_474),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_532),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_503),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_577),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_577),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_551),
.B(n_530),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_552),
.B(n_532),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_540),
.B(n_522),
.Y(n_589)
);

INVx2_ASAP7_75t_R g590 ( 
.A(n_539),
.Y(n_590)
);

OAI221xp5_ASAP7_75t_SL g591 ( 
.A1(n_564),
.A2(n_522),
.B1(n_510),
.B2(n_521),
.C(n_518),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_539),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_541),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_555),
.B(n_532),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_573),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_550),
.B(n_538),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_541),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_573),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_499),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_548),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_548),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_544),
.B(n_521),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_553),
.B(n_571),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_555),
.B(n_515),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_547),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_547),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_553),
.B(n_499),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_546),
.B(n_554),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_571),
.B(n_499),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_549),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_549),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_559),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_559),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_542),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_554),
.B(n_515),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_576),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_563),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_581),
.B(n_563),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_611),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_581),
.B(n_567),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_614),
.B(n_576),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_611),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_596),
.B(n_567),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_608),
.B(n_547),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_562),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_612),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_587),
.B(n_557),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_596),
.B(n_562),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_603),
.B(n_557),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_594),
.B(n_557),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_591),
.B(n_569),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_582),
.A2(n_578),
.B(n_575),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_612),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_603),
.B(n_568),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_595),
.B(n_568),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_599),
.B(n_562),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_613),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_602),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_613),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_617),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_584),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_599),
.B(n_562),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_617),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_598),
.B(n_570),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_602),
.B(n_570),
.Y(n_645)
);

NOR2x1_ASAP7_75t_L g646 ( 
.A(n_616),
.B(n_565),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_609),
.B(n_515),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_600),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_609),
.B(n_504),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_605),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_602),
.B(n_561),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_606),
.B(n_561),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_633),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_633),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_640),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_640),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_619),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_628),
.B(n_616),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_622),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_627),
.B(n_583),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_641),
.B(n_589),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_626),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_637),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_628),
.B(n_590),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_624),
.B(n_583),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_638),
.B(n_607),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_636),
.B(n_590),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_639),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_645),
.B(n_588),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_643),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_648),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

NOR2x1p5_ASAP7_75t_SL g673 ( 
.A(n_654),
.B(n_630),
.Y(n_673)
);

OAI32xp33_ASAP7_75t_L g674 ( 
.A1(n_661),
.A2(n_631),
.A3(n_629),
.B1(n_651),
.B2(n_634),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_665),
.B(n_620),
.Y(n_675)
);

AOI222xp33_ASAP7_75t_L g676 ( 
.A1(n_661),
.A2(n_632),
.B1(n_631),
.B2(n_618),
.C1(n_652),
.C2(n_572),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_669),
.B(n_660),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_666),
.B(n_623),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_668),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_658),
.B(n_636),
.Y(n_680)
);

OAI32xp33_ASAP7_75t_L g681 ( 
.A1(n_657),
.A2(n_644),
.A3(n_635),
.B1(n_621),
.B2(n_610),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_672),
.Y(n_682)
);

AOI211xp5_ASAP7_75t_L g683 ( 
.A1(n_659),
.A2(n_477),
.B(n_650),
.C(n_572),
.Y(n_683)
);

NAND3xp33_ASAP7_75t_SL g684 ( 
.A(n_662),
.B(n_621),
.C(n_588),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_668),
.Y(n_685)
);

AOI222xp33_ASAP7_75t_L g686 ( 
.A1(n_663),
.A2(n_649),
.B1(n_647),
.B2(n_642),
.C1(n_607),
.C2(n_615),
.Y(n_686)
);

AO21x1_ASAP7_75t_L g687 ( 
.A1(n_683),
.A2(n_670),
.B(n_653),
.Y(n_687)
);

NAND5xp2_ASAP7_75t_L g688 ( 
.A(n_676),
.B(n_664),
.C(n_667),
.D(n_658),
.E(n_642),
.Y(n_688)
);

OAI221xp5_ASAP7_75t_SL g689 ( 
.A1(n_683),
.A2(n_664),
.B1(n_667),
.B2(n_671),
.C(n_656),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_679),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_685),
.Y(n_691)
);

BUFx2_ASAP7_75t_SL g692 ( 
.A(n_682),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_674),
.A2(n_614),
.B1(n_625),
.B2(n_650),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_693),
.A2(n_684),
.B(n_681),
.Y(n_694)
);

AOI222xp33_ASAP7_75t_L g695 ( 
.A1(n_688),
.A2(n_673),
.B1(n_678),
.B2(n_671),
.C1(n_655),
.C2(n_654),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_687),
.A2(n_686),
.B1(n_677),
.B2(n_625),
.Y(n_696)
);

OAI21xp33_ASAP7_75t_L g697 ( 
.A1(n_689),
.A2(n_675),
.B(n_646),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_690),
.B(n_680),
.Y(n_698)
);

AOI221xp5_ASAP7_75t_L g699 ( 
.A1(n_687),
.A2(n_601),
.B1(n_625),
.B2(n_592),
.C(n_597),
.Y(n_699)
);

NAND4xp25_ASAP7_75t_L g700 ( 
.A(n_697),
.B(n_691),
.C(n_516),
.D(n_594),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_696),
.B(n_691),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_698),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_694),
.B(n_692),
.Y(n_703)
);

OAI211xp5_ASAP7_75t_L g704 ( 
.A1(n_695),
.A2(n_592),
.B(n_593),
.C(n_597),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_703),
.B(n_699),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_702),
.B(n_510),
.Y(n_706)
);

NOR3xp33_ASAP7_75t_L g707 ( 
.A(n_704),
.B(n_566),
.C(n_579),
.Y(n_707)
);

NOR2x1p5_ASAP7_75t_L g708 ( 
.A(n_705),
.B(n_700),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_706),
.B(n_707),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_705),
.B(n_701),
.C(n_566),
.Y(n_710)
);

XOR2xp5_ASAP7_75t_L g711 ( 
.A(n_709),
.B(n_516),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_708),
.Y(n_712)
);

AOI31xp33_ASAP7_75t_L g713 ( 
.A1(n_710),
.A2(n_486),
.A3(n_524),
.B(n_560),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_709),
.Y(n_714)
);

OAI211xp5_ASAP7_75t_SL g715 ( 
.A1(n_710),
.A2(n_543),
.B(n_556),
.C(n_558),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_712),
.Y(n_716)
);

XNOR2xp5_ASAP7_75t_L g717 ( 
.A(n_711),
.B(n_579),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_714),
.B(n_524),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_713),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_715),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_714),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_721),
.A2(n_586),
.B1(n_585),
.B2(n_580),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_721),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_716),
.B(n_593),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_720),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_719),
.A2(n_614),
.B1(n_604),
.B2(n_586),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_723),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_725),
.A2(n_718),
.B1(n_717),
.B2(n_521),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_724),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_727),
.A2(n_722),
.B1(n_518),
.B2(n_485),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_730),
.A2(n_485),
.B1(n_560),
.B2(n_537),
.Y(n_732)
);

AO21x2_ASAP7_75t_L g733 ( 
.A1(n_728),
.A2(n_474),
.B(n_492),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_732),
.A2(n_729),
.B(n_492),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_733),
.A2(n_461),
.B(n_463),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_734),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_736),
.A2(n_731),
.B(n_735),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_737),
.A2(n_467),
.B(n_534),
.Y(n_738)
);

AOI21xp33_ASAP7_75t_SL g739 ( 
.A1(n_738),
.A2(n_467),
.B(n_534),
.Y(n_739)
);


endmodule