module real_aes_17916_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_884;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_0), .Y(n_200) );
AND2x4_ASAP7_75t_L g106 ( .A(n_1), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_2), .B(n_495), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_2), .B(n_496), .C(n_504), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_2), .B(n_504), .C(n_509), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_3), .Y(n_879) );
BUFx3_ASAP7_75t_L g266 ( .A(n_4), .Y(n_266) );
INVx1_ASAP7_75t_L g107 ( .A(n_5), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_6), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g113 ( .A(n_7), .B(n_23), .Y(n_113) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_8), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_9), .B(n_155), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_10), .B(n_155), .Y(n_538) );
INVx1_ASAP7_75t_L g885 ( .A(n_11), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_12), .B(n_181), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_13), .A2(n_84), .B1(n_151), .B2(n_155), .Y(n_154) );
OAI22x1_ASAP7_75t_L g496 ( .A1(n_14), .A2(n_28), .B1(n_497), .B2(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_14), .Y(n_498) );
OAI21x1_ASAP7_75t_L g144 ( .A1(n_15), .A2(n_39), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_16), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_17), .B(n_192), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_18), .Y(n_550) );
AO32x1_ASAP7_75t_L g142 ( .A1(n_19), .A2(n_143), .A3(n_146), .B1(n_157), .B2(n_161), .Y(n_142) );
AO32x2_ASAP7_75t_L g274 ( .A1(n_19), .A2(n_143), .A3(n_146), .B1(n_157), .B2(n_161), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_20), .B(n_575), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_21), .B(n_161), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_22), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_24), .A2(n_30), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_24), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_25), .A2(n_45), .B1(n_192), .B2(n_193), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_26), .A2(n_92), .B1(n_151), .B2(n_153), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_27), .B(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g497 ( .A(n_28), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_29), .Y(n_554) );
INVx1_ASAP7_75t_L g516 ( .A(n_30), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_31), .B(n_169), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_32), .A2(n_65), .B1(n_153), .B2(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_33), .B(n_155), .Y(n_590) );
INVx2_ASAP7_75t_L g128 ( .A(n_34), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_35), .B(n_156), .Y(n_599) );
BUFx3_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
INVx1_ASAP7_75t_L g120 ( .A(n_36), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_37), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_38), .B(n_557), .Y(n_605) );
AND2x2_ASAP7_75t_L g556 ( .A(n_40), .B(n_557), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_41), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_42), .B(n_201), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_43), .B(n_575), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_44), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_46), .B(n_626), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_47), .A2(n_78), .B1(n_169), .B2(n_201), .Y(n_252) );
OAI22xp5_ASAP7_75t_SL g512 ( .A1(n_48), .A2(n_513), .B1(n_514), .B2(n_517), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_48), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_49), .B(n_213), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_50), .A2(n_147), .B(n_198), .C(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_51), .A2(n_80), .B1(n_151), .B2(n_155), .Y(n_262) );
INVx1_ASAP7_75t_L g145 ( .A(n_52), .Y(n_145) );
AND2x4_ASAP7_75t_L g159 ( .A(n_53), .B(n_160), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_54), .A2(n_55), .B1(n_153), .B2(n_193), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_56), .B(n_161), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_57), .B(n_557), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_58), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_59), .B(n_153), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_60), .B(n_151), .Y(n_240) );
INVx1_ASAP7_75t_L g160 ( .A(n_61), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_62), .B(n_161), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_63), .A2(n_173), .B(n_198), .C(n_199), .Y(n_197) );
NAND3xp33_ASAP7_75t_L g246 ( .A(n_64), .B(n_151), .C(n_245), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_66), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_67), .B(n_161), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_68), .B(n_533), .Y(n_573) );
AND2x2_ASAP7_75t_L g203 ( .A(n_69), .B(n_204), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_70), .Y(n_216) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_71), .B(n_156), .C(n_192), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_72), .A2(n_95), .B1(n_155), .B2(n_201), .Y(n_254) );
INVx2_ASAP7_75t_L g149 ( .A(n_73), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_74), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_75), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_76), .B(n_196), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_77), .B(n_155), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_79), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_81), .B(n_229), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_82), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_83), .A2(n_91), .B1(n_575), .B2(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_85), .B(n_155), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_86), .B(n_245), .Y(n_244) );
NAND2xp33_ASAP7_75t_SL g566 ( .A(n_87), .B(n_242), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_88), .B(n_225), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_89), .A2(n_102), .B1(n_153), .B2(n_193), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_90), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_93), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_94), .B(n_181), .Y(n_180) );
NAND2xp33_ASAP7_75t_L g534 ( .A(n_96), .B(n_242), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_97), .B(n_557), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_98), .B(n_196), .C(n_242), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_99), .B(n_533), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_100), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_101), .B(n_575), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_114), .B(n_884), .Y(n_103) );
BUFx8_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_105), .Y(n_887) );
AND2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_L g883 ( .A(n_108), .Y(n_883) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_109), .Y(n_872) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g121 ( .A(n_110), .Y(n_121) );
NOR2x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g877 ( .A(n_112), .Y(n_877) );
INVx1_ASAP7_75t_L g122 ( .A(n_113), .Y(n_122) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_123), .Y(n_114) );
INVxp67_ASAP7_75t_L g499 ( .A(n_115), .Y(n_499) );
AOI211xp5_ASAP7_75t_L g500 ( .A1(n_115), .A2(n_132), .B(n_496), .C(n_501), .Y(n_500) );
NOR2xp67_ASAP7_75t_SL g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx4_ASAP7_75t_L g495 ( .A(n_118), .Y(n_495) );
AND3x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .C(n_122), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g507 ( .A(n_120), .Y(n_507) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_121), .Y(n_519) );
AND2x6_ASAP7_75t_SL g505 ( .A(n_122), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_122), .B(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_510), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g875 ( .A(n_128), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_128), .B(n_883), .Y(n_882) );
OAI21xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_500), .B(n_502), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_493), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_131), .A2(n_132), .B1(n_503), .B2(n_508), .Y(n_502) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OA22x2_ASAP7_75t_L g518 ( .A1(n_133), .A2(n_519), .B1(n_520), .B2(n_871), .Y(n_518) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_380), .Y(n_133) );
AND4x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_289), .C(n_327), .D(n_365), .Y(n_134) );
NOR2x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_267), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_206), .B(n_217), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_162), .Y(n_138) );
NAND2xp5_ASAP7_75t_R g338 ( .A(n_139), .B(n_286), .Y(n_338) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g439 ( .A(n_141), .B(n_317), .Y(n_439) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g208 ( .A(n_142), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g300 ( .A(n_142), .Y(n_300) );
AND2x2_ASAP7_75t_L g314 ( .A(n_142), .B(n_209), .Y(n_314) );
INVx4_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx2_ASAP7_75t_SL g165 ( .A(n_143), .Y(n_165) );
BUFx3_ASAP7_75t_L g210 ( .A(n_143), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_143), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_143), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_SL g539 ( .A(n_143), .B(n_233), .Y(n_539) );
INVx1_ASAP7_75t_SL g559 ( .A(n_143), .Y(n_559) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B1(n_154), .B2(n_156), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_L g222 ( .A1(n_147), .A2(n_223), .B(n_224), .C(n_226), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_147), .A2(n_532), .B(n_534), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_147), .A2(n_565), .B(n_566), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_147), .A2(n_573), .B(n_574), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_147), .A2(n_589), .B(n_590), .Y(n_588) );
BUFx4f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g245 ( .A(n_148), .Y(n_245) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx8_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx2_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
INVx1_ASAP7_75t_L g196 ( .A(n_149), .Y(n_196) );
INVx2_ASAP7_75t_SL g169 ( .A(n_151), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_151), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_152), .Y(n_153) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx1_ASAP7_75t_L g198 ( .A(n_152), .Y(n_198) );
INVx1_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
INVx1_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_152), .Y(n_242) );
INVx3_ASAP7_75t_L g533 ( .A(n_152), .Y(n_533) );
INVx1_ASAP7_75t_L g576 ( .A(n_152), .Y(n_576) );
INVx2_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g553 ( .A1(n_153), .A2(n_533), .B1(n_554), .B2(n_555), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_153), .A2(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_L g612 ( .A(n_153), .Y(n_612) );
INVx3_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_155), .A2(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g604 ( .A(n_155), .Y(n_604) );
INVx6_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_156), .A2(n_240), .B(n_241), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_156), .A2(n_179), .B1(n_262), .B2(n_263), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_156), .A2(n_592), .B(n_593), .Y(n_591) );
O2A1O1Ixp5_ASAP7_75t_L g620 ( .A1(n_156), .A2(n_224), .B(n_621), .C(n_622), .Y(n_620) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_157), .A2(n_167), .B(n_175), .Y(n_166) );
INVx2_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_SL g255 ( .A(n_158), .Y(n_255) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
AO31x2_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_210), .A3(n_211), .B(n_215), .Y(n_209) );
BUFx10_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
BUFx10_ASAP7_75t_L g546 ( .A(n_159), .Y(n_546) );
INVx2_ASAP7_75t_L g260 ( .A(n_161), .Y(n_260) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_184), .Y(n_162) );
BUFx2_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
AND2x2_ASAP7_75t_L g272 ( .A(n_163), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g287 ( .A(n_163), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_163), .B(n_209), .Y(n_304) );
INVx3_ASAP7_75t_L g317 ( .A(n_163), .Y(n_317) );
AND2x2_ASAP7_75t_L g352 ( .A(n_163), .B(n_274), .Y(n_352) );
INVx2_ASAP7_75t_L g364 ( .A(n_163), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_163), .Y(n_368) );
INVxp67_ASAP7_75t_L g405 ( .A(n_163), .Y(n_405) );
OR2x2_ASAP7_75t_L g418 ( .A(n_163), .B(n_301), .Y(n_418) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_180), .Y(n_164) );
AOI21x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B(n_172), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_171), .A2(n_244), .B(n_246), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_172), .A2(n_179), .B1(n_212), .B2(n_214), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_172), .A2(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g552 ( .A(n_173), .Y(n_552) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g230 ( .A(n_174), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_179), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_179), .A2(n_252), .B1(n_253), .B2(n_254), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_179), .A2(n_552), .B1(n_611), .B2(n_613), .Y(n_610) );
INVx2_ASAP7_75t_L g187 ( .A(n_181), .Y(n_187) );
NOR2xp67_ASAP7_75t_SL g544 ( .A(n_181), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AO31x2_ASAP7_75t_L g609 ( .A1(n_182), .A2(n_546), .A3(n_610), .B(n_614), .Y(n_609) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g205 ( .A(n_183), .Y(n_205) );
INVx2_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g270 ( .A(n_185), .Y(n_270) );
INVx1_ASAP7_75t_L g357 ( .A(n_185), .Y(n_357) );
AND2x2_ASAP7_75t_L g372 ( .A(n_185), .B(n_209), .Y(n_372) );
INVx1_ASAP7_75t_L g387 ( .A(n_185), .Y(n_387) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g301 ( .A(n_186), .Y(n_301) );
AOI21x1_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_203), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_197), .B(n_202), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_190), .B(n_195), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B1(n_193), .B2(n_194), .Y(n_190) );
INVx2_ASAP7_75t_L g213 ( .A(n_192), .Y(n_213) );
INVx1_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
AOI21x1_ASAP7_75t_L g601 ( .A1(n_195), .A2(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_SL g253 ( .A(n_196), .Y(n_253) );
INVx1_ASAP7_75t_L g537 ( .A(n_198), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_205), .B(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_205), .B(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_206), .A2(n_476), .B1(n_478), .B2(n_480), .Y(n_475) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_207), .B(n_356), .Y(n_433) );
BUFx2_ASAP7_75t_L g447 ( .A(n_207), .Y(n_447) );
AND2x2_ASAP7_75t_L g465 ( .A(n_207), .B(n_321), .Y(n_465) );
INVx2_ASAP7_75t_L g347 ( .A(n_208), .Y(n_347) );
OR2x2_ASAP7_75t_L g363 ( .A(n_208), .B(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g271 ( .A(n_209), .Y(n_271) );
AND2x2_ASAP7_75t_L g356 ( .A(n_209), .B(n_357), .Y(n_356) );
AO31x2_ASAP7_75t_L g250 ( .A1(n_210), .A2(n_251), .A3(n_255), .B(n_256), .Y(n_250) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_248), .Y(n_217) );
OR2x2_ASAP7_75t_L g412 ( .A(n_218), .B(n_369), .Y(n_412) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_235), .Y(n_218) );
AND2x2_ASAP7_75t_L g283 ( .A(n_219), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g324 ( .A(n_219), .Y(n_324) );
INVx2_ASAP7_75t_SL g332 ( .A(n_219), .Y(n_332) );
BUFx2_ASAP7_75t_L g344 ( .A(n_219), .Y(n_344) );
OR2x2_ASAP7_75t_L g432 ( .A(n_219), .B(n_250), .Y(n_432) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_234), .Y(n_219) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_220), .A2(n_221), .B(n_234), .Y(n_297) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_220), .A2(n_587), .B(n_594), .Y(n_586) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_220), .A2(n_597), .B(n_605), .Y(n_596) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_220), .A2(n_587), .B(n_594), .Y(n_651) );
OA21x2_ASAP7_75t_L g654 ( .A1(n_220), .A2(n_597), .B(n_605), .Y(n_654) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_227), .B(n_233), .Y(n_221) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_230), .B1(n_231), .B2(n_232), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_229), .A2(n_624), .B(n_625), .Y(n_623) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_230), .A2(n_536), .B1(n_537), .B2(n_538), .Y(n_535) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_233), .A2(n_239), .B(n_243), .Y(n_238) );
AOI31xp67_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_260), .A3(n_261), .B(n_264), .Y(n_259) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_233), .A2(n_561), .B(n_564), .Y(n_560) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_233), .A2(n_572), .B(n_577), .Y(n_571) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_233), .A2(n_588), .B(n_591), .Y(n_587) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_233), .A2(n_598), .B(n_601), .Y(n_597) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_233), .A2(n_620), .B(n_623), .Y(n_619) );
AND2x2_ASAP7_75t_L g276 ( .A(n_235), .B(n_258), .Y(n_276) );
AND2x2_ASAP7_75t_L g312 ( .A(n_235), .B(n_297), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_238), .B(n_247), .Y(n_235) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_236), .A2(n_238), .B(n_247), .Y(n_282) );
OAI21xp33_ASAP7_75t_SL g570 ( .A1(n_236), .A2(n_571), .B(n_580), .Y(n_570) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_236), .A2(n_619), .B(n_627), .Y(n_618) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_236), .A2(n_571), .B(n_580), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_236), .A2(n_619), .B(n_627), .Y(n_702) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g557 ( .A(n_237), .Y(n_557) );
INVx2_ASAP7_75t_L g626 ( .A(n_242), .Y(n_626) );
INVx1_ASAP7_75t_L g350 ( .A(n_248), .Y(n_350) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_249), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g456 ( .A(n_249), .B(n_436), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_249), .B(n_279), .Y(n_480) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_258), .Y(n_249) );
INVx1_ASAP7_75t_L g284 ( .A(n_250), .Y(n_284) );
INVx2_ASAP7_75t_L g294 ( .A(n_250), .Y(n_294) );
AND2x2_ASAP7_75t_L g308 ( .A(n_250), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g323 ( .A(n_250), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g337 ( .A(n_250), .B(n_297), .Y(n_337) );
OR2x2_ASAP7_75t_L g369 ( .A(n_250), .B(n_309), .Y(n_369) );
INVx1_ASAP7_75t_L g453 ( .A(n_250), .Y(n_453) );
AND2x2_ASAP7_75t_L g296 ( .A(n_258), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g334 ( .A(n_258), .Y(n_334) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_266), .Y(n_265) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_275), .B1(n_277), .B2(n_285), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g414 ( .A(n_270), .Y(n_414) );
INVx1_ASAP7_75t_L g288 ( .A(n_271), .Y(n_288) );
AND2x4_ASAP7_75t_L g321 ( .A(n_271), .B(n_274), .Y(n_321) );
AND2x2_ASAP7_75t_L g430 ( .A(n_271), .B(n_301), .Y(n_430) );
AND2x2_ASAP7_75t_L g482 ( .A(n_272), .B(n_356), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_272), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g336 ( .A(n_276), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g469 ( .A(n_276), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_283), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_279), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g388 ( .A(n_279), .Y(n_388) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g454 ( .A(n_280), .Y(n_454) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g341 ( .A(n_281), .Y(n_341) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g326 ( .A(n_282), .B(n_310), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_283), .B(n_325), .Y(n_441) );
AND2x2_ASAP7_75t_L g333 ( .A(n_284), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g473 ( .A(n_288), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_298), .B1(n_305), .B2(n_313), .C(n_318), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
AND2x2_ASAP7_75t_L g391 ( .A(n_292), .B(n_312), .Y(n_391) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_293), .B(n_312), .Y(n_360) );
OR2x2_ASAP7_75t_L g375 ( .A(n_293), .B(n_326), .Y(n_375) );
INVx2_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g451 ( .A(n_296), .Y(n_451) );
INVx1_ASAP7_75t_L g411 ( .A(n_297), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
AND2x2_ASAP7_75t_L g471 ( .A(n_299), .B(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g425 ( .A(n_300), .B(n_387), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_301), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
INVx1_ASAP7_75t_L g398 ( .A(n_301), .Y(n_398) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI21xp33_ASAP7_75t_L g366 ( .A1(n_306), .A2(n_332), .B(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_311), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g361 ( .A(n_308), .B(n_344), .Y(n_361) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_308), .Y(n_401) );
AND2x2_ASAP7_75t_L g485 ( .A(n_308), .B(n_422), .Y(n_485) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g492 ( .A(n_311), .B(n_409), .Y(n_492) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_SL g393 ( .A(n_314), .Y(n_393) );
AND2x2_ASAP7_75t_L g397 ( .A(n_314), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g457 ( .A(n_314), .B(n_317), .Y(n_457) );
AND2x2_ASAP7_75t_L g479 ( .A(n_314), .B(n_404), .Y(n_479) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g376 ( .A(n_317), .B(n_321), .Y(n_376) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g370 ( .A(n_321), .B(n_346), .Y(n_370) );
AND2x2_ASAP7_75t_L g403 ( .A(n_321), .B(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g420 ( .A(n_321), .Y(n_420) );
INVx1_ASAP7_75t_L g489 ( .A(n_322), .Y(n_489) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
AND2x4_ASAP7_75t_L g353 ( .A(n_323), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g395 ( .A(n_325), .B(n_344), .Y(n_395) );
AND2x2_ASAP7_75t_L g421 ( .A(n_325), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g431 ( .A(n_326), .B(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_348), .Y(n_327) );
A2O1A1Ixp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_335), .B(n_338), .C(n_339), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_331), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_332), .B(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_332), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_333), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g354 ( .A(n_334), .B(n_341), .Y(n_354) );
INVx1_ASAP7_75t_L g409 ( .A(n_334), .Y(n_409) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B(n_345), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_341), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g422 ( .A(n_344), .Y(n_422) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AND2x4_ASAP7_75t_L g446 ( .A(n_347), .B(n_414), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_358), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B(n_353), .C(n_355), .Y(n_349) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g413 ( .A(n_352), .B(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_361), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_364), .Y(n_373) );
OR2x2_ASAP7_75t_L g392 ( .A(n_364), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g474 ( .A(n_364), .Y(n_474) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B1(n_371), .B2(n_374), .C1(n_376), .C2(n_377), .Y(n_365) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_367), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_368), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g379 ( .A(n_369), .Y(n_379) );
INVx1_ASAP7_75t_L g477 ( .A(n_369), .Y(n_477) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_372), .B(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g455 ( .A(n_372), .Y(n_455) );
AND2x4_ASAP7_75t_L g462 ( .A(n_372), .B(n_439), .Y(n_462) );
INVx2_ASAP7_75t_L g491 ( .A(n_372), .Y(n_491) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_375), .A2(n_428), .B1(n_431), .B2(n_433), .Y(n_427) );
AOI211xp5_ASAP7_75t_L g481 ( .A1(n_377), .A2(n_482), .B(n_483), .C(n_487), .Y(n_481) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NOR2xp67_ASAP7_75t_SL g380 ( .A(n_381), .B(n_442), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_399), .C(n_406), .D(n_426), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_388), .B(n_389), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B1(n_394), .B2(n_396), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_393), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_394), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g404 ( .A(n_398), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_413), .B1(n_415), .B2(n_421), .C(n_423), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_412), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_408), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g461 ( .A(n_409), .B(n_436), .Y(n_461) );
INVx2_ASAP7_75t_L g436 ( .A(n_410), .Y(n_436) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
NAND2x1_ASAP7_75t_SL g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g486 ( .A(n_417), .Y(n_486) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g488 ( .A(n_425), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_434), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_440), .B2(n_441), .Y(n_434) );
AND2x2_ASAP7_75t_L g467 ( .A(n_436), .B(n_453), .Y(n_467) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g448 ( .A(n_441), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_458), .C(n_481), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_448), .B1(n_449), .B2(n_455), .C1(n_456), .C2(n_457), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AOI211xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_463), .C(n_475), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B1(n_468), .B2(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_490), .B2(n_492), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_499), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_494), .Y(n_501) );
INVx1_ASAP7_75t_L g509 ( .A(n_496), .Y(n_509) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI21xp33_ASAP7_75t_SL g510 ( .A1(n_511), .A2(n_873), .B(n_878), .Y(n_510) );
XNOR2x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_751), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_659), .C(n_710), .Y(n_521) );
OAI211xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_581), .B(n_628), .C(n_646), .Y(n_522) );
NAND3x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_540), .C(n_568), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g719 ( .A(n_525), .B(n_698), .Y(n_719) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND3x2_ASAP7_75t_L g639 ( .A(n_526), .B(n_640), .C(n_644), .Y(n_639) );
AND2x2_ASAP7_75t_L g674 ( .A(n_526), .B(n_658), .Y(n_674) );
AND2x2_ASAP7_75t_L g680 ( .A(n_526), .B(n_676), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g821 ( .A(n_526), .B(n_644), .Y(n_821) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g723 ( .A(n_527), .B(n_644), .Y(n_723) );
AND2x2_ASAP7_75t_L g734 ( .A(n_527), .B(n_688), .Y(n_734) );
BUFx2_ASAP7_75t_L g740 ( .A(n_527), .Y(n_740) );
NAND2x1_ASAP7_75t_L g756 ( .A(n_527), .B(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g762 ( .A(n_527), .B(n_763), .Y(n_762) );
INVx4_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g656 ( .A(n_528), .Y(n_656) );
AND2x2_ASAP7_75t_L g687 ( .A(n_528), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g707 ( .A(n_528), .B(n_643), .Y(n_707) );
INVx1_ASAP7_75t_L g778 ( .A(n_528), .Y(n_778) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_535), .B(n_539), .Y(n_530) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x6_ASAP7_75t_L g755 ( .A(n_541), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g657 ( .A(n_542), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_542), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_558), .Y(n_542) );
INVx2_ASAP7_75t_L g645 ( .A(n_543), .Y(n_645) );
INVx1_ASAP7_75t_L g699 ( .A(n_543), .Y(n_699) );
AOI21x1_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .B(n_556), .Y(n_543) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g643 ( .A(n_558), .Y(n_643) );
INVx2_ASAP7_75t_L g677 ( .A(n_558), .Y(n_677) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_567), .Y(n_558) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_569), .A2(n_859), .B(n_863), .Y(n_858) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g698 ( .A(n_570), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_606), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g854 ( .A(n_583), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp67_ASAP7_75t_L g584 ( .A(n_585), .B(n_595), .Y(n_584) );
INVx3_ASAP7_75t_L g636 ( .A(n_585), .Y(n_636) );
AND2x2_ASAP7_75t_L g783 ( .A(n_585), .B(n_596), .Y(n_783) );
BUFx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g672 ( .A(n_586), .Y(n_672) );
AND2x4_ASAP7_75t_L g637 ( .A(n_595), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g696 ( .A(n_596), .Y(n_696) );
AND2x2_ASAP7_75t_L g713 ( .A(n_596), .B(n_609), .Y(n_713) );
AND2x2_ASAP7_75t_L g825 ( .A(n_596), .B(n_702), .Y(n_825) );
AND2x2_ASAP7_75t_L g847 ( .A(n_596), .B(n_617), .Y(n_847) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_616), .Y(n_607) );
INVx1_ASAP7_75t_L g667 ( .A(n_608), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_608), .B(n_857), .Y(n_856) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g638 ( .A(n_609), .Y(n_638) );
OR2x2_ASAP7_75t_L g653 ( .A(n_609), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g671 ( .A(n_609), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g725 ( .A(n_609), .B(n_651), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_609), .B(n_654), .Y(n_767) );
OR2x2_ASAP7_75t_L g837 ( .A(n_609), .B(n_651), .Y(n_837) );
INVx1_ASAP7_75t_L g665 ( .A(n_616), .Y(n_665) );
AND2x4_ASAP7_75t_L g683 ( .A(n_616), .B(n_637), .Y(n_683) );
AND2x2_ASAP7_75t_L g829 ( .A(n_616), .B(n_671), .Y(n_829) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx3_ASAP7_75t_L g631 ( .A(n_617), .Y(n_631) );
AND2x2_ASAP7_75t_L g691 ( .A(n_617), .B(n_650), .Y(n_691) );
INVx1_ASAP7_75t_L g744 ( .A(n_617), .Y(n_744) );
INVxp67_ASAP7_75t_SL g782 ( .A(n_617), .Y(n_782) );
AND2x2_ASAP7_75t_L g785 ( .A(n_617), .B(n_654), .Y(n_785) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_617), .Y(n_795) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_632), .B(n_639), .Y(n_628) );
AND2x2_ASAP7_75t_L g827 ( .A(n_629), .B(n_732), .Y(n_827) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g694 ( .A(n_630), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_630), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_631), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g774 ( .A(n_631), .B(n_637), .Y(n_774) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_636), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g772 ( .A(n_636), .B(n_713), .Y(n_772) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_636), .Y(n_803) );
INVx2_ASAP7_75t_L g737 ( .A(n_637), .Y(n_737) );
AND2x2_ASAP7_75t_L g866 ( .A(n_638), .B(n_651), .Y(n_866) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_639), .A2(n_721), .B1(n_722), .B2(n_724), .C(n_726), .Y(n_720) );
AND2x2_ASAP7_75t_L g661 ( .A(n_640), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g722 ( .A(n_640), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx2_ASAP7_75t_L g658 ( .A(n_641), .Y(n_658) );
OR2x2_ASAP7_75t_L g791 ( .A(n_641), .B(n_676), .Y(n_791) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g688 ( .A(n_642), .Y(n_688) );
INVxp67_ASAP7_75t_L g718 ( .A(n_643), .Y(n_718) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g662 ( .A(n_645), .Y(n_662) );
AND2x2_ASAP7_75t_L g675 ( .A(n_645), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g682 ( .A(n_645), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_655), .Y(n_646) );
AND2x2_ASAP7_75t_L g805 ( .A(n_647), .B(n_806), .Y(n_805) );
AND2x4_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g732 ( .A(n_649), .B(n_713), .Y(n_732) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_649), .Y(n_862) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g690 ( .A(n_652), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g840 ( .A(n_652), .Y(n_840) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g728 ( .A(n_653), .Y(n_728) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_653), .Y(n_802) );
AND2x2_ASAP7_75t_L g701 ( .A(n_654), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_655), .B(n_827), .Y(n_826) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g697 ( .A(n_656), .B(n_698), .Y(n_697) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_657), .A2(n_679), .B(n_683), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_678), .C(n_684), .D(n_692), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_663), .B(n_668), .Y(n_660) );
INVx2_ASAP7_75t_L g749 ( .A(n_662), .Y(n_749) );
AND2x2_ASAP7_75t_L g760 ( .A(n_662), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g770 ( .A(n_662), .B(n_687), .Y(n_770) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g846 ( .A(n_667), .B(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI33xp33_ASAP7_75t_L g816 ( .A1(n_670), .A2(n_707), .A3(n_817), .B1(n_819), .B2(n_822), .B3(n_823), .Y(n_816) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g849 ( .A(n_671), .B(n_701), .Y(n_849) );
BUFx2_ASAP7_75t_L g704 ( .A(n_672), .Y(n_704) );
AND2x4_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_675), .B(n_687), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_676), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_677), .Y(n_730) );
INVx1_ASAP7_75t_L g763 ( .A(n_677), .Y(n_763) );
AND2x2_ASAP7_75t_L g777 ( .A(n_677), .B(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AND2x2_ASAP7_75t_L g748 ( .A(n_680), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g800 ( .A(n_680), .Y(n_800) );
INVx1_ASAP7_75t_L g810 ( .A(n_681), .Y(n_810) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g686 ( .A(n_682), .Y(n_686) );
INVx1_ASAP7_75t_L g792 ( .A(n_682), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_689), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
OR2x2_ASAP7_75t_L g775 ( .A(n_686), .B(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g746 ( .A(n_687), .B(n_730), .Y(n_746) );
AND2x2_ASAP7_75t_L g709 ( .A(n_688), .B(n_699), .Y(n_709) );
INVx2_ASAP7_75t_L g757 ( .A(n_688), .Y(n_757) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g750 ( .A(n_691), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_697), .B1(n_700), .B2(n_705), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_695), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_697), .A2(n_780), .B1(n_784), .B2(n_786), .C(n_788), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_698), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g834 ( .A(n_698), .Y(n_834) );
AND2x2_ASAP7_75t_L g853 ( .A(n_698), .B(n_777), .Y(n_853) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g822 ( .A(n_701), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_701), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g808 ( .A(n_702), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_703), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g796 ( .A(n_703), .B(n_737), .Y(n_796) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_705), .A2(n_851), .B1(n_853), .B2(n_854), .Y(n_850) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
OR2x2_ASAP7_75t_L g867 ( .A(n_708), .B(n_762), .Y(n_867) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g815 ( .A(n_709), .B(n_777), .Y(n_815) );
OAI211xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .B(n_720), .C(n_735), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_713), .Y(n_721) );
AND2x2_ASAP7_75t_L g794 ( .A(n_713), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2x1p5_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g787 ( .A(n_719), .Y(n_787) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_725), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g784 ( .A(n_725), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g818 ( .A(n_725), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_725), .B(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B1(n_731), .B2(n_733), .Y(n_726) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI21xp33_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_738), .B(n_741), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B1(n_747), .B2(n_750), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_743), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI211xp5_ASAP7_75t_SL g828 ( .A1(n_746), .A2(n_829), .B(n_830), .C(n_838), .Y(n_828) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g843 ( .A(n_749), .B(n_777), .Y(n_843) );
NOR3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_811), .C(n_841), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_779), .C(n_799), .Y(n_752) );
O2A1O1Ixp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_758), .B(n_764), .C(n_768), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI22xp33_ASAP7_75t_SL g830 ( .A1(n_756), .A2(n_831), .B1(n_833), .B2(n_835), .Y(n_830) );
INVx1_ASAP7_75t_SL g820 ( .A(n_757), .Y(n_820) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g833 ( .A(n_762), .B(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B1(n_773), .B2(n_775), .Y(n_768) );
NAND2xp33_ASAP7_75t_SL g786 ( .A(n_769), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g852 ( .A(n_774), .Y(n_852) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g806 ( .A(n_777), .B(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_781), .B(n_815), .Y(n_814) );
AND2x4_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVx1_ASAP7_75t_L g857 ( .A(n_782), .Y(n_857) );
INVx1_ASAP7_75t_L g832 ( .A(n_785), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_793), .B1(n_796), .B2(n_797), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2x1p5_ASAP7_75t_SL g790 ( .A(n_791), .B(n_792), .Y(n_790) );
INVx1_ASAP7_75t_L g798 ( .A(n_791), .Y(n_798) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
BUFx2_ASAP7_75t_L g804 ( .A(n_795), .Y(n_804) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B(n_805), .C(n_809), .Y(n_799) );
NOR3x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .C(n_804), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_806), .B(n_861), .Y(n_860) );
AND2x2_ASAP7_75t_L g865 ( .A(n_807), .B(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND3xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_826), .C(n_828), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_816), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
BUFx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NOR2xp67_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g870 ( .A(n_839), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_850), .C(n_858), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVxp67_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVxp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVxp67_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVxp67_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_867), .B1(n_868), .B2(n_869), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx4_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
AND2x6_ASAP7_75t_SL g874 ( .A(n_875), .B(n_876), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
INVx5_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
BUFx10_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_887), .Y(n_886) );
endmodule