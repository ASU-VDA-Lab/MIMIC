module fake_jpeg_25790_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_57),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_1),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_2),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_2),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_74),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_19),
.B(n_2),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_71),
.Y(n_77)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_34),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_29),
.B1(n_25),
.B2(n_16),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_82),
.B1(n_86),
.B2(n_33),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_29),
.B1(n_25),
.B2(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_39),
.B1(n_35),
.B2(n_30),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_84),
.A2(n_17),
.B1(n_33),
.B2(n_27),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_29),
.B1(n_25),
.B2(n_16),
.Y(n_86)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_94),
.B(n_97),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_35),
.Y(n_97)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_41),
.B(n_21),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_50),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_123),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_42),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_121),
.B(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_48),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_21),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_125),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_51),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_128),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_28),
.B1(n_22),
.B2(n_24),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_30),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_78),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_134),
.Y(n_170)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_72),
.B1(n_45),
.B2(n_22),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_63),
.A3(n_24),
.B1(n_33),
.B2(n_28),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_77),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_24),
.B(n_17),
.C(n_22),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_75),
.B(n_31),
.Y(n_183)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_60),
.C(n_53),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_151),
.C(n_87),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_34),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_145),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_20),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_149),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_28),
.B1(n_27),
.B2(n_85),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_34),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_2),
.C(n_3),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_157),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_98),
.B(n_27),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_91),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_46),
.C(n_47),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_20),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_155),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_81),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_162),
.A2(n_180),
.B1(n_158),
.B2(n_129),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_85),
.B1(n_87),
.B2(n_118),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_184),
.B1(n_155),
.B2(n_157),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_109),
.B1(n_93),
.B2(n_100),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_56),
.B(n_55),
.Y(n_167)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_167),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_179),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_96),
.C(n_111),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_195),
.C(n_138),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_121),
.B(n_143),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_118),
.B1(n_117),
.B2(n_106),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_188),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_185),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_SL g240 ( 
.A1(n_183),
.A2(n_9),
.B(n_10),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_123),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_108),
.B1(n_100),
.B2(n_66),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_134),
.B1(n_148),
.B2(n_156),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_122),
.A2(n_31),
.B1(n_61),
.B2(n_54),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_126),
.B(n_3),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_6),
.Y(n_229)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_207),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_152),
.B1(n_161),
.B2(n_122),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_203),
.A2(n_204),
.B1(n_187),
.B2(n_188),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_126),
.B1(n_147),
.B2(n_135),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_206),
.A2(n_208),
.B1(n_215),
.B2(n_223),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_199),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_147),
.B1(n_154),
.B2(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_212),
.Y(n_249)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_139),
.B1(n_159),
.B2(n_151),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_224),
.B1(n_240),
.B2(n_184),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_217),
.B(n_219),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_222),
.Y(n_263)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_167),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_140),
.C(n_127),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_168),
.C(n_172),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_131),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_158),
.B1(n_119),
.B2(n_150),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_156),
.B(n_142),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_227),
.B(n_232),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_176),
.A2(n_156),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_226),
.A2(n_236),
.B1(n_165),
.B2(n_171),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_3),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_192),
.Y(n_230)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_6),
.B(n_7),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g233 ( 
.A1(n_167),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_7),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_239),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_8),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_210),
.B1(n_231),
.B2(n_207),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_253),
.B1(n_257),
.B2(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_251),
.C(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_172),
.C(n_189),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_252),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_231),
.B1(n_213),
.B2(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_189),
.C(n_191),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_200),
.B1(n_163),
.B2(n_189),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_270),
.Y(n_288)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_204),
.A2(n_200),
.B1(n_167),
.B2(n_177),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_214),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_264),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_226),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_265),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_215),
.A2(n_194),
.B1(n_178),
.B2(n_173),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_267),
.A2(n_269),
.B1(n_233),
.B2(n_227),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_183),
.B1(n_173),
.B2(n_178),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_199),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_228),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_208),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_232),
.B(n_225),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_279),
.B(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_282),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_221),
.C(n_218),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_281),
.C(n_241),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_205),
.B(n_225),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_239),
.C(n_206),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_296),
.Y(n_304)
);

HAxp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_199),
.CON(n_285),
.SN(n_285)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_285),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_235),
.Y(n_286)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_232),
.B(n_259),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_205),
.B(n_234),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_299),
.B1(n_257),
.B2(n_269),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_195),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_293),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_186),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_242),
.A2(n_236),
.B(n_233),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_298),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_247),
.A2(n_227),
.B1(n_171),
.B2(n_174),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_256),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_305),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_246),
.Y(n_305)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_246),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_311),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_247),
.B1(n_252),
.B2(n_265),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_308),
.A2(n_288),
.B1(n_298),
.B2(n_301),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_271),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_261),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_314),
.C(n_321),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_288),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_323),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_286),
.Y(n_318)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_284),
.A2(n_268),
.B1(n_254),
.B2(n_249),
.Y(n_319)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_268),
.C(n_243),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_243),
.C(n_250),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_281),
.C(n_291),
.Y(n_330)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_287),
.Y(n_323)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_294),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_332),
.C(n_333),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_293),
.C(n_280),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_280),
.C(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_315),
.Y(n_335)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_325),
.A2(n_294),
.B1(n_277),
.B2(n_295),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_336),
.B(n_343),
.C(n_347),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_300),
.C(n_283),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_322),
.C(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_308),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_340),
.B(n_342),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_255),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_295),
.B1(n_301),
.B2(n_290),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_344),
.A2(n_312),
.B1(n_299),
.B2(n_260),
.Y(n_363)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_346),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_307),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_354),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_335),
.A2(n_288),
.B1(n_316),
.B2(n_310),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_347),
.Y(n_371)
);

OAI322xp33_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_320),
.A3(n_303),
.B1(n_313),
.B2(n_282),
.C1(n_317),
.C2(n_250),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_345),
.A2(n_309),
.B(n_289),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_356),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_290),
.B(n_275),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_296),
.B1(n_255),
.B2(n_297),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_357),
.A2(n_363),
.B1(n_258),
.B2(n_237),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_338),
.C(n_330),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_202),
.Y(n_359)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_337),
.B(n_333),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_362),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_329),
.C(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_365),
.B(n_366),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_329),
.C(n_338),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_369),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_328),
.C(n_331),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_344),
.C(n_326),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_374),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_355),
.B(n_348),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_372),
.A2(n_353),
.B1(n_348),
.B2(n_352),
.Y(n_381)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_356),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_326),
.B1(n_174),
.B2(n_175),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_378),
.A2(n_382),
.B(n_370),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_371),
.A2(n_373),
.B1(n_360),
.B2(n_361),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_383),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_381),
.B(n_385),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_376),
.A2(n_361),
.B(n_352),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_367),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_351),
.B(n_11),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_365),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_384),
.B(n_366),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_392),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_391),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_394),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_175),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_10),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_386),
.A2(n_11),
.B(n_12),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_378),
.C(n_377),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_401),
.B(n_402),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_381),
.C(n_385),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_397),
.A2(n_395),
.B(n_388),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_403),
.A2(n_405),
.B(n_400),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_11),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_406),
.A2(n_407),
.B(n_11),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_404),
.A2(n_398),
.B(n_12),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_14),
.B(n_15),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_15),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_15),
.Y(n_411)
);


endmodule