module fake_jpeg_25242_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_0),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_3),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_70),
.B(n_64),
.C(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_57),
.B1(n_68),
.B2(n_65),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_69),
.B1(n_67),
.B2(n_61),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_57),
.B1(n_68),
.B2(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_91),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_53),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_62),
.B1(n_53),
.B2(n_66),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_69),
.B1(n_67),
.B2(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_66),
.B1(n_50),
.B2(n_47),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_80),
.B1(n_82),
.B2(n_52),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_55),
.B1(n_54),
.B2(n_59),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_98),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_51),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_102),
.B(n_6),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_90),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_92),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_73),
.B1(n_61),
.B2(n_7),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_113),
.B1(n_8),
.B2(n_9),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_93),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_125),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_105),
.C(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_106),
.C(n_8),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_122),
.B(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_123),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_102),
.B1(n_97),
.B2(n_31),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_110),
.B1(n_115),
.B2(n_11),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_7),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_114),
.B(n_10),
.Y(n_127)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_130),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_135),
.Y(n_140)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_134),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_133),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_132),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_139),
.C(n_10),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_110),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_32),
.B(n_44),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_143),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_129),
.C(n_34),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_128),
.B1(n_127),
.B2(n_136),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_149),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_147),
.B1(n_146),
.B2(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_145),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_150),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_140),
.A3(n_30),
.B1(n_35),
.B2(n_14),
.C1(n_15),
.C2(n_18),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_46),
.A3(n_36),
.B1(n_37),
.B2(n_20),
.C1(n_24),
.C2(n_28),
.Y(n_157)
);

AOI31xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_39),
.A3(n_40),
.B(n_42),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_43),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_11),
.Y(n_160)
);


endmodule