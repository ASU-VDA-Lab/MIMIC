module fake_jpeg_31955_n_371 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_371);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_72),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_24),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_52),
.Y(n_122)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_32),
.B1(n_20),
.B2(n_31),
.Y(n_76)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_70),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_71),
.B(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_75),
.B(n_82),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_76),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_38),
.B1(n_37),
.B2(n_21),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_91),
.B1(n_116),
.B2(n_64),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_40),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_87),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_92),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_85),
.B(n_86),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_34),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_99),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_27),
.B1(n_26),
.B2(n_33),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_95),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_15),
.B(n_18),
.C(n_29),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_73),
.B(n_96),
.C(n_78),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_15),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_19),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_102),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_44),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_68),
.B(n_0),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_5),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_44),
.B(n_23),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_63),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_66),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_66),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_120),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_23),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_124),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

HB1xp67_ASAP7_75t_SL g186 ( 
.A(n_131),
.Y(n_186)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_70),
.B1(n_61),
.B2(n_33),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_144),
.B1(n_119),
.B2(n_114),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_76),
.A2(n_1),
.B(n_2),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_136),
.A2(n_138),
.B(n_164),
.Y(n_215)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_27),
.B(n_19),
.C(n_16),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_29),
.B1(n_18),
.B2(n_16),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_143),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_16),
.B1(n_10),
.B2(n_11),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_16),
.B1(n_9),
.B2(n_12),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_147),
.B1(n_156),
.B2(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_83),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_160),
.Y(n_191)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_161),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_93),
.A2(n_9),
.B1(n_13),
.B2(n_7),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_7),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_154),
.B(n_168),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_107),
.A2(n_96),
.B1(n_74),
.B2(n_106),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_98),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_161),
.C(n_129),
.Y(n_177)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_171),
.Y(n_196)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_79),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_174),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_175),
.A2(n_201),
.B1(n_171),
.B2(n_137),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_177),
.B(n_159),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_182),
.B1(n_185),
.B2(n_194),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_140),
.A2(n_166),
.B1(n_135),
.B2(n_138),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_119),
.B1(n_125),
.B2(n_117),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_189),
.B(n_215),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_100),
.B(n_108),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_144),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_136),
.A2(n_111),
.B1(n_117),
.B2(n_125),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_129),
.A2(n_100),
.B1(n_106),
.B2(n_113),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_203),
.B1(n_164),
.B2(n_143),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_129),
.A2(n_79),
.B1(n_113),
.B2(n_115),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_147),
.A2(n_108),
.B1(n_115),
.B2(n_97),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_121),
.C(n_97),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_201),
.C(n_177),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_142),
.A2(n_79),
.B1(n_155),
.B2(n_172),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_152),
.B1(n_128),
.B2(n_167),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_153),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_212),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_127),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_204),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_132),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_216),
.B(n_221),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_217),
.A2(n_239),
.B(n_248),
.Y(n_271)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_219),
.A2(n_232),
.B1(n_197),
.B2(n_248),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_148),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_185),
.B1(n_205),
.B2(n_184),
.Y(n_251)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_151),
.B(n_130),
.C(n_133),
.D(n_174),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_243),
.CI(n_178),
.CON(n_252),
.SN(n_252)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_182),
.B(n_151),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_236),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_184),
.B1(n_179),
.B2(n_187),
.Y(n_256)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_126),
.B1(n_157),
.B2(n_170),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_134),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_242),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_150),
.B(n_215),
.C(n_189),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_227),
.Y(n_272)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_188),
.A2(n_202),
.B(n_178),
.C(n_212),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_188),
.A2(n_202),
.B1(n_200),
.B2(n_194),
.Y(n_247)
);

AOI32xp33_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_183),
.A3(n_197),
.B1(n_243),
.B2(n_234),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_203),
.A2(n_176),
.B(n_180),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_198),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_251),
.A2(n_270),
.B1(n_247),
.B2(n_230),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_252),
.B(n_273),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_211),
.C(n_205),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_272),
.C(n_277),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_256),
.A2(n_259),
.B1(n_229),
.B2(n_218),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_179),
.B1(n_197),
.B2(n_183),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_269),
.A2(n_246),
.B1(n_249),
.B2(n_217),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_225),
.C(n_234),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_219),
.A2(n_232),
.B1(n_228),
.B2(n_222),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_253),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_302),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_225),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_295),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_271),
.B(n_273),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_282),
.A2(n_258),
.B(n_275),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_283),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_284),
.A2(n_254),
.B1(n_252),
.B2(n_260),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_288),
.B1(n_291),
.B2(n_299),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_240),
.B1(n_235),
.B2(n_224),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_231),
.B1(n_237),
.B2(n_250),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_223),
.B(n_245),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g321 ( 
.A1(n_292),
.A2(n_297),
.B(n_264),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_263),
.B(n_233),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_293),
.B(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_218),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_279),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_220),
.B(n_244),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_229),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_226),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_301),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_226),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_262),
.B1(n_267),
.B2(n_266),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_299),
.B1(n_287),
.B2(n_285),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_312),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_287),
.B1(n_298),
.B2(n_292),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_315),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_255),
.C(n_265),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_290),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_295),
.B(n_275),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_276),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_322),
.B(n_301),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_319),
.Y(n_325)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_289),
.A2(n_264),
.B(n_257),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_326),
.B(n_331),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_329),
.C(n_334),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_296),
.B1(n_292),
.B2(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_281),
.B1(n_258),
.B2(n_276),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_319),
.B1(n_304),
.B2(n_308),
.Y(n_332)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_317),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_316),
.C(n_307),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_321),
.B1(n_322),
.B2(n_304),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_336),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_310),
.Y(n_337)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

A2O1A1Ixp33_ASAP7_75t_SL g340 ( 
.A1(n_327),
.A2(n_322),
.B(n_321),
.C(n_318),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_349),
.Y(n_356)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_333),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_350),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_320),
.B(n_313),
.C(n_312),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_333),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_345),
.A2(n_332),
.B1(n_338),
.B2(n_323),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_352),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_339),
.A2(n_324),
.B1(n_331),
.B2(n_336),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_357),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_325),
.B1(n_324),
.B2(n_334),
.Y(n_354)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_354),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_305),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_355),
.A2(n_343),
.B(n_342),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_342),
.C(n_341),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_356),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_363),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_359),
.A2(n_355),
.B1(n_343),
.B2(n_356),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_346),
.C(n_358),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_SL g367 ( 
.A1(n_365),
.A2(n_328),
.B(n_349),
.C(n_340),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_366),
.B(n_340),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_368),
.A2(n_354),
.B1(n_340),
.B2(n_351),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_335),
.B(n_305),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_313),
.Y(n_371)
);


endmodule