module real_jpeg_2852_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_0),
.B(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_5),
.Y(n_43)
);

OR2x4_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

AO21x1_ASAP7_75t_L g11 ( 
.A1(n_2),
.A2(n_12),
.B(n_14),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_5),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_21),
.Y(n_34)
);

NAND2x1_ASAP7_75t_SL g35 ( 
.A(n_5),
.B(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_26),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_SL g7 ( 
.A1(n_8),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_16),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_25),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_23),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_38),
.B2(n_41),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OA21x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B(n_35),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);


endmodule