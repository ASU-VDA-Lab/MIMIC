module fake_jpeg_11327_n_399 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_399);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_399;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_57),
.Y(n_88)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_17),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_64),
.B(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_15),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_15),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_14),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_69),
.Y(n_94)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_30),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_29),
.B1(n_37),
.B2(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_71),
.A2(n_79),
.B1(n_82),
.B2(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_73),
.B(n_103),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_34),
.B1(n_23),
.B2(n_29),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_93),
.B1(n_98),
.B2(n_105),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_25),
.B1(n_32),
.B2(n_20),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_25),
.B1(n_32),
.B2(n_20),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_23),
.B1(n_20),
.B2(n_28),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_40),
.B1(n_55),
.B2(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_99),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_34),
.B1(n_30),
.B2(n_33),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_33),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_52),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_33),
.B1(n_36),
.B2(n_31),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_33),
.B1(n_32),
.B2(n_36),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_36),
.B1(n_31),
.B2(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_60),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_110),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_69),
.B1(n_51),
.B2(n_59),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_132),
.B1(n_48),
.B2(n_42),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_89),
.B1(n_80),
.B2(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_72),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_130),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_126),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_69),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_131),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_26),
.B1(n_56),
.B2(n_54),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_26),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_62),
.B1(n_42),
.B2(n_44),
.Y(n_132)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_138),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_52),
.B1(n_100),
.B2(n_95),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_0),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_73),
.B(n_74),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_94),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_157),
.B1(n_116),
.B2(n_125),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_103),
.B(n_84),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_146),
.A2(n_153),
.B(n_174),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_151),
.B1(n_155),
.B2(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_94),
.B1(n_74),
.B2(n_107),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_144),
.B1(n_128),
.B2(n_115),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_84),
.C(n_94),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_14),
.C(n_13),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_111),
.B1(n_132),
.B2(n_114),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_141),
.B(n_130),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_107),
.B1(n_104),
.B2(n_81),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_84),
.C(n_104),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_134),
.C(n_52),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_108),
.A2(n_75),
.B(n_81),
.C(n_90),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_131),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_112),
.A2(n_107),
.B1(n_80),
.B2(n_44),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_142),
.B1(n_123),
.B2(n_110),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_180),
.Y(n_228)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_146),
.B(n_161),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_171),
.B(n_159),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_186),
.B(n_188),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_193),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_138),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_208),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_159),
.B1(n_167),
.B2(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_110),
.B1(n_109),
.B2(n_113),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_135),
.B(n_134),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_200),
.B(n_211),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_140),
.B1(n_127),
.B2(n_76),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_140),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_205),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_153),
.A2(n_127),
.B1(n_100),
.B2(n_95),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_204),
.A2(n_206),
.B1(n_0),
.B2(n_1),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_97),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_100),
.B1(n_97),
.B2(n_62),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_166),
.C(n_168),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_13),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_158),
.B(n_14),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_164),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_45),
.B(n_137),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_219),
.Y(n_267)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_147),
.A3(n_158),
.B1(n_171),
.B2(n_168),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_234),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_147),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_175),
.B1(n_145),
.B2(n_152),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_220),
.B(n_233),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_230),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_165),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_225),
.B(n_229),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_238),
.B1(n_206),
.B2(n_201),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_180),
.A2(n_167),
.A3(n_176),
.B1(n_172),
.B2(n_162),
.C1(n_173),
.C2(n_165),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_172),
.C(n_162),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_169),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_184),
.A2(n_139),
.B1(n_137),
.B2(n_22),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_191),
.B(n_2),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_139),
.B1(n_22),
.B2(n_2),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_22),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_241),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_1),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_1),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_255),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_227),
.A2(n_184),
.B1(n_200),
.B2(n_211),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_260),
.B1(n_262),
.B2(n_265),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_187),
.B1(n_182),
.B2(n_202),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_248),
.A2(n_252),
.B1(n_259),
.B2(n_215),
.Y(n_286)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_182),
.B(n_188),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_198),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_196),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_261),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_204),
.B1(n_195),
.B2(n_192),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_227),
.A2(n_186),
.B1(n_181),
.B2(n_189),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_191),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_266),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_264)
);

XNOR2x2_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_6),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_223),
.A2(n_5),
.B(n_6),
.Y(n_266)
);

NAND2x1p5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_6),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_271),
.Y(n_294)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_215),
.A2(n_12),
.B1(n_7),
.B2(n_8),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_238),
.B1(n_241),
.B2(n_216),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_228),
.B1(n_214),
.B2(n_220),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_282),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_219),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_287),
.Y(n_303)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_217),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_268),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_239),
.C(n_234),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_293),
.C(n_296),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_292),
.B1(n_299),
.B2(n_273),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_233),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_257),
.A2(n_272),
.B1(n_254),
.B2(n_244),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_298),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_216),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_295),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_220),
.B1(n_240),
.B2(n_222),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_222),
.C(n_236),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_231),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_231),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_231),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_297),
.B(n_253),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_257),
.A2(n_231),
.B1(n_7),
.B2(n_8),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_252),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_300),
.A2(n_253),
.B(n_264),
.Y(n_322)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_305),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_245),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_317),
.Y(n_339)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_311),
.Y(n_326)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_260),
.C(n_258),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_284),
.C(n_291),
.Y(n_324)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_288),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_318),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_269),
.B(n_262),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_259),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_287),
.B(n_268),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_323),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_286),
.A2(n_292),
.B1(n_279),
.B2(n_293),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_289),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_290),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_266),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_314),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_332),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_327),
.B(n_338),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_323),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_295),
.C(n_296),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_334),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_278),
.C(n_274),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_298),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

XOR2x2_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_306),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_324),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_301),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_350),
.Y(n_358)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_351),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_307),
.B(n_308),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_246),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_314),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_356),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_246),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_354),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_331),
.B(n_312),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_340),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_359),
.A2(n_369),
.B(n_352),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_363),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_313),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_346),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_366),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_347),
.Y(n_366)
);

INVx11_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_367),
.A2(n_321),
.B1(n_335),
.B2(n_308),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_313),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_368),
.B(n_337),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_337),
.C(n_335),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_331),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_370),
.A2(n_371),
.B(n_372),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_364),
.A2(n_307),
.B(n_330),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_369),
.A2(n_361),
.B(n_357),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_320),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_343),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_365),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_376),
.A2(n_377),
.B(n_316),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_358),
.B(n_315),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_378),
.B(n_358),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_380),
.B(n_382),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_367),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_383),
.A2(n_385),
.B(n_387),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_365),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_386),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_375),
.A2(n_318),
.B(n_271),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_305),
.C(n_270),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_390),
.Y(n_394)
);

OAI221xp5_ASAP7_75t_SL g390 ( 
.A1(n_385),
.A2(n_264),
.B1(n_269),
.B2(n_255),
.C(n_250),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_299),
.Y(n_393)
);

OAI321xp33_ASAP7_75t_L g396 ( 
.A1(n_393),
.A2(n_395),
.A3(n_391),
.B1(n_300),
.B2(n_265),
.C(n_12),
.Y(n_396)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_396),
.A2(n_394),
.B(n_9),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_397),
.B(n_8),
.C(n_9),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_398),
.A2(n_12),
.B(n_392),
.Y(n_399)
);


endmodule