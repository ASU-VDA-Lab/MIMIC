module fake_jpeg_25574_n_99 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_11),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_32),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_57),
.B(n_58),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_39),
.B(n_35),
.C(n_41),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_39),
.B(n_33),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_41),
.B1(n_37),
.B2(n_38),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_63),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_59),
.B1(n_53),
.B2(n_50),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_71),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_74),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_6),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_77),
.C(n_80),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_20),
.B1(n_28),
.B2(n_27),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_19),
.B1(n_26),
.B2(n_25),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_79),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_79),
.Y(n_90)
);

AO221x1_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_81),
.B1(n_83),
.B2(n_72),
.C(n_73),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_68),
.B(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_92),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_86),
.C(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_82),
.B1(n_64),
.B2(n_72),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_18),
.C(n_13),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_16),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_17),
.Y(n_99)
);


endmodule