module fake_jpeg_8751_n_326 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_6),
.B(n_15),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_24),
.B1(n_21),
.B2(n_29),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_56),
.B1(n_69),
.B2(n_27),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_24),
.B1(n_29),
.B2(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_24),
.B1(n_21),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_71),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_24),
.B1(n_17),
.B2(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_75),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_46),
.B(n_37),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_41),
.B(n_48),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_81),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_53),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_17),
.C(n_34),
.Y(n_136)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_91),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_48),
.B1(n_28),
.B2(n_19),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_26),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_22),
.B1(n_17),
.B2(n_34),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_41),
.B(n_20),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g129 ( 
.A(n_93),
.B(n_105),
.C(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_102),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_97),
.Y(n_134)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_39),
.B1(n_42),
.B2(n_41),
.Y(n_101)
);

OAI22x1_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_68),
.B1(n_42),
.B2(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_18),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_22),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_18),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_121),
.B1(n_102),
.B2(n_84),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_59),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_113),
.A2(n_76),
.B(n_95),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_68),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_101),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_117),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_73),
.B1(n_87),
.B2(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_98),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_129),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_83),
.C(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_137),
.B1(n_95),
.B2(n_99),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_98),
.B(n_105),
.C(n_93),
.D(n_106),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_141),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_98),
.B1(n_105),
.B2(n_80),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_144),
.A2(n_149),
.B1(n_158),
.B2(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_160),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_48),
.B1(n_101),
.B2(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_151),
.A2(n_165),
.B(n_166),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_106),
.B1(n_79),
.B2(n_83),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_109),
.B1(n_135),
.B2(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_77),
.Y(n_155)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_116),
.C(n_114),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_126),
.C(n_114),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_101),
.B1(n_99),
.B2(n_89),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_112),
.B(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_170),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_78),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_112),
.B(n_76),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_184),
.C(n_185),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_SL g221 ( 
.A(n_173),
.B(n_178),
.C(n_189),
.Y(n_221)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_177),
.B(n_180),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_122),
.B1(n_110),
.B2(n_113),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_144),
.B(n_136),
.CI(n_113),
.CON(n_180),
.SN(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_113),
.B(n_122),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_190),
.B(n_191),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_163),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_135),
.Y(n_185)
);

AOI221xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_119),
.B1(n_136),
.B2(n_115),
.C(n_97),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_133),
.B(n_33),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_97),
.B(n_33),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_97),
.B(n_33),
.C(n_137),
.D(n_81),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_23),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_162),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_158),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_148),
.A2(n_133),
.B(n_23),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_164),
.B(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_159),
.B1(n_149),
.B2(n_157),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_223),
.B1(n_28),
.B2(n_1),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_218),
.B(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_140),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_211),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_159),
.C(n_154),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_220),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_177),
.B1(n_199),
.B2(n_145),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_178),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_173),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_229),
.Y(n_235)
);

NAND2x1p5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_142),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_174),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_28),
.C(n_19),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_230),
.C(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_175),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_172),
.B(n_8),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_9),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_28),
.C(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_179),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_253),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_239),
.C(n_242),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_219),
.B1(n_229),
.B2(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_185),
.C(n_181),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_191),
.B(n_175),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_204),
.B(n_211),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_180),
.C(n_197),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_194),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_180),
.C(n_203),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_246),
.C(n_248),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_221),
.C(n_206),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_186),
.C(n_176),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_215),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_206),
.C(n_205),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_207),
.C(n_208),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_7),
.C(n_15),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_216),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_209),
.B(n_7),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_262),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_252),
.B1(n_253),
.B2(n_250),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_260),
.A2(n_266),
.B1(n_264),
.B2(n_254),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_244),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_269),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_235),
.B(n_208),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_270),
.C(n_236),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_207),
.B(n_226),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_7),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_6),
.B(n_14),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_251),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_9),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_5),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_280),
.C(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_239),
.C(n_242),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_262),
.B(n_247),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_287),
.B(n_3),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_284),
.B1(n_280),
.B2(n_273),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_266),
.B1(n_254),
.B2(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_4),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_0),
.C(n_1),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_261),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_290),
.C(n_293),
.Y(n_310)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_259),
.B1(n_5),
.B2(n_11),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_284),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_295),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_259),
.Y(n_295)
);

FAx1_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_4),
.CI(n_12),
.CON(n_296),
.SN(n_296)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_286),
.B(n_14),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_4),
.Y(n_297)
);

AOI31xp67_ASAP7_75t_SL g308 ( 
.A1(n_297),
.A2(n_13),
.A3(n_16),
.B(n_296),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_16),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_13),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

INVx11_ASAP7_75t_L g305 ( 
.A(n_300),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_276),
.Y(n_301)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_13),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_296),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_307),
.B(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_289),
.C(n_288),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_300),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_312),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_315),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_303),
.C(n_305),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_305),
.B(n_309),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_312),
.C(n_314),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_321),
.B(n_317),
.C(n_311),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_320),
.B(n_322),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_302),
.Y(n_326)
);


endmodule