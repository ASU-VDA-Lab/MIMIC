module fake_aes_11244_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx3_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_10), .B(n_2), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_8), .B(n_4), .Y(n_14) );
BUFx3_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_6), .B(n_7), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_13), .A2(n_0), .B(n_1), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
AOI22xp33_ASAP7_75t_SL g19 ( .A1(n_16), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
AOI22xp33_ASAP7_75t_SL g21 ( .A1(n_18), .A2(n_16), .B1(n_15), .B2(n_12), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_18), .A2(n_11), .B(n_14), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_12), .B(n_11), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
NOR2x1_ASAP7_75t_L g27 ( .A(n_25), .B(n_16), .Y(n_27) );
OAI21xp5_ASAP7_75t_SL g28 ( .A1(n_27), .A2(n_19), .B(n_21), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_25), .Y(n_29) );
XOR2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_3), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
OAI211xp5_ASAP7_75t_SL g32 ( .A1(n_28), .A2(n_17), .B(n_14), .C(n_13), .Y(n_32) );
AND4x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_17), .C(n_23), .D(n_7), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_16), .B1(n_12), .B2(n_13), .Y(n_34) );
NAND2x1p5_ASAP7_75t_L g35 ( .A(n_32), .B(n_16), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
AND2x4_ASAP7_75t_L g37 ( .A(n_34), .B(n_12), .Y(n_37) );
OAI22xp5_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_33), .B1(n_11), .B2(n_12), .Y(n_38) );
AOI322xp5_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_4), .A3(n_5), .B1(n_11), .B2(n_37), .C1(n_31), .C2(n_36), .Y(n_39) );
endmodule