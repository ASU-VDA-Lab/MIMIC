module real_jpeg_12863_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_53),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_5),
.A2(n_19),
.B1(n_20),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_5),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_7),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_7),
.A2(n_22),
.B1(n_44),
.B2(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_7),
.B(n_76),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_24),
.C(n_26),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_7),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_7),
.B(n_23),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_85),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_83),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_69),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_69),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_68),
.Y(n_13)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_14)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_30),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_23),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_17),
.B(n_31),
.Y(n_109)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_19),
.A2(n_20),
.B1(n_24),
.B2(n_29),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_19),
.A2(n_22),
.B(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_19),
.A2(n_20),
.B1(n_41),
.B2(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_20),
.B(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_23),
.B(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_23),
.B(n_73),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_23)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_26),
.B(n_114),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_30),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_31),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_36),
.A2(n_40),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B(n_39),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_37),
.B(n_95),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_37),
.B(n_52),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_38),
.B(n_95),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_45),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_49),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_55),
.CI(n_59),
.CON(n_49),
.SN(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_51),
.B(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_54),
.B(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.C(n_80),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_74),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_129),
.B(n_133),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_110),
.B(n_128),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_104),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_104),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_96),
.B1(n_97),
.B2(n_103),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_101),
.C(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_121),
.B(n_127),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_117),
.B(n_120),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_131),
.Y(n_133)
);


endmodule