module fake_netlist_1_10056_n_44 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_44);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_44;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g15 ( .A(n_2), .B(n_8), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_9), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_8), .B(n_7), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_10), .B(n_6), .Y(n_21) );
AO22x1_ASAP7_75t_L g22 ( .A1(n_3), .A2(n_13), .B1(n_14), .B2(n_11), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_16), .B(n_0), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_16), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_19), .B(n_1), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_24), .B(n_21), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
AOI22xp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_27), .B1(n_28), .B2(n_25), .Y(n_32) );
OAI32xp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_27), .A3(n_26), .B1(n_15), .B2(n_30), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_28), .B(n_22), .Y(n_34) );
OAI21xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_32), .B(n_15), .Y(n_35) );
AOI22xp33_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_18), .B1(n_17), .B2(n_9), .Y(n_36) );
OAI322xp33_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_17), .A3(n_18), .B1(n_10), .B2(n_11), .C1(n_4), .C2(n_5), .Y(n_37) );
XNOR2xp5_ASAP7_75t_L g38 ( .A(n_35), .B(n_4), .Y(n_38) );
AND3x2_ASAP7_75t_L g39 ( .A(n_37), .B(n_5), .C(n_17), .Y(n_39) );
NAND2x1p5_ASAP7_75t_L g40 ( .A(n_37), .B(n_17), .Y(n_40) );
CKINVDCx20_ASAP7_75t_R g41 ( .A(n_38), .Y(n_41) );
AND2x2_ASAP7_75t_L g42 ( .A(n_40), .B(n_36), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_42), .Y(n_43) );
AOI322xp5_ASAP7_75t_L g44 ( .A1(n_43), .A2(n_41), .A3(n_42), .B1(n_18), .B2(n_39), .C1(n_40), .C2(n_12), .Y(n_44) );
endmodule