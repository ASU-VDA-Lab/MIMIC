module fake_jpeg_28897_n_539 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_539);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_77),
.Y(n_115)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_67),
.B(n_107),
.Y(n_160)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_94),
.Y(n_132)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g152 ( 
.A(n_85),
.Y(n_152)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_27),
.B(n_29),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_102),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_105),
.Y(n_138)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_22),
.Y(n_165)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_108),
.B1(n_50),
.B2(n_40),
.Y(n_124)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_116),
.A2(n_133),
.B1(n_137),
.B2(n_144),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_124),
.A2(n_145),
.B1(n_127),
.B2(n_137),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_23),
.B1(n_50),
.B2(n_40),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_127),
.A2(n_53),
.B1(n_48),
.B2(n_33),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_74),
.A2(n_40),
.B1(n_50),
.B2(n_23),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_72),
.A2(n_40),
.B1(n_50),
.B2(n_23),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_41),
.B(n_49),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_22),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_81),
.A2(n_102),
.B1(n_23),
.B2(n_40),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_61),
.A2(n_18),
.B1(n_44),
.B2(n_41),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_94),
.B(n_47),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_156),
.B(n_168),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_45),
.B1(n_26),
.B2(n_28),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_162),
.B1(n_163),
.B2(n_93),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_101),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_54),
.A2(n_73),
.B1(n_97),
.B2(n_96),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_57),
.B(n_44),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_56),
.B(n_35),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_33),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_34),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_22),
.Y(n_184)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_147),
.Y(n_173)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_173),
.Y(n_240)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_176),
.Y(n_250)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

AO22x1_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_22),
.B1(n_79),
.B2(n_69),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g263 ( 
.A1(n_178),
.A2(n_111),
.A3(n_148),
.B1(n_117),
.B2(n_120),
.Y(n_263)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_180),
.Y(n_228)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_123),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_187),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_214),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_129),
.A2(n_35),
.B1(n_23),
.B2(n_50),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_185),
.A2(n_215),
.B1(n_221),
.B2(n_139),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_66),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_161),
.Y(n_229)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_189),
.B(n_191),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_80),
.B1(n_58),
.B2(n_89),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_190),
.A2(n_220),
.B1(n_118),
.B2(n_125),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_192),
.B(n_213),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_115),
.B(n_48),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_193),
.B(n_195),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_95),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_199),
.Y(n_270)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_146),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_205),
.Y(n_260)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_145),
.A2(n_71),
.B1(n_87),
.B2(n_76),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_217),
.B1(n_224),
.B2(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_134),
.Y(n_205)
);

BUFx12_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_144),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_212),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

INVx11_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_157),
.A2(n_85),
.B1(n_56),
.B2(n_84),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_152),
.B(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_216),
.B(n_226),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_157),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_222),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_85),
.B1(n_53),
.B2(n_48),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_109),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_225),
.Y(n_230)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_109),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_231),
.A2(n_199),
.B1(n_172),
.B2(n_222),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_192),
.A2(n_124),
.B1(n_112),
.B2(n_118),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_237),
.A2(n_257),
.B1(n_53),
.B2(n_48),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_112),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_243),
.A2(n_201),
.B1(n_221),
.B2(n_208),
.Y(n_281)
);

HAxp5_ASAP7_75t_SL g245 ( 
.A(n_216),
.B(n_153),
.CON(n_245),
.SN(n_245)
);

OAI21xp33_ASAP7_75t_SL g288 ( 
.A1(n_245),
.A2(n_253),
.B(n_265),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_122),
.B(n_153),
.C(n_149),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_251),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_217),
.A2(n_200),
.B1(n_218),
.B2(n_125),
.Y(n_257)
);

AO22x1_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_207),
.B1(n_53),
.B2(n_48),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_154),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_268),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_194),
.B(n_122),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_227),
.B(n_149),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_174),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_110),
.Y(n_279)
);

AOI22x1_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_263),
.B1(n_217),
.B2(n_265),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_255),
.Y(n_311)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_177),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_277),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_175),
.A3(n_224),
.B1(n_194),
.B2(n_214),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_231),
.A2(n_120),
.B1(n_117),
.B2(n_154),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_278),
.A2(n_285),
.B1(n_290),
.B2(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_282),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_281),
.A2(n_296),
.B1(n_306),
.B2(n_247),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_198),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_188),
.B(n_173),
.C(n_210),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_283),
.A2(n_230),
.B(n_233),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_252),
.B(n_213),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_284),
.B(n_287),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_257),
.A2(n_242),
.B1(n_235),
.B2(n_237),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_228),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_233),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_1),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_235),
.A2(n_197),
.B1(n_203),
.B2(n_225),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_235),
.A2(n_212),
.B1(n_196),
.B2(n_211),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_292),
.A2(n_293),
.B1(n_307),
.B2(n_270),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_53),
.B1(n_48),
.B2(n_207),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_277),
.B(n_289),
.Y(n_337)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_53),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_299),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_260),
.B(n_2),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_3),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_234),
.B(n_4),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_228),
.B(n_33),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_247),
.B1(n_267),
.B2(n_270),
.Y(n_320)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_305),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_248),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_262),
.A2(n_33),
.B1(n_7),
.B2(n_8),
.Y(n_307)
);

XOR2x2_ASAP7_75t_SL g309 ( 
.A(n_272),
.B(n_262),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_247),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_275),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_310),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_311),
.A2(n_290),
.B1(n_293),
.B2(n_307),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_329),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_260),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_266),
.C(n_246),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_316),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_296),
.A2(n_251),
.B1(n_230),
.B2(n_249),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_327),
.B1(n_334),
.B2(n_287),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_324),
.A2(n_335),
.B1(n_294),
.B2(n_306),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_274),
.A2(n_251),
.B(n_244),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_325),
.A2(n_326),
.B(n_339),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_274),
.A2(n_244),
.B(n_230),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_256),
.C(n_238),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_266),
.C(n_246),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_238),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_288),
.A2(n_239),
.B(n_259),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_331),
.A2(n_283),
.B(n_303),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_295),
.A2(n_279),
.B1(n_304),
.B2(n_273),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_278),
.A2(n_249),
.B1(n_250),
.B2(n_261),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_267),
.B(n_33),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_295),
.A2(n_250),
.B1(n_239),
.B2(n_261),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_284),
.A2(n_273),
.B(n_300),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_341),
.A2(n_342),
.B1(n_346),
.B2(n_367),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_321),
.A2(n_286),
.B1(n_298),
.B2(n_292),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_313),
.B(n_276),
.Y(n_343)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_344),
.A2(n_351),
.B(n_358),
.Y(n_375)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_321),
.A2(n_333),
.B1(n_324),
.B2(n_339),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_330),
.Y(n_353)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_364),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_313),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_356),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_331),
.A2(n_301),
.B(n_299),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_311),
.A2(n_305),
.B(n_258),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_359),
.A2(n_363),
.B(n_316),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_361),
.B(n_368),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_368),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_311),
.A2(n_297),
.B1(n_241),
.B2(n_232),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_372),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_338),
.A2(n_280),
.B1(n_236),
.B2(n_232),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_333),
.A2(n_280),
.B1(n_232),
.B2(n_254),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_369),
.A2(n_371),
.B1(n_322),
.B2(n_327),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_309),
.A2(n_254),
.B1(n_247),
.B2(n_267),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_315),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_374),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_328),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_376),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_309),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_386),
.C(n_389),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_311),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_360),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_390),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_326),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_336),
.C(n_319),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_312),
.Y(n_391)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_391),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_394),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_319),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_400),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_345),
.C(n_371),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_397),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_360),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_343),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_404),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_399),
.A2(n_372),
.B(n_366),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_342),
.A2(n_334),
.B1(n_337),
.B2(n_332),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_355),
.B(n_323),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_403),
.A2(n_357),
.B1(n_341),
.B2(n_369),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_332),
.Y(n_404)
);

BUFx12f_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_419),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_SL g410 ( 
.A1(n_378),
.A2(n_372),
.B(n_337),
.C(n_344),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_410),
.A2(n_423),
.B(n_350),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_411),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_382),
.B(n_323),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_413),
.A2(n_432),
.B1(n_379),
.B2(n_373),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_390),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_375),
.A2(n_377),
.B(n_399),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_415),
.A2(n_381),
.B(n_402),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_348),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_422),
.Y(n_435)
);

NOR3xp33_ASAP7_75t_SL g419 ( 
.A(n_377),
.B(n_358),
.C(n_312),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_375),
.A2(n_367),
.B1(n_354),
.B2(n_337),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_420),
.A2(n_425),
.B1(n_414),
.B2(n_415),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_376),
.B(n_308),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_386),
.A2(n_359),
.B(n_363),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_395),
.A2(n_351),
.B1(n_372),
.B2(n_365),
.Y(n_425)
);

INVx13_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_408),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_308),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_428),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_310),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_423),
.B(n_410),
.Y(n_452)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_393),
.Y(n_430)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_430),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_353),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_4),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_389),
.B(n_352),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_388),
.B1(n_394),
.B2(n_374),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_434),
.A2(n_438),
.B1(n_447),
.B2(n_452),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_430),
.Y(n_436)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_392),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_437),
.B(n_441),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_407),
.A2(n_388),
.B1(n_400),
.B2(n_396),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_443),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_410),
.B1(n_407),
.B2(n_429),
.Y(n_464)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_418),
.Y(n_445)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_425),
.A2(n_403),
.B1(n_335),
.B2(n_381),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_449),
.A2(n_405),
.B1(n_412),
.B2(n_421),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_410),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_452),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_317),
.C(n_318),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_454),
.C(n_455),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_317),
.C(n_318),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_318),
.C(n_267),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_422),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_405),
.C(n_417),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_467),
.C(n_442),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_462),
.Y(n_491)
);

XOR2x1_ASAP7_75t_SL g463 ( 
.A(n_450),
.B(n_419),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_463),
.B(n_465),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_464),
.A2(n_435),
.B1(n_426),
.B2(n_408),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_417),
.C(n_432),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_468),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_446),
.B(n_409),
.Y(n_469)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_410),
.B1(n_426),
.B2(n_424),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_473),
.A2(n_474),
.B1(n_444),
.B2(n_445),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_455),
.A2(n_409),
.B(n_428),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_475),
.A2(n_442),
.B(n_440),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_481),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_438),
.C(n_434),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_484),
.C(n_486),
.Y(n_500)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_479),
.Y(n_493)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_480),
.Y(n_494)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_470),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_482),
.A2(n_483),
.B1(n_457),
.B2(n_463),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_471),
.A2(n_449),
.B1(n_441),
.B2(n_413),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_437),
.C(n_435),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_467),
.C(n_472),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_468),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_457),
.B(n_461),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_424),
.C(n_427),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_439),
.C(n_456),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_464),
.A2(n_408),
.B1(n_439),
.B2(n_431),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_487),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_478),
.B(n_459),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_496),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_465),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_498),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_499),
.A2(n_492),
.B1(n_489),
.B2(n_485),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_501),
.B(n_506),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_473),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_502),
.B(n_9),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_491),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_7),
.C(n_8),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_9),
.C(n_11),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_7),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_8),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_507),
.B(n_9),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_503),
.A2(n_476),
.B(n_489),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_508),
.A2(n_509),
.B(n_497),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_494),
.B(n_501),
.Y(n_509)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_510),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_515),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_485),
.C(n_483),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_518),
.C(n_493),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_517),
.Y(n_525)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_520),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_505),
.B(n_496),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_516),
.B(n_12),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_523),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_506),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_519),
.A2(n_510),
.B(n_512),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_526),
.A2(n_527),
.B(n_525),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_529),
.B(n_524),
.Y(n_530)
);

A2O1A1O1Ixp25_ASAP7_75t_L g534 ( 
.A1(n_530),
.A2(n_531),
.B(n_13),
.C(n_14),
.D(n_16),
.Y(n_534)
);

OAI21xp33_ASAP7_75t_SL g532 ( 
.A1(n_528),
.A2(n_11),
.B(n_12),
.Y(n_532)
);

MAJx2_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_11),
.C(n_12),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_533),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_535),
.A2(n_534),
.B(n_14),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_536),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_13),
.C(n_14),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_14),
.B(n_16),
.Y(n_539)
);


endmodule