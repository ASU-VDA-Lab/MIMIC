module real_aes_7247_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_1175;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1170;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_673;
wire n_635;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_1192;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1123;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_571;
wire n_1034;
wire n_952;
wire n_429;
wire n_976;
wire n_1166;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1110;
wire n_593;
wire n_1137;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_884;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_883;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1078;
wire n_1072;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_1053;
wire n_466;
wire n_1182;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1189;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_1168;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_996;
wire n_860;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_1174;
wire n_1100;
wire n_1167;
wire n_1193;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_1006;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_563;
wire n_997;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1157;
wire n_902;
wire n_1105;
wire n_1158;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1187;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_749;
wire n_1056;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_968;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_922;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_1191;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_1172;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_686;
wire n_776;
wire n_1190;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1045;
wire n_465;
wire n_967;
wire n_473;
wire n_566;
wire n_837;
wire n_719;
wire n_871;
wire n_1159;
wire n_474;
wire n_1156;
wire n_829;
wire n_1030;
wire n_1088;
wire n_1055;
wire n_988;
wire n_921;
wire n_597;
wire n_1176;
wire n_640;
wire n_483;
wire n_611;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_652;
wire n_1040;
wire n_703;
wire n_500;
wire n_601;
wire n_1185;
wire n_1076;
wire n_463;
wire n_661;
wire n_804;
wire n_1101;
wire n_447;
wire n_1102;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1119;
wire n_1039;
wire n_802;
wire n_868;
wire n_877;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_0), .A2(n_205), .B1(n_687), .B2(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g590 ( .A(n_1), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g1090 ( .A1(n_2), .A2(n_194), .B1(n_348), .B2(n_482), .C1(n_652), .C2(n_738), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_3), .A2(n_265), .B1(n_418), .B2(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_4), .A2(n_107), .B1(n_691), .B2(n_831), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g1149 ( .A1(n_5), .A2(n_341), .B1(n_644), .B2(n_691), .C(n_1150), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_6), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_7), .A2(n_178), .B1(n_861), .B2(n_891), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_8), .A2(n_84), .B1(n_715), .B2(n_738), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_9), .A2(n_249), .B1(n_467), .B2(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_SL g1019 ( .A(n_10), .B(n_1020), .Y(n_1019) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_11), .A2(n_237), .B1(n_424), .B2(n_429), .Y(n_432) );
INVx1_ASAP7_75t_L g1139 ( .A(n_11), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_12), .A2(n_187), .B1(n_643), .B2(n_744), .Y(n_1084) );
CKINVDCx20_ASAP7_75t_R g1120 ( .A(n_13), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_14), .A2(n_173), .B1(n_597), .B2(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_15), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_16), .Y(n_897) );
INVx1_ASAP7_75t_L g521 ( .A(n_17), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_18), .A2(n_210), .B1(n_706), .B2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_19), .A2(n_111), .B1(n_437), .B2(n_691), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_20), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_21), .A2(n_334), .B1(n_437), .B2(n_837), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_22), .A2(n_335), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g959 ( .A1(n_23), .A2(n_324), .B1(n_644), .B2(n_748), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_24), .A2(n_246), .B1(n_633), .B2(n_922), .Y(n_1007) );
AOI222xp33_ASAP7_75t_L g1075 ( .A1(n_25), .A2(n_68), .B1(n_293), .B2(n_570), .C1(n_852), .C2(n_1076), .Y(n_1075) );
AOI22xp33_ASAP7_75t_SL g839 ( .A1(n_26), .A2(n_323), .B1(n_720), .B2(n_840), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_27), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g1154 ( .A1(n_28), .A2(n_39), .B1(n_706), .B2(n_940), .C(n_1155), .Y(n_1154) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_29), .A2(n_319), .B1(n_748), .B2(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_30), .A2(n_380), .B1(n_551), .B2(n_861), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g1122 ( .A(n_31), .Y(n_1122) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_32), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_33), .A2(n_258), .B1(n_604), .B2(n_744), .Y(n_799) );
AO22x2_ASAP7_75t_L g434 ( .A1(n_34), .A2(n_126), .B1(n_424), .B2(n_425), .Y(n_434) );
INVx1_ASAP7_75t_L g987 ( .A(n_35), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_36), .A2(n_190), .B1(n_445), .B2(n_634), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g1077 ( .A(n_37), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_38), .A2(n_901), .B1(n_923), .B2(n_924), .Y(n_900) );
INVx1_ASAP7_75t_L g924 ( .A(n_38), .Y(n_924) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_40), .A2(n_63), .B1(n_643), .B2(n_749), .Y(n_802) );
INVx1_ASAP7_75t_L g563 ( .A(n_41), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_42), .A2(n_301), .B1(n_738), .B2(n_792), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_43), .A2(n_64), .B1(n_453), .B2(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g477 ( .A(n_44), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_45), .A2(n_182), .B1(n_743), .B2(n_744), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g1187 ( .A(n_46), .Y(n_1187) );
INVx1_ASAP7_75t_L g1152 ( .A(n_47), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_48), .A2(n_315), .B1(n_444), .B2(n_691), .Y(n_920) );
INVx1_ASAP7_75t_L g736 ( .A(n_49), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_50), .A2(n_225), .B1(n_496), .B2(n_529), .Y(n_561) );
AOI222xp33_ASAP7_75t_L g1158 ( .A1(n_51), .A2(n_147), .B1(n_160), .B2(n_482), .C1(n_657), .C2(n_819), .Y(n_1158) );
AOI222xp33_ASAP7_75t_L g942 ( .A1(n_52), .A2(n_310), .B1(n_333), .B2(n_677), .C1(n_770), .C2(n_906), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g1091 ( .A(n_53), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_54), .A2(n_127), .B1(n_1001), .B2(n_1045), .Y(n_1103) );
AOI22xp5_ASAP7_75t_SL g596 ( .A1(n_55), .A2(n_236), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g818 ( .A1(n_56), .A2(n_79), .B1(n_495), .B2(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g531 ( .A(n_57), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_58), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_59), .A2(n_193), .B1(n_633), .B2(n_1048), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_60), .A2(n_342), .B1(n_739), .B2(n_1071), .Y(n_1070) );
CKINVDCx16_ASAP7_75t_R g873 ( .A(n_61), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_62), .A2(n_313), .B1(n_827), .B2(n_911), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_65), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_66), .A2(n_378), .B1(n_544), .B2(n_545), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_67), .A2(n_285), .B1(n_495), .B2(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_69), .A2(n_96), .B1(n_738), .B2(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g992 ( .A(n_70), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g1142 ( .A1(n_71), .A2(n_1143), .B1(n_1144), .B2(n_1159), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g1159 ( .A(n_71), .Y(n_1159) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_72), .A2(n_138), .B1(n_553), .B2(n_723), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_73), .A2(n_366), .B1(n_643), .B2(n_916), .Y(n_1003) );
INVx1_ASAP7_75t_L g588 ( .A(n_74), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g1185 ( .A(n_75), .Y(n_1185) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_76), .B(n_576), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_77), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g1172 ( .A(n_78), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_80), .A2(n_97), .B1(n_540), .B2(n_776), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_81), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_82), .A2(n_273), .B1(n_826), .B2(n_827), .Y(n_1175) );
INVx1_ASAP7_75t_L g526 ( .A(n_83), .Y(n_526) );
AOI22xp5_ASAP7_75t_SL g602 ( .A1(n_85), .A2(n_100), .B1(n_603), .B2(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g499 ( .A(n_86), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_87), .A2(n_165), .B1(n_1051), .B2(n_1053), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_88), .A2(n_172), .B1(n_463), .B2(n_467), .Y(n_462) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_89), .A2(n_274), .B1(n_424), .B2(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g1136 ( .A(n_89), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_90), .A2(n_284), .B1(n_551), .B2(n_634), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_91), .A2(n_370), .B1(n_487), .B2(n_852), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_92), .A2(n_367), .B1(n_743), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_93), .A2(n_306), .B1(n_881), .B2(n_909), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_94), .A2(n_231), .B1(n_679), .B2(n_906), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_95), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_98), .A2(n_326), .B1(n_553), .B2(n_600), .Y(n_862) );
OA22x2_ASAP7_75t_L g928 ( .A1(n_99), .A2(n_929), .B1(n_930), .B2(n_943), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_99), .Y(n_929) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_101), .A2(n_218), .B1(n_444), .B2(n_576), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_102), .A2(n_120), .B1(n_604), .B2(n_723), .Y(n_745) );
INVx1_ASAP7_75t_L g472 ( .A(n_103), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_104), .A2(n_175), .B1(n_467), .B2(n_1111), .Y(n_1183) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_105), .A2(n_112), .B1(n_734), .B2(n_770), .Y(n_794) );
INVx1_ASAP7_75t_L g593 ( .A(n_106), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_108), .A2(n_250), .B1(n_463), .B2(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g435 ( .A(n_109), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_110), .A2(n_137), .B1(n_544), .B2(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g957 ( .A1(n_113), .A2(n_227), .B1(n_822), .B2(n_940), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_114), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_115), .B(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_116), .A2(n_154), .B1(n_837), .B2(n_1006), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_117), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_118), .A2(n_256), .B1(n_548), .B2(n_551), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g1036 ( .A(n_119), .Y(n_1036) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_121), .A2(n_292), .B1(n_598), .B2(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g455 ( .A(n_122), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_123), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_124), .Y(n_966) );
INVx1_ASAP7_75t_L g712 ( .A(n_125), .Y(n_712) );
INVx1_ASAP7_75t_L g1140 ( .A(n_126), .Y(n_1140) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_128), .A2(n_159), .B1(n_633), .B2(n_834), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_129), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_130), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g1107 ( .A(n_131), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_132), .A2(n_215), .B1(n_533), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_133), .A2(n_141), .B1(n_444), .B2(n_689), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_134), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_135), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_136), .A2(n_322), .B1(n_693), .B2(n_1182), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_139), .A2(n_217), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_140), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_142), .A2(n_275), .B1(n_827), .B2(n_911), .Y(n_1117) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_143), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g875 ( .A1(n_144), .A2(n_677), .B(n_876), .C(n_883), .Y(n_875) );
INVx1_ASAP7_75t_L g725 ( .A(n_145), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_146), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g1035 ( .A(n_148), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_149), .B(n_1174), .Y(n_1173) );
CKINVDCx20_ASAP7_75t_R g1102 ( .A(n_150), .Y(n_1102) );
INVx1_ASAP7_75t_L g751 ( .A(n_151), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_152), .A2(n_189), .B1(n_538), .B2(n_723), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_153), .A2(n_352), .B1(n_724), .B2(n_782), .Y(n_937) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_155), .A2(n_271), .B1(n_495), .B2(n_528), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g1000 ( .A1(n_156), .A2(n_254), .B1(n_840), .B2(n_1001), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g960 ( .A1(n_157), .A2(n_235), .B1(n_639), .B2(n_864), .Y(n_960) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_158), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_161), .A2(n_376), .B1(n_570), .B2(n_734), .Y(n_733) );
AOI211xp5_ASAP7_75t_L g961 ( .A1(n_162), .A2(n_544), .B(n_962), .C(n_967), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_163), .A2(n_414), .B1(n_511), .B2(n_512), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_163), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_164), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_166), .A2(n_201), .B1(n_634), .B2(n_749), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_167), .A2(n_375), .B1(n_826), .B2(n_827), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g1167 ( .A(n_168), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_169), .A2(n_287), .B1(n_529), .B2(n_826), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_170), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_171), .A2(n_247), .B1(n_467), .B2(n_922), .Y(n_921) );
AND2x6_ASAP7_75t_L g403 ( .A(n_174), .B(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_174), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_176), .A2(n_318), .B1(n_444), .B2(n_447), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_177), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_179), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_180), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_181), .A2(n_272), .B1(n_657), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g747 ( .A1(n_183), .A2(n_372), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_184), .A2(n_387), .B1(n_604), .B2(n_744), .Y(n_1026) );
AO22x1_ASAP7_75t_L g1147 ( .A1(n_185), .A2(n_197), .B1(n_1006), .B2(n_1148), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_186), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_188), .A2(n_351), .B1(n_418), .B2(n_778), .C(n_1147), .Y(n_1146) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_191), .A2(n_395), .B1(n_658), .B2(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g672 ( .A(n_192), .Y(n_672) );
INVx1_ASAP7_75t_L g492 ( .A(n_195), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_196), .Y(n_641) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_198), .A2(n_202), .B1(n_689), .B2(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g836 ( .A1(n_199), .A2(n_281), .B1(n_837), .B2(n_838), .Y(n_836) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_200), .A2(n_260), .B1(n_424), .B2(n_425), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g1137 ( .A(n_200), .B(n_1138), .Y(n_1137) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_203), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_204), .Y(n_1190) );
AOI211xp5_ASAP7_75t_L g1170 ( .A1(n_206), .A2(n_677), .B(n_1171), .C(n_1176), .Y(n_1170) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_207), .A2(n_280), .B1(n_778), .B2(n_859), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_208), .A2(n_262), .B1(n_538), .B2(n_600), .Y(n_1081) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_209), .A2(n_362), .B1(n_538), .B2(n_597), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g1178 ( .A(n_211), .Y(n_1178) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_212), .A2(n_350), .B1(n_538), .B2(n_540), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_213), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_214), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_216), .A2(n_251), .B1(n_744), .B2(n_864), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_219), .A2(n_358), .B1(n_634), .B2(n_782), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_220), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_221), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_222), .B(n_702), .Y(n_1088) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_223), .A2(n_369), .B1(n_739), .B2(n_826), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_224), .A2(n_625), .B1(n_664), .B2(n_665), .Y(n_624) );
INVx1_ASAP7_75t_L g664 ( .A(n_224), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g1115 ( .A(n_226), .Y(n_1115) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_228), .A2(n_261), .B1(n_826), .B2(n_827), .Y(n_825) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_229), .A2(n_399), .B(n_408), .C(n_1141), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_230), .A2(n_389), .B1(n_598), .B2(n_691), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_232), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_233), .Y(n_850) );
INVx1_ASAP7_75t_L g990 ( .A(n_234), .Y(n_990) );
CKINVDCx20_ASAP7_75t_R g1116 ( .A(n_238), .Y(n_1116) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_239), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_240), .A2(n_253), .B1(n_643), .B2(n_644), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_241), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_242), .A2(n_373), .B1(n_724), .B2(n_782), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_243), .B(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_244), .A2(n_308), .B1(n_827), .B2(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_245), .A2(n_384), .B1(n_720), .B2(n_864), .Y(n_1085) );
XNOR2xp5_ASAP7_75t_L g813 ( .A(n_248), .B(n_814), .Y(n_813) );
AOI22xp5_ASAP7_75t_SL g982 ( .A1(n_252), .A2(n_983), .B1(n_1008), .B2(n_1009), .Y(n_982) );
INVx1_ASAP7_75t_L g1009 ( .A(n_252), .Y(n_1009) );
INVx2_ASAP7_75t_L g407 ( .A(n_255), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g1016 ( .A1(n_257), .A2(n_340), .B1(n_496), .B2(n_570), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_259), .Y(n_950) );
INVx1_ASAP7_75t_L g986 ( .A(n_263), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_264), .A2(n_279), .B1(n_718), .B2(n_778), .Y(n_1067) );
OA22x2_ASAP7_75t_L g515 ( .A1(n_266), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_266), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_267), .A2(n_298), .B1(n_553), .B2(n_554), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_268), .A2(n_1095), .B1(n_1123), .B2(n_1124), .Y(n_1094) );
INVx1_ASAP7_75t_L g1123 ( .A(n_268), .Y(n_1123) );
INVx1_ASAP7_75t_L g996 ( .A(n_269), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_270), .A2(n_329), .B1(n_640), .B2(n_723), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_276), .A2(n_328), .B1(n_467), .B2(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_277), .A2(n_377), .B1(n_540), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g560 ( .A(n_278), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_282), .A2(n_397), .B1(n_834), .B2(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_283), .A2(n_365), .B1(n_686), .B2(n_687), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_286), .A2(n_332), .B1(n_909), .B2(n_940), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g1018 ( .A(n_288), .B(n_706), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_289), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_290), .A2(n_345), .B1(n_1001), .B2(n_1055), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_291), .A2(n_381), .B1(n_706), .B2(n_881), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_294), .Y(n_612) );
INVx1_ASAP7_75t_L g424 ( .A(n_295), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_295), .Y(n_426) );
INVx1_ASAP7_75t_L g763 ( .A(n_296), .Y(n_763) );
INVx1_ASAP7_75t_L g485 ( .A(n_297), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g1031 ( .A1(n_299), .A2(n_1032), .B1(n_1056), .B2(n_1057), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_299), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_300), .Y(n_964) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_302), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_303), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g1156 ( .A(n_304), .Y(n_1156) );
CKINVDCx20_ASAP7_75t_R g1189 ( .A(n_305), .Y(n_1189) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_307), .A2(n_354), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g762 ( .A(n_309), .Y(n_762) );
INVx1_ASAP7_75t_L g461 ( .A(n_311), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_312), .Y(n_620) );
INVx1_ASAP7_75t_L g673 ( .A(n_314), .Y(n_673) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_316), .A2(n_364), .B1(n_709), .B2(n_739), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g1119 ( .A(n_317), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_320), .B(n_657), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_321), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_325), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_327), .A2(n_355), .B1(n_528), .B2(n_734), .Y(n_1089) );
NAND2xp5_ASAP7_75t_SL g824 ( .A(n_330), .B(n_796), .Y(n_824) );
AO22x2_ASAP7_75t_L g842 ( .A1(n_331), .A2(n_843), .B1(n_865), .B2(n_866), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_331), .Y(n_866) );
INVx1_ASAP7_75t_L g406 ( .A(n_336), .Y(n_406) );
AOI22xp5_ASAP7_75t_SL g668 ( .A1(n_337), .A2(n_669), .B1(n_694), .B2(n_695), .Y(n_668) );
INVx1_ASAP7_75t_L g695 ( .A(n_337), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_338), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g404 ( .A(n_339), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_343), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_344), .B(n_702), .Y(n_732) );
INVx1_ASAP7_75t_L g504 ( .A(n_346), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_347), .B(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g591 ( .A(n_349), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_353), .B(n_881), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g1177 ( .A(n_356), .Y(n_1177) );
INVx1_ASAP7_75t_L g534 ( .A(n_357), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g1109 ( .A(n_359), .Y(n_1109) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_360), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_361), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g1087 ( .A(n_363), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_368), .Y(n_771) );
INVx1_ASAP7_75t_L g898 ( .A(n_371), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_374), .B(n_702), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_379), .Y(n_895) );
INVx1_ASAP7_75t_L g523 ( .A(n_382), .Y(n_523) );
INVx1_ASAP7_75t_L g995 ( .A(n_383), .Y(n_995) );
INVx1_ASAP7_75t_L g1151 ( .A(n_385), .Y(n_1151) );
XNOR2xp5_ASAP7_75t_L g945 ( .A(n_386), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g442 ( .A(n_388), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_390), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_391), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g1157 ( .A(n_392), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_393), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_394), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_396), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_404), .Y(n_1132) );
OAI21xp5_ASAP7_75t_L g1165 ( .A1(n_405), .A2(n_1131), .B(n_1166), .Y(n_1165) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_975), .B1(n_1126), .B2(n_1127), .C(n_1128), .Y(n_408) );
INVx1_ASAP7_75t_L g1126 ( .A(n_409), .Y(n_1126) );
XOR2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_808), .Y(n_409) );
XOR2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_622), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
XNOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_513), .Y(n_412) );
INVx1_ASAP7_75t_L g512 ( .A(n_414), .Y(n_512) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_415), .B(n_470), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_451), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_435), .B1(n_436), .B2(n_442), .C(n_443), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_417), .A2(n_456), .B1(n_897), .B2(n_898), .Y(n_896) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g636 ( .A(n_419), .Y(n_636) );
BUFx3_ASAP7_75t_L g837 ( .A(n_419), .Y(n_837) );
BUFx3_ASAP7_75t_L g1045 ( .A(n_419), .Y(n_1045) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_SL g544 ( .A(n_420), .Y(n_544) );
INVx2_ASAP7_75t_L g578 ( .A(n_420), .Y(n_578) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_430), .Y(n_420) );
AND2x6_ASAP7_75t_L g439 ( .A(n_421), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g453 ( .A(n_421), .B(n_454), .Y(n_453) );
AND2x6_ASAP7_75t_L g483 ( .A(n_421), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g446 ( .A(n_422), .B(n_428), .Y(n_446) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_423), .B(n_428), .Y(n_450) );
AND2x2_ASAP7_75t_L g459 ( .A(n_423), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g491 ( .A(n_423), .B(n_432), .Y(n_491) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_426), .Y(n_429) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
INVx1_ASAP7_75t_L g490 ( .A(n_428), .Y(n_490) );
AND2x4_ASAP7_75t_L g445 ( .A(n_430), .B(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g448 ( .A(n_430), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_430), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g542 ( .A(n_430), .B(n_459), .Y(n_542) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
OR2x2_ASAP7_75t_L g441 ( .A(n_431), .B(n_434), .Y(n_441) );
AND2x2_ASAP7_75t_L g454 ( .A(n_431), .B(n_434), .Y(n_454) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g484 ( .A(n_432), .B(n_434), .Y(n_484) );
AND2x2_ASAP7_75t_L g489 ( .A(n_433), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g503 ( .A(n_433), .Y(n_503) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g469 ( .A(n_434), .Y(n_469) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g603 ( .A(n_438), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g627 ( .A1(n_438), .A2(n_628), .B1(n_629), .B2(n_630), .C(n_631), .Y(n_627) );
INVx3_ASAP7_75t_L g778 ( .A(n_438), .Y(n_778) );
INVx11_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx11_ASAP7_75t_L g539 ( .A(n_439), .Y(n_539) );
AND2x4_ASAP7_75t_L g704 ( .A(n_440), .B(n_446), .Y(n_704) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g475 ( .A(n_441), .B(n_476), .Y(n_475) );
INVx4_ASAP7_75t_L g783 ( .A(n_444), .Y(n_783) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g553 ( .A(n_445), .Y(n_553) );
INVx2_ASAP7_75t_L g573 ( .A(n_445), .Y(n_573) );
BUFx3_ASAP7_75t_L g640 ( .A(n_445), .Y(n_640) );
BUFx3_ASAP7_75t_L g720 ( .A(n_445), .Y(n_720) );
INVx1_ASAP7_75t_L g476 ( .A(n_446), .Y(n_476) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_446), .B(n_454), .Y(n_479) );
AND2x6_ASAP7_75t_L g707 ( .A(n_446), .B(n_454), .Y(n_707) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx3_ASAP7_75t_L g545 ( .A(n_448), .Y(n_545) );
INVx1_ASAP7_75t_L g584 ( .A(n_448), .Y(n_584) );
BUFx3_ASAP7_75t_L g604 ( .A(n_448), .Y(n_604) );
BUFx2_ASAP7_75t_SL g687 ( .A(n_448), .Y(n_687) );
BUFx2_ASAP7_75t_L g724 ( .A(n_448), .Y(n_724) );
BUFx2_ASAP7_75t_SL g776 ( .A(n_448), .Y(n_776) );
BUFx3_ASAP7_75t_L g864 ( .A(n_448), .Y(n_864) );
AND2x2_ASAP7_75t_L g576 ( .A(n_449), .B(n_503), .Y(n_576) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x6_ASAP7_75t_L g468 ( .A(n_450), .B(n_469), .Y(n_468) );
OAI221xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_455), .B1(n_456), .B2(n_461), .C(n_462), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g577 ( .A1(n_452), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_577) );
INVx3_ASAP7_75t_L g643 ( .A(n_452), .Y(n_643) );
INVx2_ASAP7_75t_L g691 ( .A(n_452), .Y(n_691) );
INVx2_ASAP7_75t_L g718 ( .A(n_452), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_452), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_892) );
INVx2_ASAP7_75t_L g1053 ( .A(n_452), .Y(n_1053) );
INVx6_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g550 ( .A(n_453), .Y(n_550) );
BUFx3_ASAP7_75t_L g748 ( .A(n_453), .Y(n_748) );
BUFx3_ASAP7_75t_L g859 ( .A(n_453), .Y(n_859) );
AND2x2_ASAP7_75t_L g466 ( .A(n_454), .B(n_459), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_454), .B(n_459), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_456), .A2(n_1185), .B1(n_1186), .B2(n_1187), .Y(n_1184) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_458), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g510 ( .A(n_460), .Y(n_510) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g551 ( .A(n_465), .Y(n_551) );
INVx3_ASAP7_75t_L g598 ( .A(n_465), .Y(n_598) );
INVx5_ASAP7_75t_L g749 ( .A(n_465), .Y(n_749) );
INVx4_ASAP7_75t_L g835 ( .A(n_465), .Y(n_835) );
INVx1_ASAP7_75t_L g891 ( .A(n_465), .Y(n_891) );
INVx8_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g554 ( .A(n_468), .Y(n_554) );
INVx6_ASAP7_75t_SL g634 ( .A(n_468), .Y(n_634) );
INVx1_ASAP7_75t_SL g689 ( .A(n_468), .Y(n_689) );
INVx1_ASAP7_75t_L g710 ( .A(n_469), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .C(n_498), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_477), .B2(n_478), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_473), .A2(n_478), .B1(n_762), .B2(n_763), .Y(n_761) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g648 ( .A(n_474), .Y(n_648) );
INVx2_ASAP7_75t_L g847 ( .A(n_474), .Y(n_847) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_475), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_475), .A2(n_560), .B(n_561), .Y(n_559) );
BUFx3_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_478), .A2(n_502), .B1(n_563), .B2(n_564), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_478), .A2(n_648), .B1(n_672), .B2(n_673), .Y(n_671) );
INVx2_ASAP7_75t_L g879 ( .A(n_478), .Y(n_879) );
OA211x2_ASAP7_75t_L g1086 ( .A1(n_478), .A2(n_1087), .B(n_1088), .C(n_1089), .Y(n_1086) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g609 ( .A(n_479), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_485), .B1(n_486), .B2(n_492), .C(n_493), .Y(n_480) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_481), .A2(n_526), .B(n_527), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g764 ( .A1(n_481), .A2(n_765), .B(n_766), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g989 ( .A1(n_481), .A2(n_990), .B1(n_991), .B2(n_992), .C(n_993), .Y(n_989) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g654 ( .A(n_482), .Y(n_654) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_SL g567 ( .A(n_483), .Y(n_567) );
INVx4_ASAP7_75t_L g617 ( .A(n_483), .Y(n_617) );
BUFx3_ASAP7_75t_L g677 ( .A(n_483), .Y(n_677) );
INVx2_ASAP7_75t_L g713 ( .A(n_483), .Y(n_713) );
INVx2_ASAP7_75t_L g949 ( .A(n_483), .Y(n_949) );
INVx1_ASAP7_75t_L g508 ( .A(n_484), .Y(n_508) );
AND2x4_ASAP7_75t_L g529 ( .A(n_484), .B(n_510), .Y(n_529) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_488), .Y(n_533) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_488), .Y(n_570) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_488), .Y(n_652) );
BUFx4f_ASAP7_75t_SL g770 ( .A(n_488), .Y(n_770) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g497 ( .A(n_490), .Y(n_497) );
AND2x4_ASAP7_75t_L g496 ( .A(n_491), .B(n_497), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_491), .B(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g709 ( .A(n_491), .B(n_710), .Y(n_709) );
BUFx4f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g953 ( .A(n_495), .Y(n_953) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_496), .Y(n_658) );
BUFx12f_ASAP7_75t_L g738 ( .A(n_496), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_504), .B2(n_505), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_500), .A2(n_507), .B1(n_855), .B2(n_856), .Y(n_854) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx3_ASAP7_75t_SL g611 ( .A(n_501), .Y(n_611) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_502), .A2(n_531), .B1(n_532), .B2(n_534), .Y(n_530) );
BUFx3_ASAP7_75t_L g662 ( .A(n_502), .Y(n_662) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_502), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_502), .A2(n_505), .B1(n_1156), .B2(n_1157), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_505), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g683 ( .A(n_506), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g997 ( .A(n_507), .Y(n_997) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AO22x2_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_555), .B2(n_621), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_535), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .C(n_530), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g613 ( .A1(n_522), .A2(n_614), .B(n_615), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g985 ( .A1(n_522), .A2(n_986), .B1(n_987), .B2(n_988), .Y(n_985) );
OAI221xp5_ASAP7_75t_SL g1114 ( .A1(n_524), .A2(n_648), .B1(n_1115), .B2(n_1116), .C(n_1117), .Y(n_1114) );
OAI211xp5_ASAP7_75t_L g1171 ( .A1(n_524), .A2(n_1172), .B(n_1173), .C(n_1175), .Y(n_1171) );
INVx1_ASAP7_75t_SL g828 ( .A(n_528), .Y(n_828) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_SL g715 ( .A(n_529), .Y(n_715) );
BUFx3_ASAP7_75t_L g739 ( .A(n_529), .Y(n_739) );
BUFx2_ASAP7_75t_SL g792 ( .A(n_529), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_532), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_883) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_533), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_546), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .Y(n_536) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_538), .Y(n_1182) );
INVx5_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_539), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_SL g743 ( .A(n_539), .Y(n_743) );
INVx4_ASAP7_75t_L g838 ( .A(n_539), .Y(n_838) );
INVx2_ASAP7_75t_L g916 ( .A(n_539), .Y(n_916) );
INVx1_ASAP7_75t_L g1099 ( .A(n_539), .Y(n_1099) );
BUFx4f_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g1002 ( .A(n_541), .Y(n_1002) );
BUFx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g597 ( .A(n_542), .Y(n_597) );
BUFx3_ASAP7_75t_L g744 ( .A(n_542), .Y(n_744) );
BUFx3_ASAP7_75t_L g918 ( .A(n_542), .Y(n_918) );
INVx2_ASAP7_75t_L g629 ( .A(n_545), .Y(n_629) );
HB1xp67_ASAP7_75t_L g1148 ( .A(n_545), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_552), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_551), .Y(n_632) );
BUFx2_ASAP7_75t_L g1106 ( .A(n_553), .Y(n_1106) );
INVx2_ASAP7_75t_L g621 ( .A(n_555), .Y(n_621) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_592), .Y(n_555) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_591), .Y(n_556) );
AND3x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_571), .C(n_581), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .C(n_565), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_565) );
OAI222xp33_ASAP7_75t_L g1118 ( .A1(n_567), .A2(n_769), .B1(n_1119), .B2(n_1120), .C1(n_1121), .C2(n_1122), .Y(n_1118) );
INVx3_ASAP7_75t_L g819 ( .A(n_569), .Y(n_819) );
INVx4_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g619 ( .A(n_570), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_577), .Y(n_571) );
OAI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B(n_575), .Y(n_572) );
INVx2_ASAP7_75t_L g686 ( .A(n_573), .Y(n_686) );
INVx1_ASAP7_75t_L g1046 ( .A(n_573), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_573), .A2(n_1189), .B1(n_1190), .B2(n_1191), .Y(n_1188) );
INVx3_ASAP7_75t_L g600 ( .A(n_578), .Y(n_600) );
INVx3_ASAP7_75t_L g723 ( .A(n_578), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_587), .C(n_589), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_582) );
BUFx2_ASAP7_75t_R g963 ( .A(n_586), .Y(n_963) );
XNOR2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND3x1_ASAP7_75t_SL g594 ( .A(n_595), .B(n_601), .C(n_606), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
BUFx2_ASAP7_75t_L g644 ( .A(n_597), .Y(n_644) );
INVx1_ASAP7_75t_L g832 ( .A(n_597), .Y(n_832) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g969 ( .A(n_603), .Y(n_969) );
BUFx2_ASAP7_75t_L g1055 ( .A(n_604), .Y(n_1055) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_613), .C(n_616), .Y(n_606) );
OAI22xp5_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_610), .B1(n_611), .B2(n_612), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_608), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_608), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_845) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g988 ( .A(n_609), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_611), .A2(n_995), .B1(n_996), .B2(n_997), .Y(n_994) );
OAI22xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_616) );
INVx4_ASAP7_75t_L g1076 ( .A(n_617), .Y(n_1076) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_666), .B1(n_806), .B2(n_807), .Y(n_622) );
INVx3_ASAP7_75t_L g806 ( .A(n_623), .Y(n_806) );
BUFx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g665 ( .A(n_625), .Y(n_665) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_626), .B(n_645), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_635), .Y(n_626) );
INVx2_ASAP7_75t_L g840 ( .A(n_629), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g1153 ( .A(n_633), .Y(n_1153) );
BUFx4f_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g861 ( .A(n_634), .Y(n_861) );
BUFx2_ASAP7_75t_L g934 ( .A(n_634), .Y(n_934) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_637), .B1(n_638), .B2(n_641), .C(n_642), .Y(n_635) );
INVx2_ASAP7_75t_L g693 ( .A(n_636), .Y(n_693) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_650), .C(n_660), .Y(n_645) );
OAI222xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_654), .B2(n_655), .C1(n_656), .C2(n_659), .Y(n_650) );
OAI222xp33_ASAP7_75t_L g1038 ( .A1(n_651), .A2(n_656), .B1(n_713), .B2(n_1039), .C1(n_1040), .C2(n_1041), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g816 ( .A1(n_654), .A2(n_817), .B(n_818), .Y(n_816) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g1121 ( .A(n_658), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_662), .A2(n_681), .B1(n_682), .B2(n_683), .Y(n_680) );
INVx1_ASAP7_75t_L g807 ( .A(n_666), .Y(n_807) );
XOR2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_754), .Y(n_666) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_696), .B1(n_752), .B2(n_753), .Y(n_667) );
INVx1_ASAP7_75t_L g752 ( .A(n_668), .Y(n_752) );
INVx2_ASAP7_75t_SL g694 ( .A(n_669), .Y(n_694) );
AND2x2_ASAP7_75t_SL g669 ( .A(n_670), .B(n_684), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .C(n_680), .Y(n_670) );
OAI21xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B(n_678), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g849 ( .A1(n_676), .A2(n_850), .B(n_851), .Y(n_849) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g951 ( .A(n_679), .Y(n_951) );
AND4x1_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .C(n_690), .D(n_692), .Y(n_684) );
INVx1_ASAP7_75t_L g753 ( .A(n_696), .Y(n_753) );
XOR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_726), .Y(n_696) );
OA22x2_ASAP7_75t_L g754 ( .A1(n_697), .A2(n_755), .B1(n_756), .B2(n_805), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_697), .Y(n_755) );
XOR2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_725), .Y(n_697) );
NAND4xp75_ASAP7_75t_SL g698 ( .A(n_699), .B(n_716), .C(n_721), .D(n_722), .Y(n_698) );
NOR2xp67_ASAP7_75t_SL g699 ( .A(n_700), .B(n_711), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_705), .C(n_708), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx5_ASAP7_75t_L g796 ( .A(n_703), .Y(n_796) );
INVx2_ASAP7_75t_L g881 ( .A(n_703), .Y(n_881) );
INVx2_ASAP7_75t_L g1020 ( .A(n_703), .Y(n_1020) );
INVx4_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g823 ( .A(n_706), .Y(n_823) );
BUFx4f_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g731 ( .A(n_707), .Y(n_731) );
BUFx2_ASAP7_75t_L g909 ( .A(n_707), .Y(n_909) );
BUFx3_ASAP7_75t_L g734 ( .A(n_709), .Y(n_734) );
BUFx2_ASAP7_75t_L g826 ( .A(n_709), .Y(n_826) );
INVx1_ASAP7_75t_L g912 ( .A(n_709), .Y(n_912) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_709), .Y(n_1071) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B(n_714), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g735 ( .A1(n_713), .A2(n_736), .B(n_737), .Y(n_735) );
OAI21xp5_ASAP7_75t_L g789 ( .A1(n_713), .A2(n_790), .B(n_791), .Y(n_789) );
OAI21xp5_ASAP7_75t_SL g903 ( .A1(n_713), .A2(n_904), .B(n_905), .Y(n_903) );
OAI21xp5_ASAP7_75t_SL g1014 ( .A1(n_713), .A2(n_1015), .B(n_1016), .Y(n_1014) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_720), .Y(n_1006) );
XOR2x2_ASAP7_75t_SL g726 ( .A(n_727), .B(n_751), .Y(n_726) );
NAND2x1p5_ASAP7_75t_L g727 ( .A(n_728), .B(n_740), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_735), .Y(n_728) );
NAND3xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .C(n_733), .Y(n_729) );
INVx2_ASAP7_75t_L g853 ( .A(n_738), .Y(n_853) );
BUFx4f_ASAP7_75t_SL g906 ( .A(n_738), .Y(n_906) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_746), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g1052 ( .A(n_743), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_750), .Y(n_746) );
BUFx6f_ASAP7_75t_L g922 ( .A(n_749), .Y(n_922) );
BUFx2_ASAP7_75t_L g1048 ( .A(n_749), .Y(n_1048) );
INVx1_ASAP7_75t_L g805 ( .A(n_756), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_785), .B2(n_786), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
XNOR2x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_784), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_773), .Y(n_759) );
NOR3xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_764), .C(n_767), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B1(n_771), .B2(n_772), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_774), .B(n_779), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g1108 ( .A(n_776), .Y(n_1108) );
INVx1_ASAP7_75t_L g894 ( .A(n_778), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx3_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
XOR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_804), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g787 ( .A(n_788), .B(n_797), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_793), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
BUFx6f_ASAP7_75t_L g940 ( .A(n_796), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_867), .B1(n_868), .B2(n_974), .Y(n_808) );
INVx1_ASAP7_75t_L g974 ( .A(n_809), .Y(n_974) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AO22x1_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B1(n_841), .B2(n_842), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND4xp75_ASAP7_75t_SL g814 ( .A(n_815), .B(n_829), .C(n_836), .D(n_839), .Y(n_814) );
NOR2xp67_ASAP7_75t_L g815 ( .A(n_816), .B(n_820), .Y(n_815) );
INVx1_ASAP7_75t_L g991 ( .A(n_819), .Y(n_991) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .C(n_825), .Y(n_820) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AND2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g1112 ( .A(n_835), .Y(n_1112) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
XNOR2x2_ASAP7_75t_L g899 ( .A(n_842), .B(n_900), .Y(n_899) );
INVx1_ASAP7_75t_SL g865 ( .A(n_843), .Y(n_865) );
AND2x2_ASAP7_75t_SL g843 ( .A(n_844), .B(n_857), .Y(n_843) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_849), .C(n_854), .Y(n_844) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_847), .A2(n_878), .B1(n_1035), .B2(n_1036), .C(n_1037), .Y(n_1034) );
INVx1_ASAP7_75t_L g886 ( .A(n_852), .Y(n_886) );
INVx3_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
AND4x1_ASAP7_75t_L g857 ( .A(n_858), .B(n_860), .C(n_862), .D(n_863), .Y(n_857) );
INVx1_ASAP7_75t_L g1101 ( .A(n_859), .Y(n_1101) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OAI22xp5_ASAP7_75t_SL g868 ( .A1(n_869), .A2(n_926), .B1(n_927), .B2(n_973), .Y(n_868) );
INVx2_ASAP7_75t_SL g973 ( .A(n_869), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_871), .B1(n_899), .B2(n_925), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_871), .A2(n_872), .B1(n_945), .B2(n_970), .Y(n_944) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
XNOR2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_887), .Y(n_874) );
OAI211xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_878), .B(n_880), .C(n_882), .Y(n_876) );
INVx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_886), .A2(n_951), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
NOR3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_892), .C(n_896), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
INVx2_ASAP7_75t_L g925 ( .A(n_899), .Y(n_925) );
INVx2_ASAP7_75t_SL g923 ( .A(n_901), .Y(n_923) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_913), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_907), .Y(n_902) );
NAND2xp5_ASAP7_75t_SL g907 ( .A(n_908), .B(n_910), .Y(n_907) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_919), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_917), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_944), .B1(n_971), .B2(n_972), .Y(n_927) );
INVx1_ASAP7_75t_L g972 ( .A(n_928), .Y(n_972) );
INVx1_ASAP7_75t_SL g943 ( .A(n_930), .Y(n_943) );
NAND4xp75_ASAP7_75t_L g930 ( .A(n_931), .B(n_935), .C(n_938), .D(n_942), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_932), .B(n_933), .Y(n_931) );
INVx1_ASAP7_75t_L g965 ( .A(n_934), .Y(n_965) );
AND2x2_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
AND2x2_ASAP7_75t_SL g938 ( .A(n_939), .B(n_941), .Y(n_938) );
INVx1_ASAP7_75t_L g971 ( .A(n_944), .Y(n_971) );
INVx1_ASAP7_75t_L g970 ( .A(n_945), .Y(n_970) );
NAND3x1_ASAP7_75t_L g946 ( .A(n_947), .B(n_958), .C(n_961), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_955), .Y(n_947) );
OAI222xp33_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_950), .B1(n_951), .B2(n_952), .C1(n_953), .C2(n_954), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
OAI22xp5_ASAP7_75t_SL g962 ( .A1(n_963), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_963), .A2(n_1151), .B1(n_1152), .B2(n_1153), .Y(n_1150) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
INVx1_ASAP7_75t_L g1127 ( .A(n_975), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_977), .B1(n_1058), .B2(n_1059), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
BUFx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OAI22xp5_ASAP7_75t_SL g979 ( .A1(n_980), .A2(n_981), .B1(n_1030), .B2(n_1031), .Y(n_979) );
INVx2_ASAP7_75t_SL g980 ( .A(n_981), .Y(n_980) );
OA22x2_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_1010), .B1(n_1011), .B2(n_1029), .Y(n_981) );
INVx1_ASAP7_75t_L g1029 ( .A(n_982), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_983), .Y(n_1008) );
AND2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_998), .Y(n_983) );
NOR3xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_989), .C(n_994), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1004), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1003), .Y(n_999) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1007), .Y(n_1004) );
INVx4_ASAP7_75t_SL g1010 ( .A(n_1011), .Y(n_1010) );
XOR2x2_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1028), .Y(n_1011) );
NAND3x1_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1022), .C(n_1025), .Y(n_1012) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1017), .Y(n_1013) );
NAND3xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .C(n_1021), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1174 ( .A(n_1020), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_SL g1057 ( .A(n_1032), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1042), .Y(n_1032) );
NOR2xp33_ASAP7_75t_SL g1033 ( .A(n_1034), .B(n_1038), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1049), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1047), .Y(n_1043) );
NAND2xp5_ASAP7_75t_SL g1049 ( .A(n_1050), .B(n_1054), .Y(n_1049) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVxp67_ASAP7_75t_L g1186 ( .A(n_1053), .Y(n_1186) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1055), .Y(n_1191) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
AOI22xp5_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1062), .B1(n_1094), .B2(n_1125), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
AO22x1_ASAP7_75t_SL g1062 ( .A1(n_1063), .A2(n_1078), .B1(n_1092), .B2(n_1093), .Y(n_1062) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_1063), .Y(n_1092) );
XOR2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1077), .Y(n_1063) );
NAND4xp75_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1068), .C(n_1072), .D(n_1075), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
AND2x2_ASAP7_75t_SL g1068 ( .A(n_1069), .B(n_1070), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1074), .Y(n_1072) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_1078), .Y(n_1093) );
XOR2x2_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1091), .Y(n_1078) );
NAND4xp75_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1083), .C(n_1086), .D(n_1090), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1094), .Y(n_1125) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1095), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1113), .Y(n_1095) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1104), .Y(n_1096) );
OAI221xp5_ASAP7_75t_SL g1097 ( .A1(n_1098), .A2(n_1100), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
OAI221xp5_ASAP7_75t_SL g1104 ( .A1(n_1105), .A2(n_1107), .B1(n_1108), .B2(n_1109), .C(n_1110), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx3_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
NOR2xp33_ASAP7_75t_SL g1113 ( .A(n_1114), .B(n_1118), .Y(n_1113) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_1129), .Y(n_1128) );
NOR2x1_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1134), .Y(n_1129) );
OR2x2_ASAP7_75t_SL g1194 ( .A(n_1130), .B(n_1135), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1133), .Y(n_1130) );
CKINVDCx20_ASAP7_75t_R g1161 ( .A(n_1131), .Y(n_1161) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1132), .B(n_1163), .Y(n_1166) );
CKINVDCx16_ASAP7_75t_R g1163 ( .A(n_1133), .Y(n_1163) );
CKINVDCx20_ASAP7_75t_R g1134 ( .A(n_1135), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1140), .Y(n_1138) );
OAI322xp33_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1160), .A3(n_1162), .B1(n_1164), .B2(n_1167), .C1(n_1168), .C2(n_1192), .Y(n_1141) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AND4x1_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1149), .C(n_1154), .D(n_1158), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
CKINVDCx20_ASAP7_75t_R g1164 ( .A(n_1165), .Y(n_1164) );
XNOR2x1_ASAP7_75t_L g1168 ( .A(n_1167), .B(n_1169), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1179), .Y(n_1169) );
NOR3xp33_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1184), .C(n_1188), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1183), .Y(n_1180) );
CKINVDCx20_ASAP7_75t_R g1192 ( .A(n_1193), .Y(n_1192) );
CKINVDCx20_ASAP7_75t_R g1193 ( .A(n_1194), .Y(n_1193) );
endmodule