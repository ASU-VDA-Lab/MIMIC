module real_aes_6766_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g442 ( .A(n_0), .Y(n_442) );
INVx1_ASAP7_75t_L g481 ( .A(n_1), .Y(n_481) );
INVx1_ASAP7_75t_L g191 ( .A(n_2), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_3), .A2(n_79), .B1(n_749), .B2(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_3), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_4), .A2(n_39), .B1(n_147), .B2(n_497), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g171 ( .A1(n_5), .A2(n_128), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_6), .B(n_121), .Y(n_472) );
AND2x6_ASAP7_75t_L g133 ( .A(n_7), .B(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_8), .A2(n_230), .B(n_231), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_9), .B(n_40), .Y(n_443) );
INVx1_ASAP7_75t_L g178 ( .A(n_10), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_11), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
INVx1_ASAP7_75t_L g476 ( .A(n_13), .Y(n_476) );
INVx1_ASAP7_75t_L g236 ( .A(n_14), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_15), .B(n_159), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_16), .B(n_122), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_17), .Y(n_756) );
AO32x2_ASAP7_75t_L g505 ( .A1(n_18), .A2(n_121), .A3(n_156), .B1(n_459), .B2(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_19), .B(n_147), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_20), .B(n_142), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_21), .B(n_122), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_22), .A2(n_52), .B1(n_147), .B2(n_497), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_23), .B(n_128), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_24), .A2(n_76), .B1(n_147), .B2(n_159), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_25), .B(n_147), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_26), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_27), .A2(n_234), .B(n_235), .C(n_237), .Y(n_233) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_28), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_29), .B(n_180), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_30), .B(n_176), .Y(n_193) );
AOI222xp33_ASAP7_75t_SL g104 ( .A1(n_31), .A2(n_105), .B1(n_111), .B2(n_723), .C1(n_724), .C2(n_729), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_32), .A2(n_43), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_32), .Y(n_107) );
INVx1_ASAP7_75t_L g165 ( .A(n_33), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_34), .B(n_180), .Y(n_520) );
INVx2_ASAP7_75t_L g131 ( .A(n_35), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_36), .B(n_147), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_37), .B(n_180), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_38), .A2(n_133), .B(n_137), .C(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g163 ( .A(n_41), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_42), .B(n_176), .Y(n_246) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_43), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_44), .B(n_147), .Y(n_466) );
OAI22xp5_ASAP7_75t_SL g105 ( .A1(n_45), .A2(n_106), .B1(n_109), .B2(n_110), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_45), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_46), .A2(n_87), .B1(n_209), .B2(n_497), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_47), .B(n_147), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_48), .B(n_147), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g166 ( .A(n_49), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_50), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_51), .B(n_128), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_53), .A2(n_62), .B1(n_147), .B2(n_159), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_54), .A2(n_137), .B1(n_159), .B2(n_161), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_55), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_56), .B(n_147), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_57), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_58), .B(n_147), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_59), .A2(n_146), .B(n_175), .C(n_177), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_60), .Y(n_250) );
INVx1_ASAP7_75t_L g173 ( .A(n_61), .Y(n_173) );
INVx1_ASAP7_75t_L g134 ( .A(n_63), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_64), .B(n_147), .Y(n_482) );
INVx1_ASAP7_75t_L g125 ( .A(n_65), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_66), .Y(n_738) );
AO32x2_ASAP7_75t_L g500 ( .A1(n_67), .A2(n_121), .A3(n_216), .B1(n_459), .B2(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g539 ( .A(n_68), .Y(n_539) );
INVx1_ASAP7_75t_L g515 ( .A(n_69), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_SL g141 ( .A1(n_70), .A2(n_142), .B(n_143), .C(n_146), .Y(n_141) );
INVxp67_ASAP7_75t_L g144 ( .A(n_71), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_72), .B(n_159), .Y(n_516) );
INVx1_ASAP7_75t_L g737 ( .A(n_73), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_74), .Y(n_169) );
INVx1_ASAP7_75t_L g243 ( .A(n_75), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_77), .A2(n_133), .B(n_137), .C(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_78), .B(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_79), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_80), .B(n_159), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_81), .B(n_192), .Y(n_205) );
INVx2_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_83), .B(n_142), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_84), .B(n_159), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_85), .A2(n_133), .B(n_137), .C(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g440 ( .A(n_86), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g445 ( .A(n_86), .Y(n_445) );
OR2x2_ASAP7_75t_L g741 ( .A(n_86), .B(n_732), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_88), .A2(n_101), .B1(n_159), .B2(n_160), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_89), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_90), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_91), .A2(n_133), .B(n_137), .C(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_92), .Y(n_226) );
INVx1_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_94), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_95), .B(n_192), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_96), .B(n_159), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_97), .B(n_121), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_98), .A2(n_128), .B(n_135), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_99), .B(n_737), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_100), .A2(n_103), .B1(n_733), .B2(n_742), .C1(n_757), .C2(n_763), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_100), .A2(n_747), .B1(n_748), .B2(n_751), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_100), .Y(n_751) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g723 ( .A(n_105), .Y(n_723) );
INVx1_ASAP7_75t_L g109 ( .A(n_106), .Y(n_109) );
OAI22x1_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_438), .B1(n_444), .B2(n_446), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_112), .A2(n_113), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_113), .A2(n_725), .B1(n_726), .B2(n_728), .Y(n_724) );
AND2x2_ASAP7_75t_SL g113 ( .A(n_114), .B(n_375), .Y(n_113) );
NOR4xp25_ASAP7_75t_L g114 ( .A(n_115), .B(n_305), .C(n_336), .D(n_355), .Y(n_114) );
NAND4xp25_ASAP7_75t_L g115 ( .A(n_116), .B(n_263), .C(n_278), .D(n_296), .Y(n_115) );
AOI222xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_198), .B1(n_239), .B2(n_251), .C1(n_256), .C2(n_258), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_181), .Y(n_117) );
INVx1_ASAP7_75t_L g319 ( .A(n_118), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_152), .Y(n_118) );
AND2x2_ASAP7_75t_L g182 ( .A(n_119), .B(n_170), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_119), .B(n_185), .Y(n_348) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g255 ( .A(n_120), .B(n_154), .Y(n_255) );
AND2x2_ASAP7_75t_L g264 ( .A(n_120), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g290 ( .A(n_120), .Y(n_290) );
AND2x2_ASAP7_75t_L g311 ( .A(n_120), .B(n_154), .Y(n_311) );
BUFx2_ASAP7_75t_L g334 ( .A(n_120), .Y(n_334) );
AND2x2_ASAP7_75t_L g358 ( .A(n_120), .B(n_155), .Y(n_358) );
AND2x2_ASAP7_75t_L g422 ( .A(n_120), .B(n_170), .Y(n_422) );
OA21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_127), .B(n_149), .Y(n_120) );
INVx4_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_121), .A2(n_464), .B(n_472), .Y(n_463) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_123), .B(n_124), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
BUFx2_ASAP7_75t_L g230 ( .A(n_128), .Y(n_230) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_129), .B(n_133), .Y(n_167) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g471 ( .A(n_130), .Y(n_471) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g138 ( .A(n_131), .Y(n_138) );
INVx1_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
INVx1_ASAP7_75t_L g139 ( .A(n_132), .Y(n_139) );
INVx1_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
INVx3_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
INVx4_ASAP7_75t_SL g148 ( .A(n_133), .Y(n_148) );
BUFx3_ASAP7_75t_L g459 ( .A(n_133), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_133), .A2(n_465), .B(n_468), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_133), .A2(n_475), .B(n_479), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_133), .A2(n_490), .B(n_494), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_133), .A2(n_514), .B(n_517), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B(n_141), .C(n_148), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_136), .A2(n_148), .B(n_173), .C(n_174), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_136), .A2(n_148), .B(n_232), .C(n_233), .Y(n_231) );
INVx5_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_138), .Y(n_147) );
BUFx3_ASAP7_75t_L g209 ( .A(n_138), .Y(n_209) );
INVx1_ASAP7_75t_L g497 ( .A(n_138), .Y(n_497) );
INVx1_ASAP7_75t_L g493 ( .A(n_142), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_145), .B(n_178), .Y(n_177) );
INVx5_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g501 ( .A1(n_145), .A2(n_176), .B1(n_502), .B2(n_503), .Y(n_501) );
O2A1O1Ixp5_ASAP7_75t_SL g514 ( .A1(n_146), .A2(n_192), .B(n_515), .C(n_516), .Y(n_514) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g157 ( .A1(n_148), .A2(n_158), .B1(n_166), .B2(n_167), .Y(n_157) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_150), .A2(n_171), .B(n_179), .Y(n_170) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_151), .B(n_212), .Y(n_211) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_151), .B(n_455), .C(n_459), .Y(n_454) );
AO21x1_ASAP7_75t_L g547 ( .A1(n_151), .A2(n_455), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g323 ( .A(n_152), .B(n_254), .Y(n_323) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_153), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_170), .Y(n_153) );
OR2x2_ASAP7_75t_L g283 ( .A(n_154), .B(n_186), .Y(n_283) );
AND2x2_ASAP7_75t_L g295 ( .A(n_154), .B(n_254), .Y(n_295) );
BUFx2_ASAP7_75t_L g427 ( .A(n_154), .Y(n_427) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OR2x2_ASAP7_75t_L g184 ( .A(n_155), .B(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g277 ( .A(n_155), .B(n_186), .Y(n_277) );
AND2x2_ASAP7_75t_L g330 ( .A(n_155), .B(n_170), .Y(n_330) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_155), .Y(n_366) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_168), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_156), .B(n_169), .Y(n_168) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_156), .A2(n_187), .B(n_195), .Y(n_186) );
INVx2_ASAP7_75t_L g210 ( .A(n_156), .Y(n_210) );
INVx2_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g161 ( .A1(n_162), .A2(n_163), .B1(n_164), .B2(n_165), .Y(n_161) );
INVx2_ASAP7_75t_L g164 ( .A(n_162), .Y(n_164) );
INVx4_ASAP7_75t_L g234 ( .A(n_162), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_167), .A2(n_188), .B(n_189), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_167), .A2(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g253 ( .A(n_170), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_SL g265 ( .A(n_170), .Y(n_265) );
INVx2_ASAP7_75t_L g276 ( .A(n_170), .Y(n_276) );
BUFx2_ASAP7_75t_L g300 ( .A(n_170), .Y(n_300) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_170), .B(n_358), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_175), .A2(n_495), .B(n_496), .Y(n_494) );
O2A1O1Ixp5_ASAP7_75t_L g538 ( .A1(n_175), .A2(n_480), .B(n_539), .C(n_540), .Y(n_538) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g222 ( .A(n_176), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_176), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_176), .A2(n_457), .B1(n_507), .B2(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g197 ( .A(n_180), .Y(n_197) );
INVx2_ASAP7_75t_L g216 ( .A(n_180), .Y(n_216) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_180), .A2(n_229), .B(n_238), .Y(n_228) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_180), .A2(n_489), .B(n_498), .Y(n_488) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_180), .A2(n_513), .B(n_520), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
AOI332xp33_ASAP7_75t_L g278 ( .A1(n_182), .A2(n_279), .A3(n_283), .B1(n_284), .B2(n_288), .B3(n_291), .C1(n_292), .C2(n_294), .Y(n_278) );
NAND2x1_ASAP7_75t_L g363 ( .A(n_182), .B(n_254), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_182), .B(n_268), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_SL g296 ( .A1(n_183), .A2(n_297), .B(n_300), .C(n_301), .Y(n_296) );
AND2x2_ASAP7_75t_L g435 ( .A(n_183), .B(n_276), .Y(n_435) );
INVx3_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g332 ( .A(n_184), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g337 ( .A(n_184), .B(n_334), .Y(n_337) );
INVx1_ASAP7_75t_L g268 ( .A(n_185), .Y(n_268) );
AND2x2_ASAP7_75t_L g371 ( .A(n_185), .B(n_330), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_185), .B(n_311), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_185), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_185), .B(n_289), .Y(n_397) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx3_ASAP7_75t_L g254 ( .A(n_186), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .C(n_194), .Y(n_190) );
INVx2_ASAP7_75t_L g457 ( .A(n_192), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_192), .A2(n_466), .B(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_192), .A2(n_536), .B(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_194), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_197), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_197), .B(n_250), .Y(n_249) );
OAI31xp33_ASAP7_75t_L g436 ( .A1(n_198), .A2(n_357), .A3(n_364), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
AND2x2_ASAP7_75t_L g239 ( .A(n_199), .B(n_240), .Y(n_239) );
NAND2x1_ASAP7_75t_SL g259 ( .A(n_199), .B(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_199), .Y(n_346) );
AND2x2_ASAP7_75t_L g351 ( .A(n_199), .B(n_262), .Y(n_351) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_200), .A2(n_264), .B(n_266), .C(n_269), .Y(n_263) );
OR2x2_ASAP7_75t_L g280 ( .A(n_200), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g293 ( .A(n_200), .Y(n_293) );
AND2x2_ASAP7_75t_L g299 ( .A(n_200), .B(n_241), .Y(n_299) );
INVx2_ASAP7_75t_L g317 ( .A(n_200), .Y(n_317) );
AND2x2_ASAP7_75t_L g328 ( .A(n_200), .B(n_282), .Y(n_328) );
AND2x2_ASAP7_75t_L g360 ( .A(n_200), .B(n_318), .Y(n_360) );
AND2x2_ASAP7_75t_L g364 ( .A(n_200), .B(n_287), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_200), .B(n_213), .Y(n_369) );
AND2x2_ASAP7_75t_L g403 ( .A(n_200), .B(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_200), .B(n_306), .Y(n_437) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AOI21xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_203), .B(n_210), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_207), .A2(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g237 ( .A(n_209), .Y(n_237) );
INVx1_ASAP7_75t_L g248 ( .A(n_210), .Y(n_248) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_210), .A2(n_474), .B(n_483), .Y(n_473) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_210), .A2(n_534), .B(n_541), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_213), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g345 ( .A(n_213), .Y(n_345) );
AND2x2_ASAP7_75t_L g407 ( .A(n_213), .B(n_328), .Y(n_407) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_227), .Y(n_213) );
OR2x2_ASAP7_75t_L g261 ( .A(n_214), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g271 ( .A(n_214), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_214), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g379 ( .A(n_214), .Y(n_379) );
AND2x2_ASAP7_75t_L g396 ( .A(n_214), .B(n_241), .Y(n_396) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g287 ( .A(n_215), .B(n_227), .Y(n_287) );
AND2x2_ASAP7_75t_L g316 ( .A(n_215), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g327 ( .A(n_215), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_215), .B(n_282), .Y(n_418) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_225), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_224), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_223), .Y(n_219) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g240 ( .A(n_228), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g262 ( .A(n_228), .Y(n_262) );
AND2x2_ASAP7_75t_L g318 ( .A(n_228), .B(n_282), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_234), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g478 ( .A(n_234), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_234), .A2(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g420 ( .A(n_239), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_240), .Y(n_424) );
INVx2_ASAP7_75t_L g282 ( .A(n_241), .Y(n_282) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_248), .B(n_249), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_253), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_253), .B(n_358), .Y(n_416) );
OR2x2_ASAP7_75t_L g257 ( .A(n_254), .B(n_255), .Y(n_257) );
INVx1_ASAP7_75t_SL g309 ( .A(n_254), .Y(n_309) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_260), .A2(n_313), .B1(n_315), .B2(n_319), .C(n_320), .Y(n_312) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g340 ( .A(n_261), .B(n_304), .Y(n_340) );
INVx2_ASAP7_75t_L g272 ( .A(n_262), .Y(n_272) );
INVx1_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_262), .B(n_282), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_262), .B(n_285), .Y(n_392) );
INVx1_ASAP7_75t_L g400 ( .A(n_262), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_264), .B(n_268), .Y(n_314) );
AND2x4_ASAP7_75t_L g289 ( .A(n_265), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g402 ( .A(n_268), .B(n_358), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_271), .B(n_303), .Y(n_302) );
INVxp67_ASAP7_75t_L g410 ( .A(n_272), .Y(n_410) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g310 ( .A(n_276), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g382 ( .A(n_276), .B(n_358), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_276), .B(n_295), .Y(n_388) );
AOI322xp5_ASAP7_75t_L g342 ( .A1(n_277), .A2(n_311), .A3(n_318), .B1(n_343), .B2(n_346), .C1(n_347), .C2(n_349), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_277), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g408 ( .A(n_280), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g354 ( .A(n_281), .Y(n_354) );
INVx2_ASAP7_75t_L g285 ( .A(n_282), .Y(n_285) );
INVx1_ASAP7_75t_L g344 ( .A(n_282), .Y(n_344) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_283), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g380 ( .A(n_285), .B(n_293), .Y(n_380) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g292 ( .A(n_287), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g335 ( .A(n_287), .B(n_328), .Y(n_335) );
AND2x2_ASAP7_75t_L g339 ( .A(n_287), .B(n_299), .Y(n_339) );
OAI21xp33_ASAP7_75t_SL g349 ( .A1(n_288), .A2(n_350), .B(n_352), .Y(n_349) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_288), .A2(n_420), .B1(n_421), .B2(n_423), .Y(n_419) );
INVx3_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g294 ( .A(n_289), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_289), .B(n_309), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_291), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g431 ( .A(n_298), .Y(n_431) );
INVx4_ASAP7_75t_L g304 ( .A(n_299), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_299), .B(n_326), .Y(n_374) );
INVx1_ASAP7_75t_SL g386 ( .A(n_300), .Y(n_386) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_304), .B(n_400), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_307), .B(n_312), .C(n_329), .Y(n_305) );
OAI221xp5_ASAP7_75t_SL g425 ( .A1(n_307), .A2(n_345), .B1(n_424), .B2(n_426), .C(n_428), .Y(n_425) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_309), .B(n_422), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g401 ( .A1(n_310), .A2(n_387), .A3(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g391 ( .A(n_316), .Y(n_391) );
AND2x2_ASAP7_75t_L g404 ( .A(n_318), .B(n_327), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_328), .B(n_431), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI221xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_338), .B1(n_340), .B2(n_341), .C(n_342), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_337), .A2(n_406), .B(n_408), .C(n_411), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_340), .B(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g353 ( .A(n_351), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g395 ( .A(n_351), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B(n_361), .C(n_370), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_359), .A2(n_369), .B1(n_433), .B2(n_434), .C(n_436), .Y(n_432) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B1(n_365), .B2(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_372), .B(n_373), .Y(n_370) );
INVx1_ASAP7_75t_SL g433 ( .A(n_372), .Y(n_433) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NOR4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_405), .C(n_425), .D(n_432), .Y(n_375) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B(n_383), .C(n_401), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B(n_389), .C(n_393), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g412 ( .A(n_390), .Y(n_412) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
OR2x2_ASAP7_75t_L g423 ( .A(n_391), .B(n_424), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_415), .B2(n_417), .C(n_419), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_422), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g725 ( .A(n_439), .Y(n_725) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g444 ( .A(n_441), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g732 ( .A(n_441), .Y(n_732) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g727 ( .A(n_444), .Y(n_727) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_445), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g728 ( .A(n_446), .Y(n_728) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_448), .B(n_657), .Y(n_447) );
NOR5xp2_ASAP7_75t_L g448 ( .A(n_449), .B(n_570), .C(n_616), .D(n_629), .E(n_641), .Y(n_448) );
OAI211xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_484), .B(n_524), .C(n_551), .Y(n_449) );
INVx1_ASAP7_75t_SL g652 ( .A(n_450), .Y(n_652) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
AND2x2_ASAP7_75t_L g576 ( .A(n_451), .B(n_461), .Y(n_576) );
AND2x2_ASAP7_75t_L g604 ( .A(n_451), .B(n_550), .Y(n_604) );
AND2x2_ASAP7_75t_L g612 ( .A(n_451), .B(n_555), .Y(n_612) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g542 ( .A(n_452), .B(n_462), .Y(n_542) );
INVx2_ASAP7_75t_L g554 ( .A(n_452), .Y(n_554) );
AND2x2_ASAP7_75t_L g679 ( .A(n_452), .B(n_621), .Y(n_679) );
OR2x2_ASAP7_75t_L g681 ( .A(n_452), .B(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g548 ( .A(n_453), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_457), .A2(n_469), .B(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_457), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_459), .A2(n_535), .B(n_538), .Y(n_534) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g592 ( .A(n_461), .B(n_564), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_461), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g706 ( .A(n_461), .B(n_546), .Y(n_706) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
AND2x2_ASAP7_75t_L g549 ( .A(n_462), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g596 ( .A(n_462), .Y(n_596) );
AND2x2_ASAP7_75t_L g621 ( .A(n_462), .B(n_533), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_462), .B(n_654), .Y(n_691) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g555 ( .A(n_463), .B(n_533), .Y(n_555) );
AND2x2_ASAP7_75t_L g569 ( .A(n_463), .B(n_532), .Y(n_569) );
AND2x2_ASAP7_75t_L g586 ( .A(n_463), .B(n_473), .Y(n_586) );
AND2x2_ASAP7_75t_L g643 ( .A(n_463), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_463), .B(n_550), .Y(n_656) );
AND2x2_ASAP7_75t_L g708 ( .A(n_463), .B(n_633), .Y(n_708) );
INVx2_ASAP7_75t_L g480 ( .A(n_471), .Y(n_480) );
AND2x2_ASAP7_75t_L g531 ( .A(n_473), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g550 ( .A(n_473), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_473), .B(n_533), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_509), .B(n_521), .Y(n_484) );
INVx1_ASAP7_75t_SL g640 ( .A(n_485), .Y(n_640) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_499), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_SL g528 ( .A(n_487), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g523 ( .A(n_488), .Y(n_523) );
INVx1_ASAP7_75t_L g560 ( .A(n_488), .Y(n_560) );
AND2x2_ASAP7_75t_L g581 ( .A(n_488), .B(n_504), .Y(n_581) );
AND2x2_ASAP7_75t_L g615 ( .A(n_488), .B(n_505), .Y(n_615) );
OR2x2_ASAP7_75t_L g634 ( .A(n_488), .B(n_511), .Y(n_634) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_488), .Y(n_648) );
AND2x2_ASAP7_75t_L g661 ( .A(n_488), .B(n_662), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_493), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_499), .A2(n_583), .B1(n_584), .B2(n_593), .Y(n_582) );
AND2x2_ASAP7_75t_L g666 ( .A(n_499), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_504), .Y(n_499) );
INVx1_ASAP7_75t_L g527 ( .A(n_500), .Y(n_527) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_500), .Y(n_564) );
INVx1_ASAP7_75t_L g575 ( .A(n_500), .Y(n_575) );
AND2x2_ASAP7_75t_L g590 ( .A(n_500), .B(n_505), .Y(n_590) );
OR2x2_ASAP7_75t_L g544 ( .A(n_504), .B(n_529), .Y(n_544) );
AND2x2_ASAP7_75t_L g574 ( .A(n_504), .B(n_575), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g662 ( .A(n_504), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g522 ( .A(n_505), .B(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g631 ( .A(n_505), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_509), .B(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g609 ( .A(n_510), .B(n_575), .Y(n_609) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g521 ( .A(n_511), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g529 ( .A(n_512), .Y(n_529) );
OR2x2_ASAP7_75t_L g559 ( .A(n_512), .B(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_512), .Y(n_614) );
AOI32xp33_ASAP7_75t_L g651 ( .A1(n_521), .A2(n_581), .A3(n_652), .B1(n_653), .B2(n_655), .Y(n_651) );
AND2x2_ASAP7_75t_L g577 ( .A(n_522), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_522), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_522), .B(n_609), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_522), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_530), .B1(n_543), .B2(n_545), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
AND2x2_ASAP7_75t_L g630 ( .A(n_526), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_527), .B(n_529), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_528), .A2(n_552), .B1(n_556), .B2(n_566), .Y(n_551) );
AND2x2_ASAP7_75t_L g573 ( .A(n_528), .B(n_574), .Y(n_573) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_528), .A2(n_542), .B(n_590), .C(n_625), .Y(n_624) );
OAI332xp33_ASAP7_75t_L g629 ( .A1(n_528), .A2(n_630), .A3(n_632), .B1(n_634), .B2(n_635), .B3(n_637), .C1(n_638), .C2(n_640), .Y(n_629) );
INVx2_ASAP7_75t_L g670 ( .A(n_528), .Y(n_670) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_529), .Y(n_588) );
INVx1_ASAP7_75t_L g663 ( .A(n_529), .Y(n_663) );
AND2x2_ASAP7_75t_L g717 ( .A(n_529), .B(n_581), .Y(n_717) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .Y(n_530) );
AND2x2_ASAP7_75t_L g597 ( .A(n_532), .B(n_547), .Y(n_597) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g546 ( .A(n_533), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g645 ( .A(n_533), .B(n_547), .Y(n_645) );
INVx1_ASAP7_75t_L g654 ( .A(n_533), .Y(n_654) );
INVx1_ASAP7_75t_L g628 ( .A(n_542), .Y(n_628) );
INVxp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g712 ( .A(n_544), .B(n_564), .Y(n_712) );
INVx1_ASAP7_75t_SL g623 ( .A(n_545), .Y(n_623) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
AND2x2_ASAP7_75t_L g650 ( .A(n_546), .B(n_608), .Y(n_650) );
INVx1_ASAP7_75t_L g669 ( .A(n_546), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_546), .B(n_636), .Y(n_671) );
INVx1_ASAP7_75t_L g568 ( .A(n_547), .Y(n_568) );
AND2x2_ASAP7_75t_L g572 ( .A(n_549), .B(n_553), .Y(n_572) );
AND2x2_ASAP7_75t_L g639 ( .A(n_549), .B(n_597), .Y(n_639) );
INVx2_ASAP7_75t_L g682 ( .A(n_549), .Y(n_682) );
INVx2_ASAP7_75t_L g565 ( .A(n_550), .Y(n_565) );
AND2x2_ASAP7_75t_L g567 ( .A(n_550), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx1_ASAP7_75t_L g583 ( .A(n_553), .Y(n_583) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_554), .B(n_627), .Y(n_633) );
OR2x2_ASAP7_75t_L g697 ( .A(n_554), .B(n_656), .Y(n_697) );
INVx1_ASAP7_75t_L g721 ( .A(n_554), .Y(n_721) );
INVx1_ASAP7_75t_L g677 ( .A(n_555), .Y(n_677) );
AND2x2_ASAP7_75t_L g722 ( .A(n_555), .B(n_565), .Y(n_722) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_559), .A2(n_585), .B1(n_587), .B2(n_591), .Y(n_584) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI322xp33_ASAP7_75t_SL g668 ( .A1(n_562), .A2(n_669), .A3(n_670), .B1(n_671), .B2(n_672), .C1(n_675), .C2(n_677), .Y(n_668) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
AND2x2_ASAP7_75t_L g665 ( .A(n_563), .B(n_581), .Y(n_665) );
OR2x2_ASAP7_75t_L g699 ( .A(n_563), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g702 ( .A(n_563), .B(n_634), .Y(n_702) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g647 ( .A(n_564), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g703 ( .A(n_564), .B(n_634), .Y(n_703) );
INVx3_ASAP7_75t_L g636 ( .A(n_565), .Y(n_636) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g692 ( .A(n_567), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g571 ( .A1(n_569), .A2(n_572), .B1(n_573), .B2(n_576), .C1(n_577), .C2(n_579), .Y(n_571) );
INVx1_ASAP7_75t_L g602 ( .A(n_569), .Y(n_602) );
NAND3xp33_ASAP7_75t_SL g570 ( .A(n_571), .B(n_582), .C(n_599), .Y(n_570) );
AND2x2_ASAP7_75t_L g687 ( .A(n_574), .B(n_588), .Y(n_687) );
BUFx2_ASAP7_75t_L g578 ( .A(n_575), .Y(n_578) );
INVx1_ASAP7_75t_L g619 ( .A(n_575), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_576), .A2(n_612), .B1(n_665), .B2(n_666), .C(n_668), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_578), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_581), .Y(n_605) );
AND2x2_ASAP7_75t_L g618 ( .A(n_581), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_586), .B(n_597), .Y(n_598) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g593 ( .A1(n_588), .A2(n_594), .B(n_598), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_588), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g685 ( .A(n_590), .B(n_667), .Y(n_685) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g608 ( .A(n_596), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_597), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g714 ( .A(n_597), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_605), .B1(n_606), .B2(n_609), .C(n_610), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_601), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g710 ( .A(n_609), .B(n_615), .Y(n_710) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
OAI31xp33_ASAP7_75t_SL g678 ( .A1(n_613), .A2(n_652), .A3(n_679), .B(n_680), .Y(n_678) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g667 ( .A(n_614), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_615), .B(n_619), .Y(n_718) );
OAI221xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_620), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_616) );
INVx1_ASAP7_75t_L g622 ( .A(n_618), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_621), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g637 ( .A(n_630), .Y(n_637) );
INVx2_ASAP7_75t_L g673 ( .A(n_631), .Y(n_673) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g659 ( .A(n_636), .B(n_645), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g709 ( .A1(n_636), .A2(n_653), .B(n_710), .C(n_711), .Y(n_709) );
OAI221xp5_ASAP7_75t_SL g641 ( .A1(n_637), .A2(n_642), .B1(n_646), .B2(n_649), .C(n_651), .Y(n_641) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_640), .A2(n_705), .B(n_707), .C(n_709), .Y(n_704) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_643), .A2(n_694), .B1(n_696), .B2(n_698), .C(n_701), .Y(n_693) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
NOR4xp25_ASAP7_75t_L g657 ( .A(n_658), .B(n_683), .C(n_704), .D(n_715), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_660), .B(n_664), .C(n_678), .Y(n_658) );
INVx1_ASAP7_75t_SL g713 ( .A(n_665), .Y(n_713) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_SL g676 ( .A(n_674), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_681), .A2(n_690), .B1(n_702), .B2(n_703), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B(n_688), .C(n_693), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI31xp33_ASAP7_75t_L g715 ( .A1(n_686), .A2(n_716), .A3(n_718), .B(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_739), .Y(n_734) );
NOR2xp33_ASAP7_75t_SL g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_SL g762 ( .A(n_736), .Y(n_762) );
INVx1_ASAP7_75t_L g761 ( .A(n_738), .Y(n_761) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_738), .A2(n_762), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g753 ( .A(n_741), .Y(n_753) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_741), .Y(n_755) );
BUFx2_ASAP7_75t_L g765 ( .A(n_741), .Y(n_765) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_752), .B(n_754), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_SL g754 ( .A(n_755), .B(n_756), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
endmodule