module real_jpeg_12402_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_3),
.A2(n_35),
.B1(n_67),
.B2(n_68),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_3),
.A2(n_35),
.B1(n_62),
.B2(n_64),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_4),
.A2(n_62),
.B1(n_64),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_4),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_72),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_72),
.Y(n_216)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_40),
.B1(n_67),
.B2(n_68),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_6),
.A2(n_40),
.B1(n_62),
.B2(n_64),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_62),
.B1(n_64),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_113),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_113),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_9),
.A2(n_62),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_70),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_11),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_11),
.B(n_128),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_11),
.B(n_30),
.C(n_46),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_103),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_11),
.A2(n_27),
.B1(n_38),
.B2(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_11),
.B(n_109),
.Y(n_233)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_81),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_13),
.A2(n_62),
.B1(n_64),
.B2(n_81),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_81),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_14),
.A2(n_50),
.B1(n_67),
.B2(n_68),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_14),
.A2(n_50),
.B1(n_62),
.B2(n_64),
.Y(n_286)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_332),
.C(n_338),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_330),
.B(n_335),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_318),
.B(n_329),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_280),
.B(n_315),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_257),
.B(n_279),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_139),
.B(n_256),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_114),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_23),
.B(n_114),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_84),
.C(n_94),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_24),
.B(n_84),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_56),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_25),
.B(n_57),
.C(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_26),
.B(n_41),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_27),
.A2(n_38),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_27),
.A2(n_38),
.B1(n_214),
.B2(n_222),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_27),
.A2(n_89),
.B(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_28),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_28),
.A2(n_37),
.B(n_90),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_28),
.A2(n_32),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_30),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_29),
.B(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_32),
.B(n_90),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_38),
.A2(n_87),
.B(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_38),
.B(n_103),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_51),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_42),
.A2(n_47),
.B1(n_54),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_42),
.A2(n_54),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_42),
.B(n_103),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_42),
.A2(n_54),
.B1(n_186),
.B2(n_211),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_42),
.A2(n_54),
.B(n_150),
.Y(n_293)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_43),
.B(n_52),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_43),
.A2(n_53),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_43),
.B(n_197),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OA22x2_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_49),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_48),
.B(n_68),
.C(n_78),
.Y(n_182)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_49),
.A2(n_77),
.B(n_181),
.C(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_49),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_51),
.B(n_196),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_54),
.A2(n_93),
.B(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_54),
.A2(n_136),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_54),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_59),
.A2(n_66),
.B1(n_69),
.B2(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_59),
.A2(n_71),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_59),
.B(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_68),
.B(n_102),
.C(n_104),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_103),
.CON(n_102),
.SN(n_102)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_65),
.C(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_66),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_68),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

HAxp5_ASAP7_75t_SL g181 ( 
.A(n_68),
.B(n_103),
.CON(n_181),
.SN(n_181)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_80),
.B(n_82),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_75),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_75),
.A2(n_109),
.B1(n_158),
.B2(n_181),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_75),
.A2(n_109),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_75),
.A2(n_80),
.B(n_109),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_79),
.A2(n_106),
.B1(n_107),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_79),
.A2(n_107),
.B1(n_148),
.B2(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_82),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_94),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_105),
.C(n_110),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_95),
.A2(n_96),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_112),
.B1(n_128),
.B2(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_110),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_108),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_107),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_108),
.B(n_124),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_138),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_130),
.B2(n_131),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_116),
.B(n_131),
.C(n_138),
.Y(n_278)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_118),
.B(n_122),
.C(n_126),
.Y(n_260)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_123),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_127),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_128),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_128),
.A2(n_144),
.B1(n_286),
.B2(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_128),
.A2(n_129),
.B(n_144),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_129),
.A2(n_144),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_137),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_132),
.A2(n_133),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_133),
.B(n_135),
.Y(n_265)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_133),
.A2(n_265),
.B(n_268),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_135),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_169),
.B(n_251),
.C(n_255),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_162),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_162),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_152),
.C(n_155),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_142),
.B(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_146),
.C(n_151),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_144),
.A2(n_269),
.B(n_304),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_151),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_155),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_163),
.B(n_167),
.C(n_168),
.Y(n_252)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_245),
.B(n_250),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_200),
.B(n_244),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_188),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_174),
.B(n_188),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_183),
.C(n_184),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_175),
.A2(n_176),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_184),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_189),
.B(n_194),
.C(n_198),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_238),
.B(n_243),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_228),
.B(n_237),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_217),
.B(n_227),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_223),
.B(n_226),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_242),
.Y(n_243)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_249),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_278),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_278),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_263),
.C(n_272),
.Y(n_311)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_271),
.B2(n_272),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B(n_277),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_283),
.C(n_297),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_277),
.A2(n_283),
.B1(n_284),
.B2(n_314),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_310),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_298),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_288),
.B1(n_295),
.B2(n_296),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_290),
.C(n_293),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_295),
.B1(n_302),
.B2(n_308),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_294),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_294),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_303),
.C(n_307),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_299),
.C(n_308),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_309),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_320)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_324),
.C(n_326),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_334),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule