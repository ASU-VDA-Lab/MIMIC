module real_jpeg_26855_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_244;
wire n_128;
wire n_213;
wire n_167;
wire n_179;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g63 ( 
.A(n_0),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_1),
.Y(n_122)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_1),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_65),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_40),
.B1(n_61),
.B2(n_62),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_8),
.A2(n_11),
.B(n_62),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_9),
.A2(n_29),
.B1(n_61),
.B2(n_62),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_9),
.A2(n_29),
.B1(n_42),
.B2(n_44),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_32),
.B1(n_42),
.B2(n_44),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_11),
.A2(n_22),
.B(n_25),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_11),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_11),
.B(n_21),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_11),
.A2(n_42),
.B(n_50),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_11),
.B(n_41),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_106),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_105),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_16),
.B(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_66),
.C(n_74),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_17),
.B(n_66),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_35),
.B2(n_36),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_18),
.A2(n_19),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_18),
.A2(n_19),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_18),
.A2(n_19),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_18),
.B(n_225),
.C(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_38),
.C(n_52),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_19),
.B(n_126),
.C(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_26),
.B(n_30),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_33),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_21),
.A2(n_31),
.B1(n_33),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_22),
.A2(n_32),
.B(n_51),
.C(n_162),
.Y(n_161)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_24),
.A2(n_28),
.B(n_32),
.C(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_31),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_32),
.A2(n_42),
.B(n_59),
.C(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_32),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_32),
.B(n_60),
.Y(n_200)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B(n_45),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_39),
.A2(n_41),
.B1(n_48),
.B2(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_41),
.B(n_48),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_46),
.A2(n_71),
.B(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_53),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_60),
.B1(n_64),
.B2(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_56),
.A2(n_60),
.B1(n_87),
.B2(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_68),
.B(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_61),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_96),
.B1(n_97),
.B2(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_69),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_69),
.B(n_152),
.C(n_153),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_69),
.A2(n_114),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_72),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_74),
.A2(n_75),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_83),
.B(n_88),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_76),
.A2(n_84),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_76),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_76),
.A2(n_88),
.B1(n_89),
.B2(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_77),
.A2(n_80),
.B1(n_122),
.B2(n_139),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_79),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_83),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_84),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_86),
.A2(n_134),
.B(n_136),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_96),
.A2(n_97),
.B1(n_126),
.B2(n_147),
.Y(n_240)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_97),
.B(n_114),
.C(n_115),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_97),
.B(n_147),
.C(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_258),
.B(n_263),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_247),
.B(n_257),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_233),
.B(n_246),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_155),
.B(n_216),
.C(n_232),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_144),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_111),
.B(n_144),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_123),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_112),
.B(n_124),
.C(n_131),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_119),
.A2(n_150),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_119),
.B(n_200),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_119),
.B(n_175),
.C(n_187),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_122),
.B(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_126),
.A2(n_132),
.B1(n_133),
.B2(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_132),
.A2(n_133),
.B1(n_182),
.B2(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_132),
.B(n_138),
.Y(n_225)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_147),
.C(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_133),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_151),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_146),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_149),
.B(n_151),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_215),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_210),
.B(n_214),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_209),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_166),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_165),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_173),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_175),
.C(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_177),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_177),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_175),
.B(n_222),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_204),
.B(n_208),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_189),
.B(n_203),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_184),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B(n_202),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_199),
.B(n_201),
.Y(n_193)
);

INVx5_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_206),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_212),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_230),
.B2(n_231),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_224),
.C(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_230),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_242),
.C(n_245),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_248),
.B(n_249),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_255),
.B2(n_256),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_253),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_255),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);


endmodule