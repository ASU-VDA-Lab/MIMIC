module fake_jpeg_17796_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_43),
.Y(n_61)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_17),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_50),
.Y(n_82)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_53),
.B1(n_39),
.B2(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_64),
.B(n_24),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_29),
.B1(n_25),
.B2(n_32),
.Y(n_53)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_66),
.B1(n_18),
.B2(n_44),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_14),
.B1(n_16),
.B2(n_15),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_72),
.Y(n_103)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_31),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_90),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_84),
.B1(n_97),
.B2(n_50),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_81),
.B1(n_93),
.B2(n_64),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_77),
.B(n_75),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_34),
.B1(n_22),
.B2(n_20),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_37),
.B1(n_22),
.B2(n_20),
.Y(n_84)
);

NOR2x1_ASAP7_75t_R g121 ( 
.A(n_86),
.B(n_99),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_37),
.B1(n_24),
.B2(n_26),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_45),
.B(n_37),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_61),
.C(n_49),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_33),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_102),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_6),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_105),
.B(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_98),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_117),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_56),
.B1(n_55),
.B2(n_48),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_53),
.B1(n_57),
.B2(n_48),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_57),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_76),
.C(n_93),
.Y(n_144)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_7),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_48),
.B1(n_37),
.B2(n_58),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_7),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_26),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx6p67_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_77),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_83),
.B1(n_79),
.B2(n_88),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_121),
.B(n_111),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_139),
.B(n_150),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_107),
.B(n_120),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_74),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_144),
.C(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_108),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_90),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_154),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_83),
.B1(n_70),
.B2(n_96),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_24),
.B1(n_62),
.B2(n_122),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_27),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_91),
.B(n_80),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_40),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_91),
.B(n_80),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_157),
.B(n_27),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_71),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_62),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_70),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_33),
.C(n_87),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_123),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_170),
.B(n_180),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_108),
.B1(n_89),
.B2(n_91),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_176),
.B1(n_183),
.B2(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_26),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_174),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_91),
.B(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_177),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_173),
.B(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_26),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_40),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_87),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_157),
.B1(n_152),
.B2(n_129),
.Y(n_192)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_26),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_28),
.B(n_30),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_134),
.B(n_26),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_188),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_28),
.B(n_30),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_33),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_33),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_33),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_195),
.B1(n_179),
.B2(n_190),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_148),
.B1(n_156),
.B2(n_147),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_177),
.B(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_141),
.C(n_157),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_198),
.C(n_217),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_43),
.C(n_40),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_185),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_205),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_164),
.B1(n_179),
.B2(n_178),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_28),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_196),
.Y(n_228)
);

XNOR2x2_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_180),
.Y(n_224)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_132),
.A3(n_33),
.B1(n_24),
.B2(n_40),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_211),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_132),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_216),
.B1(n_162),
.B2(n_188),
.Y(n_239)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

NOR4xp25_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_132),
.C(n_62),
.D(n_43),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_183),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_237),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_227),
.B1(n_230),
.B2(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_160),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_217),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_195),
.B1(n_213),
.B2(n_192),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_175),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_232),
.C(n_241),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_176),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_167),
.B1(n_173),
.B2(n_161),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_187),
.B1(n_174),
.B2(n_169),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_238),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_212),
.B1(n_193),
.B2(n_207),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_216),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_242),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_167),
.C(n_162),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_189),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_260),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_202),
.C(n_206),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_251),
.C(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_241),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_202),
.C(n_210),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_163),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_207),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_257),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_186),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_204),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_227),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_186),
.C(n_163),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_233),
.B1(n_214),
.B2(n_223),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_271),
.B1(n_273),
.B2(n_7),
.Y(n_290)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_247),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_256),
.B1(n_254),
.B2(n_214),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_235),
.C(n_223),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_43),
.C(n_38),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_224),
.B1(n_225),
.B2(n_231),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_122),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_11),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_260),
.B1(n_244),
.B2(n_255),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_10),
.B1(n_15),
.B2(n_3),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_287),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_288),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_245),
.B(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_289),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_122),
.B1(n_1),
.B2(n_2),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_282),
.A2(n_1),
.B1(n_2),
.B2(n_62),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_266),
.C(n_274),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_263),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_0),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_10),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_5),
.B1(n_13),
.B2(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_300),
.B1(n_282),
.B2(n_284),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_277),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_288),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_12),
.B(n_13),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_289),
.B(n_5),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_286),
.B1(n_287),
.B2(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_302),
.C(n_294),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_304),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_294),
.A3(n_297),
.B1(n_298),
.B2(n_296),
.C1(n_43),
.C2(n_5),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_310),
.A3(n_311),
.B1(n_312),
.B2(n_4),
.C1(n_38),
.C2(n_222),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_297),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_62),
.A3(n_3),
.B1(n_4),
.B2(n_2),
.C1(n_1),
.C2(n_38),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_307),
.B(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_38),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);


endmodule