module real_aes_1439_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_0), .B(n_117), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_1), .A2(n_126), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_2), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_3), .B(n_117), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_4), .B(n_133), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_5), .B(n_133), .Y(n_529) );
INVx1_ASAP7_75t_L g124 ( .A(n_6), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_7), .B(n_133), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_8), .Y(n_464) );
NAND2xp33_ASAP7_75t_L g510 ( .A(n_9), .B(n_135), .Y(n_510) );
AND2x2_ASAP7_75t_L g153 ( .A(n_10), .B(n_142), .Y(n_153) );
AND2x2_ASAP7_75t_L g162 ( .A(n_11), .B(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g139 ( .A(n_12), .Y(n_139) );
AOI221x1_ASAP7_75t_L g551 ( .A1(n_13), .A2(n_25), .B1(n_117), .B2(n_126), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_14), .B(n_133), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_15), .B(n_460), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_16), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_17), .B(n_117), .Y(n_506) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_18), .A2(n_142), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_19), .B(n_137), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_20), .B(n_133), .Y(n_489) );
AO21x1_ASAP7_75t_L g524 ( .A1(n_21), .A2(n_117), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_22), .B(n_117), .Y(n_187) );
INVx1_ASAP7_75t_L g457 ( .A(n_23), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_24), .A2(n_92), .B1(n_117), .B2(n_226), .Y(n_225) );
NAND2x1_ASAP7_75t_L g538 ( .A(n_26), .B(n_133), .Y(n_538) );
NAND2x1_ASAP7_75t_L g499 ( .A(n_27), .B(n_135), .Y(n_499) );
OR2x2_ASAP7_75t_L g140 ( .A(n_28), .B(n_89), .Y(n_140) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_28), .A2(n_89), .B(n_139), .Y(n_143) );
OAI22x1_ASAP7_75t_R g444 ( .A1(n_29), .A2(n_445), .B1(n_446), .B2(n_449), .Y(n_444) );
INVx1_ASAP7_75t_L g449 ( .A(n_29), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_30), .B(n_135), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_31), .B(n_133), .Y(n_509) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_32), .A2(n_163), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_33), .B(n_135), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_34), .A2(n_126), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g777 ( .A(n_35), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_36), .B(n_133), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_37), .A2(n_126), .B(n_570), .Y(n_569) );
XNOR2x2_ASAP7_75t_SL g470 ( .A(n_38), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g123 ( .A(n_39), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g127 ( .A(n_39), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g234 ( .A(n_39), .Y(n_234) );
OR2x6_ASAP7_75t_L g455 ( .A(n_40), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_41), .B(n_117), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_42), .B(n_117), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_43), .B(n_133), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_44), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_45), .B(n_135), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_46), .B(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_47), .A2(n_126), .B(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_48), .A2(n_126), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_49), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_50), .B(n_135), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_51), .B(n_117), .Y(n_169) );
INVx1_ASAP7_75t_L g120 ( .A(n_52), .Y(n_120) );
INVx1_ASAP7_75t_L g130 ( .A(n_52), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_53), .A2(n_68), .B1(n_447), .B2(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_53), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_54), .B(n_133), .Y(n_160) );
AND2x2_ASAP7_75t_L g198 ( .A(n_55), .B(n_137), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_56), .B(n_135), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_57), .B(n_133), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_58), .B(n_135), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_59), .A2(n_126), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_60), .B(n_117), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_61), .B(n_117), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_62), .A2(n_126), .B(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g193 ( .A(n_63), .B(n_138), .Y(n_193) );
AO21x1_ASAP7_75t_L g526 ( .A1(n_64), .A2(n_126), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_65), .B(n_117), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_66), .A2(n_84), .B1(n_472), .B2(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_66), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_67), .B(n_135), .Y(n_204) );
INVx1_ASAP7_75t_L g448 ( .A(n_68), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_69), .B(n_117), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_70), .B(n_135), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_71), .A2(n_97), .B1(n_126), .B2(n_232), .Y(n_231) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_72), .A2(n_104), .B1(n_461), .B2(n_466), .C1(n_780), .C2(n_784), .Y(n_103) );
XNOR2xp5_ASAP7_75t_L g105 ( .A(n_72), .B(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g574 ( .A(n_72), .B(n_138), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_73), .B(n_133), .Y(n_190) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
INVx1_ASAP7_75t_L g128 ( .A(n_74), .Y(n_128) );
AND2x2_ASAP7_75t_L g502 ( .A(n_75), .B(n_163), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_76), .B(n_135), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_77), .A2(n_126), .B(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_78), .A2(n_126), .B(n_131), .Y(n_125) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_79), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_80), .A2(n_126), .B(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g184 ( .A(n_81), .B(n_138), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_82), .B(n_137), .Y(n_223) );
INVx1_ASAP7_75t_L g458 ( .A(n_83), .Y(n_458) );
INVx1_ASAP7_75t_L g473 ( .A(n_84), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_85), .B(n_117), .Y(n_491) );
AND2x2_ASAP7_75t_L g512 ( .A(n_86), .B(n_163), .Y(n_512) );
AND2x2_ASAP7_75t_L g141 ( .A(n_87), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g525 ( .A(n_88), .B(n_174), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_90), .B(n_135), .Y(n_490) );
AND2x2_ASAP7_75t_L g541 ( .A(n_91), .B(n_163), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_93), .B(n_133), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_94), .A2(n_126), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_95), .B(n_135), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_96), .A2(n_126), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_98), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_99), .B(n_133), .Y(n_517) );
BUFx2_ASAP7_75t_L g192 ( .A(n_100), .Y(n_192) );
BUFx2_ASAP7_75t_L g465 ( .A(n_101), .Y(n_465) );
BUFx2_ASAP7_75t_SL g788 ( .A(n_101), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_102), .A2(n_126), .B(n_508), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_450), .B(n_459), .Y(n_104) );
OAI22x1_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_108), .B1(n_443), .B2(n_444), .Y(n_106) );
INVx5_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_108), .A2(n_475), .B1(n_477), .B2(n_768), .Y(n_474) );
INVx1_ASAP7_75t_L g773 ( .A(n_108), .Y(n_773) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_347), .Y(n_108) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_272), .C(n_308), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_246), .Y(n_110) );
AOI211xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_164), .B(n_194), .C(n_219), .Y(n_111) );
AND2x2_ASAP7_75t_L g337 ( .A(n_112), .B(n_196), .Y(n_337) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_144), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_113), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g370 ( .A(n_113), .B(n_252), .Y(n_370) );
AND2x2_ASAP7_75t_L g386 ( .A(n_113), .B(n_211), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_113), .B(n_396), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_113), .B(n_420), .Y(n_419) );
INVx4_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_SL g206 ( .A(n_114), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g241 ( .A(n_114), .Y(n_241) );
AND2x2_ASAP7_75t_L g288 ( .A(n_114), .B(n_221), .Y(n_288) );
AND2x2_ASAP7_75t_L g307 ( .A(n_114), .B(n_144), .Y(n_307) );
BUFx2_ASAP7_75t_L g312 ( .A(n_114), .Y(n_312) );
AND2x2_ASAP7_75t_L g356 ( .A(n_114), .B(n_154), .Y(n_356) );
AND2x4_ASAP7_75t_L g428 ( .A(n_114), .B(n_429), .Y(n_428) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_114), .B(n_210), .Y(n_440) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_141), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_125), .B(n_137), .Y(n_115) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_123), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
AND2x6_ASAP7_75t_L g135 ( .A(n_119), .B(n_128), .Y(n_135) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g133 ( .A(n_121), .B(n_130), .Y(n_133) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx5_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
AND2x2_ASAP7_75t_L g129 ( .A(n_124), .B(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_124), .Y(n_229) );
AND2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
BUFx3_ASAP7_75t_L g230 ( .A(n_127), .Y(n_230) );
INVx2_ASAP7_75t_L g236 ( .A(n_128), .Y(n_236) );
AND2x4_ASAP7_75t_L g232 ( .A(n_129), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g228 ( .A(n_130), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_134), .B(n_136), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_135), .B(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_136), .A2(n_150), .B(n_151), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_136), .A2(n_159), .B(n_160), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_136), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_136), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_136), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_136), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_136), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_136), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_136), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_136), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_136), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_136), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_136), .A2(n_553), .B(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_136), .A2(n_571), .B(n_572), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_137), .Y(n_146) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_137), .A2(n_225), .B(n_231), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_137), .A2(n_514), .B(n_515), .Y(n_513) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_137), .A2(n_551), .B(n_555), .Y(n_550) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_137), .A2(n_551), .B(n_555), .Y(n_562) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g174 ( .A(n_139), .B(n_140), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_142), .A2(n_187), .B(n_188), .Y(n_186) );
BUFx4f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx3_ASAP7_75t_L g155 ( .A(n_143), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_144), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g359 ( .A(n_144), .Y(n_359) );
BUFx2_ASAP7_75t_L g408 ( .A(n_144), .Y(n_408) );
INVx1_ASAP7_75t_L g430 ( .A(n_144), .Y(n_430) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_154), .Y(n_144) );
INVx3_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_145), .Y(n_396) );
AOI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_153), .Y(n_145) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_146), .A2(n_496), .B(n_502), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
INVx2_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_154), .B(n_207), .Y(n_211) );
INVx2_ASAP7_75t_L g296 ( .A(n_154), .Y(n_296) );
OR2x2_ASAP7_75t_L g303 ( .A(n_154), .B(n_252), .Y(n_303) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_162), .Y(n_154) );
INVx4_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_161), .Y(n_156) );
INVx3_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
AND2x2_ASAP7_75t_L g258 ( .A(n_164), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g292 ( .A(n_164), .B(n_255), .Y(n_292) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_175), .Y(n_164) );
AND2x2_ASAP7_75t_L g328 ( .A(n_165), .B(n_217), .Y(n_328) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g285 ( .A(n_166), .B(n_176), .Y(n_285) );
AND2x2_ASAP7_75t_L g404 ( .A(n_166), .B(n_185), .Y(n_404) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
INVx1_ASAP7_75t_L g244 ( .A(n_167), .Y(n_244) );
AND2x2_ASAP7_75t_L g300 ( .A(n_167), .B(n_176), .Y(n_300) );
AND2x2_ASAP7_75t_L g305 ( .A(n_167), .B(n_197), .Y(n_305) );
OR2x2_ASAP7_75t_L g368 ( .A(n_167), .B(n_185), .Y(n_368) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_167), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_174), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_174), .A2(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_SL g485 ( .A(n_174), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_174), .A2(n_506), .B(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_174), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g196 ( .A(n_175), .B(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g245 ( .A(n_175), .Y(n_245) );
NOR2x1_ASAP7_75t_SL g175 ( .A(n_176), .B(n_185), .Y(n_175) );
AO21x1_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_178), .B(n_184), .Y(n_176) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_177), .A2(n_178), .B(n_184), .Y(n_218) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_177), .A2(n_535), .B(n_541), .Y(n_534) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_177), .A2(n_568), .B(n_574), .Y(n_567) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_177), .A2(n_568), .B(n_574), .Y(n_603) );
AO21x2_ASAP7_75t_L g606 ( .A1(n_177), .A2(n_535), .B(n_541), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_183), .Y(n_178) );
AND2x2_ASAP7_75t_L g213 ( .A(n_185), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_SL g271 ( .A(n_185), .Y(n_271) );
NAND2x1_ASAP7_75t_L g281 ( .A(n_185), .B(n_197), .Y(n_281) );
OR2x2_ASAP7_75t_L g286 ( .A(n_185), .B(n_214), .Y(n_286) );
BUFx2_ASAP7_75t_L g342 ( .A(n_185), .Y(n_342) );
AND2x2_ASAP7_75t_L g378 ( .A(n_185), .B(n_257), .Y(n_378) );
AND2x2_ASAP7_75t_L g389 ( .A(n_185), .B(n_217), .Y(n_389) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_193), .Y(n_185) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_205), .B1(n_211), .B2(n_212), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_196), .A2(n_386), .B1(n_436), .B2(n_441), .Y(n_435) );
INVx4_ASAP7_75t_L g214 ( .A(n_197), .Y(n_214) );
INVx2_ASAP7_75t_L g255 ( .A(n_197), .Y(n_255) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_197), .Y(n_326) );
OR2x2_ASAP7_75t_L g341 ( .A(n_197), .B(n_217), .Y(n_341) );
OR2x2_ASAP7_75t_SL g367 ( .A(n_197), .B(n_368), .Y(n_367) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_206), .B(n_208), .Y(n_205) );
INVx2_ASAP7_75t_SL g248 ( .A(n_206), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_206), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g316 ( .A(n_206), .B(n_264), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_206), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g238 ( .A(n_207), .Y(n_238) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
AND2x2_ASAP7_75t_L g319 ( .A(n_207), .B(n_296), .Y(n_319) );
INVx1_ASAP7_75t_L g429 ( .A(n_207), .Y(n_429) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_209), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_209), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g237 ( .A(n_210), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_211), .B(n_370), .Y(n_369) );
AOI321xp33_ASAP7_75t_L g391 ( .A1(n_212), .A2(n_293), .A3(n_361), .B1(n_392), .B2(n_393), .C(n_397), .Y(n_391) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_215), .Y(n_212) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_213), .Y(n_290) );
AND2x2_ASAP7_75t_L g315 ( .A(n_213), .B(n_244), .Y(n_315) );
AND2x2_ASAP7_75t_L g390 ( .A(n_213), .B(n_300), .Y(n_390) );
INVx1_ASAP7_75t_L g259 ( .A(n_214), .Y(n_259) );
BUFx2_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
NOR2xp67_ASAP7_75t_L g376 ( .A(n_214), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g314 ( .A(n_215), .Y(n_314) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
BUFx2_ASAP7_75t_L g321 ( .A(n_216), .Y(n_321) );
INVx2_ASAP7_75t_L g257 ( .A(n_217), .Y(n_257) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_217), .Y(n_280) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AOI21xp33_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_239), .B(n_242), .Y(n_219) );
NOR2xp67_ASAP7_75t_L g373 ( .A(n_220), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_237), .Y(n_221) );
INVx3_ASAP7_75t_L g264 ( .A(n_222), .Y(n_264) );
AND2x2_ASAP7_75t_L g295 ( .A(n_222), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
AND2x4_ASAP7_75t_L g252 ( .A(n_223), .B(n_224), .Y(n_252) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_230), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
NOR2x1p5_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g335 ( .A(n_237), .Y(n_335) );
INVx1_ASAP7_75t_SL g420 ( .A(n_238), .Y(n_420) );
INVxp33_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_241), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g346 ( .A(n_241), .B(n_303), .Y(n_346) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_245), .Y(n_242) );
AND2x2_ASAP7_75t_L g350 ( .A(n_243), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_243), .B(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_244), .B(n_281), .Y(n_336) );
NOR4xp25_ASAP7_75t_L g431 ( .A(n_244), .B(n_275), .C(n_432), .D(n_433), .Y(n_431) );
OR2x2_ASAP7_75t_L g399 ( .A(n_245), .B(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_253), .B1(n_258), .B2(n_260), .C(n_265), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_L g274 ( .A(n_249), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g311 ( .A(n_250), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g331 ( .A(n_251), .Y(n_331) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
BUFx3_ASAP7_75t_L g354 ( .A(n_252), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_252), .B(n_362), .Y(n_361) );
INVxp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OR2x2_ASAP7_75t_L g298 ( .A(n_255), .B(n_299), .Y(n_298) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_257), .B(n_271), .Y(n_270) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
INVx2_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_262), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g267 ( .A(n_264), .Y(n_267) );
OAI321xp33_ASAP7_75t_L g379 ( .A1(n_264), .A2(n_372), .A3(n_380), .B1(n_385), .B2(n_387), .C(n_391), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
OR2x2_ASAP7_75t_L g334 ( .A(n_267), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g434 ( .A(n_270), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_271), .B(n_314), .Y(n_313) );
NAND2xp33_ASAP7_75t_SL g414 ( .A(n_271), .B(n_285), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_287), .C(n_291), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2x1_ASAP7_75t_L g276 ( .A(n_277), .B(n_282), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g383 ( .A(n_280), .Y(n_383) );
INVx3_ASAP7_75t_L g322 ( .A(n_281), .Y(n_322) );
OR2x2_ASAP7_75t_L g425 ( .A(n_281), .B(n_299), .Y(n_425) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_283), .A2(n_367), .B1(n_369), .B2(n_371), .Y(n_366) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_SL g365 ( .A(n_286), .Y(n_365) );
OR2x2_ASAP7_75t_L g442 ( .A(n_286), .B(n_299), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI21xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_293), .B(n_297), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_295), .B(n_312), .Y(n_411) );
AND2x2_ASAP7_75t_L g417 ( .A(n_295), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g362 ( .A(n_296), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_304), .B2(n_306), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_299), .A2(n_342), .B(n_344), .C(n_346), .Y(n_343) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_302), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_302), .B(n_394), .Y(n_416) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g388 ( .A(n_305), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_307), .A2(n_339), .B(n_342), .C(n_343), .Y(n_338) );
NAND3xp33_ASAP7_75t_SL g308 ( .A(n_309), .B(n_323), .C(n_338), .Y(n_308) );
AOI222xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .B1(n_315), .B2(n_316), .C1(n_317), .C2(n_320), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g372 ( .A(n_312), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_312), .B(n_345), .Y(n_398) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g332 ( .A(n_319), .Y(n_332) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
OR2x2_ASAP7_75t_L g437 ( .A(n_321), .B(n_354), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_322), .A2(n_413), .B1(n_415), .B2(n_417), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_329), .B1(n_333), .B2(n_336), .C(n_337), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI21xp5_ASAP7_75t_SL g397 ( .A1(n_330), .A2(n_398), .B(n_399), .Y(n_397) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx2_ASAP7_75t_L g345 ( .A(n_331), .Y(n_345) );
AND2x2_ASAP7_75t_L g439 ( .A(n_331), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g423 ( .A(n_335), .Y(n_423) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g352 ( .A(n_341), .B(n_342), .Y(n_352) );
INVx1_ASAP7_75t_L g405 ( .A(n_341), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_379), .C(n_401), .Y(n_347) );
OAI211xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B(n_355), .C(n_360), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_350), .A2(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI211xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B(n_366), .C(n_373), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g384 ( .A(n_367), .Y(n_384) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_368), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_370), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g432 ( .A(n_370), .Y(n_432) );
AND2x2_ASAP7_75t_L g422 ( .A(n_372), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g392 ( .A(n_374), .Y(n_392) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g400 ( .A(n_376), .Y(n_400) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_388), .A2(n_422), .B1(n_424), .B2(n_426), .C(n_431), .Y(n_421) );
OAI21xp33_ASAP7_75t_SL g436 ( .A1(n_393), .A2(n_437), .B(n_438), .Y(n_436) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_402), .B(n_412), .C(n_421), .D(n_435), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_406), .B1(n_409), .B2(n_410), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_430), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g460 ( .A(n_451), .Y(n_460) );
AND2x2_ASAP7_75t_L g780 ( .A(n_451), .B(n_781), .Y(n_780) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g790 ( .A(n_452), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x6_ASAP7_75t_SL g476 ( .A(n_453), .B(n_455), .Y(n_476) );
OR2x6_ASAP7_75t_SL g770 ( .A(n_453), .B(n_454), .Y(n_770) );
OR2x2_ASAP7_75t_L g779 ( .A(n_453), .B(n_455), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_SL g462 ( .A(n_463), .B(n_465), .Y(n_462) );
INVx2_ASAP7_75t_L g783 ( .A(n_463), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_463), .A2(n_786), .B(n_789), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g782 ( .A(n_465), .B(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_771), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_474), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI21xp33_ASAP7_75t_L g771 ( .A1(n_469), .A2(n_772), .B(n_776), .Y(n_771) );
INVx3_ASAP7_75t_SL g775 ( .A(n_475), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_478), .A2(n_770), .B1(n_773), .B2(n_774), .Y(n_772) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_666), .Y(n_478) );
NAND3xp33_ASAP7_75t_SL g479 ( .A(n_480), .B(n_578), .C(n_633), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_519), .B1(n_542), .B2(n_546), .C(n_556), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_503), .Y(n_481) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_482), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g577 ( .A(n_482), .Y(n_577) );
AND2x2_ASAP7_75t_L g622 ( .A(n_482), .B(n_559), .Y(n_622) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g610 ( .A(n_484), .Y(n_610) );
INVx1_ASAP7_75t_L g620 ( .A(n_484), .Y(n_620) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_492), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_485), .B(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_485), .A2(n_486), .B(n_492), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_491), .Y(n_486) );
OR2x2_ASAP7_75t_L g599 ( .A(n_494), .B(n_504), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_494), .B(n_545), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_494), .B(n_511), .Y(n_643) );
INVx2_ASAP7_75t_L g652 ( .A(n_494), .Y(n_652) );
AND2x2_ASAP7_75t_L g673 ( .A(n_494), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g757 ( .A(n_494), .B(n_576), .Y(n_757) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g585 ( .A(n_495), .B(n_511), .Y(n_585) );
AND2x2_ASAP7_75t_L g718 ( .A(n_495), .B(n_545), .Y(n_718) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_495), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
AND2x4_ASAP7_75t_L g672 ( .A(n_503), .B(n_673), .Y(n_672) );
AOI321xp33_ASAP7_75t_L g686 ( .A1(n_503), .A2(n_615), .A3(n_616), .B1(n_648), .B2(n_687), .C(n_690), .Y(n_686) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_511), .Y(n_503) );
BUFx3_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
INVx2_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_504), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g609 ( .A(n_504), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g642 ( .A(n_504), .Y(n_642) );
INVx5_ASAP7_75t_L g545 ( .A(n_511), .Y(n_545) );
NOR2x1_ASAP7_75t_SL g594 ( .A(n_511), .B(n_584), .Y(n_594) );
BUFx2_ASAP7_75t_L g689 ( .A(n_511), .Y(n_689) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVxp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
NOR2xp33_ASAP7_75t_SL g587 ( .A(n_521), .B(n_588), .Y(n_587) );
NOR4xp25_ASAP7_75t_L g690 ( .A(n_521), .B(n_684), .C(n_688), .D(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g728 ( .A(n_521), .Y(n_728) );
AND2x2_ASAP7_75t_L g762 ( .A(n_521), .B(n_702), .Y(n_762) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g563 ( .A(n_522), .Y(n_563) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g617 ( .A(n_523), .Y(n_617) );
OAI21x1_ASAP7_75t_SL g523 ( .A1(n_524), .A2(n_526), .B(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g531 ( .A(n_525), .Y(n_531) );
AOI33xp33_ASAP7_75t_L g758 ( .A1(n_532), .A2(n_560), .A3(n_591), .B1(n_607), .B2(n_713), .B3(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g548 ( .A(n_533), .B(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g558 ( .A(n_533), .B(n_559), .Y(n_558) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g565 ( .A(n_534), .Y(n_565) );
INVxp67_ASAP7_75t_L g646 ( .A(n_534), .Y(n_646) );
AND2x2_ASAP7_75t_L g702 ( .A(n_534), .B(n_567), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_540), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_542), .A2(n_724), .B(n_725), .Y(n_723) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_L g711 ( .A(n_543), .B(n_585), .Y(n_711) );
AND3x2_ASAP7_75t_L g713 ( .A(n_543), .B(n_597), .C(n_652), .Y(n_713) );
INVx3_ASAP7_75t_SL g665 ( .A(n_544), .Y(n_665) );
INVx4_ASAP7_75t_L g559 ( .A(n_545), .Y(n_559) );
AND2x2_ASAP7_75t_L g597 ( .A(n_545), .B(n_584), .Y(n_597) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g591 ( .A(n_549), .Y(n_591) );
AND2x4_ASAP7_75t_L g616 ( .A(n_549), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g679 ( .A(n_549), .B(n_567), .Y(n_679) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g649 ( .A(n_550), .Y(n_649) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_550), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_R g556 ( .A1(n_557), .A2(n_560), .B(n_564), .C(n_575), .Y(n_556) );
CKINVDCx16_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g608 ( .A(n_559), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_559), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_559), .B(n_576), .Y(n_737) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g719 ( .A(n_561), .B(n_709), .Y(n_719) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g566 ( .A(n_562), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g588 ( .A(n_562), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g604 ( .A(n_562), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g637 ( .A(n_562), .B(n_617), .Y(n_637) );
AND2x4_ASAP7_75t_L g602 ( .A(n_563), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g626 ( .A(n_563), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g664 ( .A(n_563), .B(n_589), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g592 ( .A(n_565), .B(n_589), .Y(n_592) );
AND2x2_ASAP7_75t_L g607 ( .A(n_565), .B(n_567), .Y(n_607) );
BUFx2_ASAP7_75t_L g663 ( .A(n_565), .Y(n_663) );
AND2x2_ASAP7_75t_L g677 ( .A(n_565), .B(n_588), .Y(n_677) );
INVx2_ASAP7_75t_L g589 ( .A(n_567), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_573), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_575), .A2(n_626), .B1(n_628), .B2(n_632), .Y(n_625) );
INVx2_ASAP7_75t_SL g656 ( .A(n_575), .Y(n_656) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g631 ( .A(n_576), .B(n_584), .Y(n_631) );
INVx1_ASAP7_75t_L g738 ( .A(n_577), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_611), .C(n_625), .Y(n_578) );
OAI221xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_586), .B1(n_590), .B2(n_593), .C(n_595), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
INVxp67_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g639 ( .A(n_583), .Y(n_639) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_583), .Y(n_767) );
INVx1_ASAP7_75t_L g730 ( .A(n_585), .Y(n_730) );
AND2x2_ASAP7_75t_SL g740 ( .A(n_585), .B(n_609), .Y(n_740) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_589), .B(n_617), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
OR2x2_ASAP7_75t_L g623 ( .A(n_591), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g701 ( .A(n_591), .Y(n_701) );
AND2x2_ASAP7_75t_L g636 ( .A(n_592), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g682 ( .A(n_594), .B(n_642), .Y(n_682) );
AND2x2_ASAP7_75t_L g759 ( .A(n_594), .B(n_757), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_600), .B1(n_607), .B2(n_608), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g618 ( .A(n_599), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx2_ASAP7_75t_L g624 ( .A(n_602), .Y(n_624) );
AND2x4_ASAP7_75t_L g648 ( .A(n_602), .B(n_649), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g678 ( .A1(n_602), .A2(n_679), .B(n_680), .Y(n_678) );
AND2x2_ASAP7_75t_L g705 ( .A(n_602), .B(n_663), .Y(n_705) );
INVx2_ASAP7_75t_L g627 ( .A(n_603), .Y(n_627) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_603), .Y(n_660) );
INVx1_ASAP7_75t_SL g684 ( .A(n_604), .Y(n_684) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g615 ( .A(n_606), .Y(n_615) );
AND2x4_ASAP7_75t_SL g709 ( .A(n_606), .B(n_627), .Y(n_709) );
AND2x2_ASAP7_75t_L g706 ( .A(n_609), .B(n_652), .Y(n_706) );
AND2x2_ASAP7_75t_L g732 ( .A(n_609), .B(n_718), .Y(n_732) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_610), .Y(n_654) );
INVx1_ASAP7_75t_L g674 ( .A(n_610), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_618), .B1(n_621), .B2(n_623), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_616), .B(n_627), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_616), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g755 ( .A(n_616), .Y(n_755) );
INVx2_ASAP7_75t_SL g680 ( .A(n_618), .Y(n_680) );
AND2x2_ASAP7_75t_L g692 ( .A(n_620), .B(n_652), .Y(n_692) );
INVx2_ASAP7_75t_L g698 ( .A(n_620), .Y(n_698) );
INVxp33_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_626), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g748 ( .A(n_626), .Y(n_748) );
INVx1_ASAP7_75t_L g676 ( .A(n_628), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_629), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g687 ( .A(n_631), .B(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_631), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_655), .C(n_658), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B1(n_640), .B2(n_644), .C(n_647), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g753 ( .A(n_638), .Y(n_753) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g722 ( .A(n_639), .B(n_688), .Y(n_722) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g653 ( .A(n_642), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g724 ( .A(n_644), .Y(n_724) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g721 ( .A(n_645), .Y(n_721) );
INVx1_ASAP7_75t_L g727 ( .A(n_646), .Y(n_727) );
OR2x2_ASAP7_75t_L g750 ( .A(n_646), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_SL g659 ( .A(n_649), .Y(n_659) );
AND2x2_ASAP7_75t_L g729 ( .A(n_649), .B(n_709), .Y(n_729) );
AND2x2_ASAP7_75t_SL g761 ( .A(n_649), .B(n_662), .Y(n_761) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g766 ( .A(n_652), .Y(n_766) );
INVx1_ASAP7_75t_L g716 ( .A(n_654), .Y(n_716) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B(n_661), .C(n_665), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_659), .B(n_709), .Y(n_733) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_662), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AND2x2_ASAP7_75t_L g670 ( .A(n_664), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g751 ( .A(n_664), .Y(n_751) );
NAND4xp75_ASAP7_75t_L g666 ( .A(n_667), .B(n_723), .C(n_739), .D(n_760), .Y(n_666) );
NOR3x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_685), .C(n_707), .Y(n_667) );
NAND4xp75_ASAP7_75t_L g668 ( .A(n_669), .B(n_675), .C(n_678), .D(n_681), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_670), .B(n_672), .Y(n_669) );
AND2x2_ASAP7_75t_L g720 ( .A(n_671), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g745 ( .A(n_672), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_SL g734 ( .A(n_677), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_693), .Y(n_685) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_689), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_699), .B(n_703), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI322xp33_ASAP7_75t_L g725 ( .A1(n_697), .A2(n_726), .A3(n_730), .B1(n_731), .B2(n_733), .C1(n_734), .C2(n_735), .Y(n_725) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_698), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_701), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_702), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_712), .C(n_714), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_719), .B1(n_720), .B2(n_722), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B(n_729), .Y(n_726) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_732), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g742 ( .A(n_737), .B(n_743), .Y(n_742) );
O2A1O1Ixp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_746), .C(n_749), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_742), .B(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI221xp5_ASAP7_75t_SL g749 ( .A1(n_750), .A2(n_752), .B1(n_754), .B2(n_756), .C(n_758), .Y(n_749) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx11_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
CKINVDCx6p67_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
BUFx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVxp67_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx8_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
endmodule