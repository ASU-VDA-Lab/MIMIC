module fake_jpeg_27517_n_294 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_38),
.B(n_32),
.C(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_23),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_31),
.B1(n_16),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_39),
.B1(n_40),
.B2(n_33),
.Y(n_72)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_77),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_36),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_80),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_31),
.B1(n_23),
.B2(n_16),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_69),
.B1(n_74),
.B2(n_27),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_56),
.B1(n_43),
.B2(n_25),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_31),
.B1(n_16),
.B2(n_29),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_86),
.B1(n_39),
.B2(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_29),
.B1(n_28),
.B2(n_21),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_40),
.C(n_36),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_20),
.C(n_37),
.Y(n_111)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_39),
.B1(n_33),
.B2(n_30),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_95),
.B1(n_106),
.B2(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_56),
.B1(n_43),
.B2(n_17),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_84),
.B1(n_62),
.B2(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_21),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_92),
.B(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_98),
.Y(n_132)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_112),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_21),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_30),
.B1(n_20),
.B2(n_51),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_66),
.B1(n_65),
.B2(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_28),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_17),
.B1(n_27),
.B2(n_24),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_22),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_70),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_30),
.B1(n_20),
.B2(n_22),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_34),
.C(n_35),
.Y(n_119)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

AO21x2_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_85),
.B(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_126),
.B1(n_109),
.B2(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_117),
.B(n_125),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_122),
.B1(n_129),
.B2(n_95),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_133),
.C(n_111),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_75),
.A3(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_75),
.B(n_66),
.C(n_19),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_131),
.B(n_35),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_19),
.B1(n_24),
.B2(n_30),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_135),
.Y(n_153)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_128),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_81),
.B(n_37),
.C(n_35),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_81),
.C(n_37),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_26),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_155),
.B1(n_157),
.B2(n_164),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_96),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_160),
.B(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_146),
.C(n_149),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_93),
.C(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_93),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_92),
.C(n_81),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_156),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_90),
.B1(n_101),
.B2(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_101),
.B1(n_99),
.B2(n_106),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_159),
.B1(n_121),
.B2(n_130),
.Y(n_180)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_109),
.B1(n_97),
.B2(n_26),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_112),
.B(n_35),
.C(n_50),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_115),
.B1(n_139),
.B2(n_123),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_50),
.B(n_26),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_166),
.B(n_131),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_115),
.A2(n_22),
.B(n_1),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_22),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_167),
.B(n_119),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_22),
.C(n_15),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_2),
.C(n_3),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_191),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_184),
.B(n_189),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_117),
.B1(n_135),
.B2(n_125),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_174),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_137),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_170),
.C(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_179),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_131),
.B1(n_126),
.B2(n_120),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_190),
.B1(n_148),
.B2(n_163),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_134),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_12),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_127),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_193),
.C(n_191),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_134),
.B(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_128),
.B1(n_15),
.B2(n_14),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_143),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_13),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_154),
.B1(n_148),
.B2(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_12),
.C(n_11),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_193),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_197),
.A2(n_206),
.B1(n_209),
.B2(n_188),
.Y(n_226)
);

NAND2x1p5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_165),
.Y(n_199)
);

XOR2x1_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_210),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_144),
.C(n_149),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_203),
.C(n_207),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_167),
.C(n_152),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_9),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_156),
.B1(n_150),
.B2(n_140),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_140),
.C(n_166),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_162),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_217),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_162),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_3),
.Y(n_212)
);

FAx1_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_189),
.CI(n_171),
.CON(n_221),
.SN(n_221)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_224),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_228),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_169),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_177),
.B1(n_190),
.B2(n_182),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_194),
.B1(n_182),
.B2(n_173),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_192),
.B1(n_11),
.B2(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_210),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_9),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_234),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_4),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_235),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_198),
.B1(n_199),
.B2(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_245),
.B1(n_221),
.B2(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_212),
.B1(n_200),
.B2(n_201),
.Y(n_245)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_212),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_205),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_205),
.C(n_195),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_223),
.C(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_251),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_220),
.C(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_224),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_256),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_221),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_255),
.A2(n_241),
.B(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_261),
.B1(n_241),
.B2(n_245),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_247),
.B(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_267),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_249),
.B1(n_243),
.B2(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_243),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_277),
.B1(n_279),
.B2(n_4),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_276),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_242),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_255),
.B1(n_257),
.B2(n_251),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_5),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_254),
.B1(n_5),
.B2(n_6),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_262),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_283),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_262),
.B(n_267),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_277),
.C(n_279),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_265),
.B(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_288),
.B(n_281),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_287),
.B(n_283),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_7),
.C(n_8),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_291),
.A2(n_7),
.B(n_8),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_7),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_8),
.B(n_292),
.Y(n_294)
);


endmodule