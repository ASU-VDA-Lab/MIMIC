module fake_aes_7459_n_1461 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1461);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1461;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1117;
wire n_1007;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1291;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1335;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1442;
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_183), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_93), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_143), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_118), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_298), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_241), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_242), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_50), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_6), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_259), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_156), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_263), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_22), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_240), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_178), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_102), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_194), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_64), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_227), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_155), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_39), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_179), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_145), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_330), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_246), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_80), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_232), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_86), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_37), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_223), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_73), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_147), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_182), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_214), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_276), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_312), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_0), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_180), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_317), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_34), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_50), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_206), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_248), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_104), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_85), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_141), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_22), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_150), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_74), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_260), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_77), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_288), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_153), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_323), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_230), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_117), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_262), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_31), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_13), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_255), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_200), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_207), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_188), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_43), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_327), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_104), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_51), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_134), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_258), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_161), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_116), .Y(n_412) );
INVxp33_ASAP7_75t_SL g413 ( .A(n_30), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_213), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_37), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_303), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_46), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_315), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_266), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_139), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_269), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_296), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_105), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_17), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_25), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_116), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_5), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_292), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_201), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_75), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_61), .Y(n_431) );
BUFx2_ASAP7_75t_SL g432 ( .A(n_203), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_226), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_282), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_316), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_208), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_101), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_307), .Y(n_438) );
INVxp33_ASAP7_75t_L g439 ( .A(n_294), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_61), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_314), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_299), .Y(n_442) );
BUFx10_ASAP7_75t_L g443 ( .A(n_270), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_215), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_278), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_52), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_159), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_12), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_285), .Y(n_449) );
CKINVDCx14_ASAP7_75t_R g450 ( .A(n_334), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_231), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_176), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_88), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_17), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_341), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_275), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_338), .B(n_123), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_186), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_273), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_162), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_233), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_157), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_319), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_181), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_277), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_297), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_244), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_52), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_217), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_89), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_142), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_211), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_144), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_98), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_225), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_170), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_117), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_283), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_247), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_151), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_138), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_295), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_106), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_306), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_311), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_331), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_66), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_189), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_11), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_221), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_219), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_27), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_102), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_46), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_71), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_129), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_91), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_148), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_53), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_174), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_89), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_320), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_106), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_264), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_75), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_228), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_229), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_202), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_41), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_304), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_51), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_290), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_80), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_329), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_69), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_308), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g517 ( .A(n_103), .B(n_133), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_128), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_101), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_318), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_325), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_83), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_172), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_163), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_279), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_83), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_191), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_272), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_152), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_251), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_345), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_345), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_461), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_499), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_461), .Y(n_535) );
BUFx3_ASAP7_75t_L g536 ( .A(n_364), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_443), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_419), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_492), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_419), .Y(n_540) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_347), .A2(n_135), .B(n_132), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_499), .Y(n_542) );
NOR2xp33_ASAP7_75t_SL g543 ( .A(n_411), .B(n_136), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_419), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_503), .Y(n_545) );
OR2x6_ASAP7_75t_L g546 ( .A(n_432), .B(n_0), .Y(n_546) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_419), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_503), .Y(n_548) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_347), .A2(n_140), .B(n_137), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_422), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_343), .B(n_1), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_360), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_526), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_422), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_439), .B(n_1), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_422), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_511), .B(n_2), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_526), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_413), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_422), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_379), .B(n_4), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_520), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_520), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_344), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_348), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_520), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_413), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_520), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_500), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_500), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_439), .B(n_7), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_351), .Y(n_574) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_544), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_537), .B(n_472), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_544), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_539), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_544), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_555), .A2(n_350), .B1(n_359), .B2(n_354), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_537), .B(n_527), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_533), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_571), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_571), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_537), .B(n_443), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_571), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_533), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_572), .Y(n_588) );
HAxp5_ASAP7_75t_SL g589 ( .A(n_559), .B(n_390), .CON(n_589), .SN(n_589) );
BUFx6f_ASAP7_75t_SL g590 ( .A(n_546), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_544), .Y(n_591) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_544), .Y(n_592) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_555), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_544), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_572), .Y(n_595) );
INVxp33_ASAP7_75t_L g596 ( .A(n_539), .Y(n_596) );
AND2x6_ASAP7_75t_L g597 ( .A(n_573), .B(n_533), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_566), .B(n_372), .Y(n_598) );
INVx4_ASAP7_75t_L g599 ( .A(n_546), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_566), .B(n_398), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_567), .B(n_401), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_572), .Y(n_602) );
BUFx10_ASAP7_75t_L g603 ( .A(n_567), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_574), .B(n_443), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_535), .B(n_362), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_547), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_573), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_574), .B(n_372), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_546), .A2(n_367), .B1(n_370), .B2(n_369), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_535), .Y(n_610) );
INVx6_ASAP7_75t_L g611 ( .A(n_536), .Y(n_611) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_547), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_562), .B(n_441), .Y(n_613) );
INVx4_ASAP7_75t_L g614 ( .A(n_546), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_535), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_536), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_557), .A2(n_382), .B1(n_388), .B2(n_386), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_593), .B(n_536), .Y(n_618) );
INVx4_ASAP7_75t_L g619 ( .A(n_603), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_610), .Y(n_620) );
NOR2x2_ASAP7_75t_L g621 ( .A(n_589), .B(n_552), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_603), .B(n_562), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_603), .B(n_563), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_611), .Y(n_624) );
NOR2xp67_ASAP7_75t_SL g625 ( .A(n_599), .B(n_342), .Y(n_625) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_596), .Y(n_626) );
AO22x1_ASAP7_75t_L g627 ( .A1(n_599), .A2(n_519), .B1(n_518), .B2(n_365), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_603), .B(n_563), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_578), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_599), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_599), .Y(n_631) );
AND2x6_ASAP7_75t_SL g632 ( .A(n_589), .B(n_561), .Y(n_632) );
NAND2xp33_ASAP7_75t_L g633 ( .A(n_597), .B(n_342), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_614), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_607), .B(n_551), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_607), .B(n_551), .Y(n_636) );
INVx5_ASAP7_75t_L g637 ( .A(n_597), .Y(n_637) );
NOR2x2_ASAP7_75t_L g638 ( .A(n_590), .B(n_390), .Y(n_638) );
BUFx12f_ASAP7_75t_L g639 ( .A(n_614), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_614), .B(n_543), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_598), .B(n_426), .Y(n_641) );
NOR2xp67_ASAP7_75t_L g642 ( .A(n_614), .B(n_559), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_610), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_597), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_597), .B(n_365), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_597), .B(n_371), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_590), .A2(n_543), .B1(n_450), .B2(n_392), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_597), .B(n_433), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_611), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_611), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_609), .B(n_433), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_604), .B(n_569), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_608), .B(n_521), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_576), .Y(n_654) );
BUFx3_ASAP7_75t_L g655 ( .A(n_597), .Y(n_655) );
BUFx3_ASAP7_75t_L g656 ( .A(n_597), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_616), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_600), .B(n_521), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_581), .B(n_524), .Y(n_659) );
NOR2xp33_ASAP7_75t_SL g660 ( .A(n_590), .B(n_360), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_585), .B(n_569), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_582), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_616), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_580), .B(n_524), .Y(n_664) );
AND2x6_ASAP7_75t_L g665 ( .A(n_590), .B(n_605), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_582), .Y(n_666) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_605), .B(n_397), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_601), .A2(n_541), .B(n_549), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_613), .B(n_452), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_605), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_605), .B(n_531), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_617), .B(n_529), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_583), .B(n_531), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_582), .B(n_366), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_582), .B(n_541), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_587), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_611), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_615), .A2(n_405), .B1(n_408), .B2(n_407), .Y(n_678) );
OAI22xp5_ASAP7_75t_SL g679 ( .A1(n_583), .A2(n_487), .B1(n_415), .B2(n_477), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_587), .A2(n_374), .B1(n_377), .B2(n_366), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_587), .A2(n_377), .B1(n_383), .B2(n_374), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_587), .B(n_358), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_615), .B(n_417), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_584), .A2(n_549), .B(n_502), .Y(n_684) );
INVx5_ASAP7_75t_L g685 ( .A(n_611), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_615), .B(n_463), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_584), .A2(n_423), .B1(n_431), .B2(n_424), .Y(n_687) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_586), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_586), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_588), .B(n_346), .Y(n_690) );
INVx5_ASAP7_75t_L g691 ( .A(n_575), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_588), .A2(n_448), .B1(n_454), .B2(n_437), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_595), .A2(n_418), .B1(n_420), .B2(n_383), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_595), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_602), .B(n_549), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_602), .A2(n_420), .B1(n_429), .B2(n_418), .Y(n_696) );
INVxp33_ASAP7_75t_SL g697 ( .A(n_577), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_577), .Y(n_698) );
BUFx3_ASAP7_75t_L g699 ( .A(n_575), .Y(n_699) );
INVx3_ASAP7_75t_L g700 ( .A(n_575), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_575), .B(n_391), .Y(n_701) );
INVx3_ASAP7_75t_L g702 ( .A(n_575), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_577), .B(n_532), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_579), .A2(n_429), .B1(n_451), .B2(n_445), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_579), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_575), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_579), .A2(n_470), .B1(n_474), .B2(n_468), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g708 ( .A(n_660), .Y(n_708) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_619), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_622), .A2(n_628), .B(n_623), .Y(n_710) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_619), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_629), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_704), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_654), .B(n_415), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_642), .A2(n_451), .B1(n_459), .B2(n_445), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_635), .B(n_518), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_636), .B(n_519), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_622), .A2(n_549), .B(n_353), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_626), .B(n_487), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_689), .Y(n_720) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_704), .Y(n_721) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_665), .Y(n_722) );
BUFx12f_ASAP7_75t_L g723 ( .A(n_639), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_620), .A2(n_494), .B(n_496), .C(n_495), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_623), .A2(n_355), .B(n_352), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_641), .A2(n_497), .B(n_522), .C(n_505), .Y(n_726) );
O2A1O1Ixp33_ASAP7_75t_L g727 ( .A1(n_664), .A2(n_453), .B(n_534), .C(n_532), .Y(n_727) );
AO21x2_ASAP7_75t_L g728 ( .A1(n_668), .A2(n_361), .B(n_356), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_657), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_628), .A2(n_368), .B(n_363), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_667), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_661), .B(n_459), .Y(n_732) );
O2A1O1Ixp33_ASAP7_75t_L g733 ( .A1(n_672), .A2(n_542), .B(n_545), .C(n_534), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_695), .A2(n_376), .B(n_375), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_637), .B(n_393), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_670), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_679), .B(n_378), .C(n_357), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_670), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_627), .B(n_381), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_695), .A2(n_384), .B(n_380), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_661), .B(n_385), .Y(n_741) );
CKINVDCx14_ASAP7_75t_R g742 ( .A(n_693), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_668), .B(n_430), .C(n_349), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_707), .B(n_430), .C(n_349), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_674), .B(n_399), .Y(n_745) );
O2A1O1Ixp33_ASAP7_75t_L g746 ( .A1(n_618), .A2(n_545), .B(n_548), .C(n_542), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_652), .A2(n_558), .B1(n_553), .B2(n_548), .C(n_412), .Y(n_747) );
INVx3_ASAP7_75t_L g748 ( .A(n_670), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_696), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_652), .B(n_400), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_680), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_658), .B(n_425), .Y(n_752) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_665), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_637), .B(n_396), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_631), .A2(n_440), .B1(n_446), .B2(n_427), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_658), .B(n_483), .Y(n_756) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_665), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_643), .A2(n_517), .B(n_457), .C(n_389), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_665), .Y(n_759) );
BUFx2_ASAP7_75t_L g760 ( .A(n_665), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_681), .Y(n_761) );
NOR2xp67_ASAP7_75t_L g762 ( .A(n_669), .B(n_8), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_647), .A2(n_509), .B1(n_513), .B2(n_501), .Y(n_763) );
OA22x2_ASAP7_75t_L g764 ( .A1(n_638), .A2(n_515), .B1(n_395), .B2(n_402), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_688), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_675), .A2(n_403), .B(n_394), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_659), .B(n_406), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_653), .B(n_373), .Y(n_768) );
BUFx2_ASAP7_75t_L g769 ( .A(n_663), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_640), .A2(n_410), .B(n_404), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_637), .B(n_409), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_694), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_655), .A2(n_430), .B1(n_493), .B2(n_349), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_683), .B(n_414), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g775 ( .A1(n_684), .A2(n_428), .B(n_416), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_634), .B(n_421), .Y(n_776) );
CKINVDCx8_ASAP7_75t_R g777 ( .A(n_632), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_656), .A2(n_430), .B1(n_493), .B2(n_349), .Y(n_778) );
NOR2xp33_ASAP7_75t_SL g779 ( .A(n_625), .B(n_434), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_683), .B(n_444), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_662), .Y(n_781) );
NOR3xp33_ASAP7_75t_SL g782 ( .A(n_651), .B(n_476), .C(n_467), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_645), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_644), .B(n_387), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_666), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_700), .A2(n_606), .B(n_594), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_645), .B(n_484), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_673), .A2(n_435), .B1(n_442), .B2(n_438), .Y(n_788) );
OAI21xp33_ASAP7_75t_L g789 ( .A1(n_646), .A2(n_507), .B(n_490), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_646), .A2(n_449), .B(n_447), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_682), .A2(n_456), .B(n_455), .Y(n_791) );
O2A1O1Ixp33_ASAP7_75t_L g792 ( .A1(n_671), .A2(n_460), .B(n_462), .C(n_458), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_687), .A2(n_493), .B1(n_464), .B2(n_469), .C(n_466), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_648), .B(n_512), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_676), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_663), .A2(n_493), .B1(n_465), .B2(n_473), .Y(n_796) );
OR2x6_ASAP7_75t_L g797 ( .A(n_630), .B(n_471), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_648), .B(n_516), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_692), .B(n_8), .Y(n_799) );
INVx3_ASAP7_75t_L g800 ( .A(n_630), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_682), .A2(n_475), .B(n_479), .C(n_478), .Y(n_801) );
INVx2_ASAP7_75t_SL g802 ( .A(n_686), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_633), .A2(n_481), .B(n_480), .Y(n_803) );
INVxp67_ASAP7_75t_L g804 ( .A(n_686), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_703), .Y(n_805) );
O2A1O1Ixp5_ASAP7_75t_L g806 ( .A1(n_701), .A2(n_502), .B(n_482), .C(n_486), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_678), .Y(n_807) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_685), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g809 ( .A(n_685), .B(n_530), .Y(n_809) );
NOR2xp33_ASAP7_75t_SL g810 ( .A(n_685), .B(n_364), .Y(n_810) );
A2O1A1Ixp33_ASAP7_75t_L g811 ( .A1(n_624), .A2(n_485), .B(n_491), .C(n_488), .Y(n_811) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_685), .Y(n_812) );
INVx3_ASAP7_75t_SL g813 ( .A(n_621), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_649), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_690), .A2(n_498), .B1(n_506), .B2(n_504), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_650), .A2(n_508), .B(n_514), .C(n_510), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_677), .B(n_697), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_691), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_L g819 ( .A1(n_698), .A2(n_523), .B(n_528), .C(n_525), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_705), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_691), .B(n_9), .Y(n_821) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_702), .B(n_436), .Y(n_822) );
CKINVDCx8_ASAP7_75t_R g823 ( .A(n_691), .Y(n_823) );
O2A1O1Ixp33_ASAP7_75t_L g824 ( .A1(n_706), .A2(n_540), .B(n_550), .C(n_538), .Y(n_824) );
BUFx2_ASAP7_75t_L g825 ( .A(n_691), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_702), .B(n_554), .C(n_547), .Y(n_826) );
INVxp67_ASAP7_75t_L g827 ( .A(n_699), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_654), .B(n_9), .Y(n_828) );
AND2x4_ASAP7_75t_L g829 ( .A(n_642), .B(n_10), .Y(n_829) );
NAND2xp33_ASAP7_75t_L g830 ( .A(n_665), .B(n_547), .Y(n_830) );
O2A1O1Ixp33_ASAP7_75t_L g831 ( .A1(n_654), .A2(n_540), .B(n_550), .C(n_538), .Y(n_831) );
OAI22xp5_ASAP7_75t_SL g832 ( .A1(n_679), .A2(n_12), .B1(n_10), .B2(n_11), .Y(n_832) );
OR2x2_ASAP7_75t_L g833 ( .A(n_629), .B(n_13), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_688), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_642), .A2(n_540), .B1(n_550), .B2(n_538), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_629), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_642), .A2(n_565), .B1(n_568), .B2(n_560), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_688), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_622), .A2(n_606), .B(n_594), .Y(n_839) );
BUFx8_ASAP7_75t_L g840 ( .A(n_674), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_629), .Y(n_841) );
NAND2x1_ASAP7_75t_L g842 ( .A(n_665), .B(n_560), .Y(n_842) );
NOR3xp33_ASAP7_75t_L g843 ( .A(n_704), .B(n_568), .C(n_565), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_629), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_714), .A2(n_568), .B1(n_565), .B2(n_554), .Y(n_845) );
OAI21xp5_ASAP7_75t_L g846 ( .A1(n_710), .A2(n_554), .B(n_547), .Y(n_846) );
BUFx12f_ASAP7_75t_L g847 ( .A(n_723), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_720), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_804), .B(n_14), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_732), .B(n_15), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_747), .B(n_15), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_836), .A2(n_556), .B1(n_564), .B2(n_554), .Y(n_852) );
AO31x2_ASAP7_75t_L g853 ( .A1(n_718), .A2(n_556), .A3(n_564), .B(n_554), .Y(n_853) );
OAI21x1_ASAP7_75t_L g854 ( .A1(n_786), .A2(n_556), .B(n_554), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_708), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_731), .B(n_16), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_725), .A2(n_564), .B(n_570), .C(n_556), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_749), .B(n_16), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_802), .B(n_18), .Y(n_859) );
OR2x6_ASAP7_75t_L g860 ( .A(n_729), .B(n_18), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_712), .B(n_19), .Y(n_861) );
O2A1O1Ixp33_ASAP7_75t_L g862 ( .A1(n_726), .A2(n_23), .B(n_20), .C(n_21), .Y(n_862) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_715), .A2(n_23), .B1(n_20), .B2(n_21), .Y(n_863) );
AO31x2_ASAP7_75t_L g864 ( .A1(n_758), .A2(n_564), .A3(n_570), .B(n_556), .Y(n_864) );
OAI21xp33_ASAP7_75t_L g865 ( .A1(n_752), .A2(n_570), .B(n_564), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_775), .A2(n_592), .B(n_591), .Y(n_866) );
BUFx2_ASAP7_75t_L g867 ( .A(n_841), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_751), .A2(n_26), .B1(n_24), .B2(n_25), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_772), .Y(n_869) );
O2A1O1Ixp33_ASAP7_75t_L g870 ( .A1(n_724), .A2(n_27), .B(n_24), .C(n_26), .Y(n_870) );
BUFx3_ASAP7_75t_L g871 ( .A(n_844), .Y(n_871) );
BUFx2_ASAP7_75t_SL g872 ( .A(n_823), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_730), .A2(n_570), .B(n_592), .C(n_591), .Y(n_873) );
OAI21xp5_ASAP7_75t_L g874 ( .A1(n_766), .A2(n_149), .B(n_146), .Y(n_874) );
AO31x2_ASAP7_75t_L g875 ( .A1(n_734), .A2(n_592), .A3(n_612), .B(n_591), .Y(n_875) );
AO32x2_ASAP7_75t_L g876 ( .A1(n_837), .A2(n_28), .A3(n_29), .B1(n_30), .B2(n_31), .Y(n_876) );
AO31x2_ASAP7_75t_L g877 ( .A1(n_740), .A2(n_837), .A3(n_801), .B(n_788), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_807), .B(n_28), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_839), .A2(n_592), .B(n_591), .Y(n_879) );
O2A1O1Ixp33_ASAP7_75t_L g880 ( .A1(n_721), .A2(n_33), .B(n_29), .C(n_32), .Y(n_880) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_722), .Y(n_881) );
O2A1O1Ixp33_ASAP7_75t_L g882 ( .A1(n_811), .A2(n_34), .B(n_32), .C(n_33), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_761), .B(n_35), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_799), .Y(n_884) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_790), .A2(n_612), .B(n_158), .Y(n_885) );
O2A1O1Ixp33_ASAP7_75t_L g886 ( .A1(n_816), .A2(n_38), .B(n_35), .C(n_36), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_719), .A2(n_612), .B1(n_39), .B2(n_36), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_750), .A2(n_612), .B1(n_41), .B2(n_38), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_805), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_833), .Y(n_890) );
O2A1O1Ixp33_ASAP7_75t_L g891 ( .A1(n_792), .A2(n_43), .B(n_40), .C(n_42), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_716), .B(n_40), .Y(n_892) );
OAI21x1_ASAP7_75t_L g893 ( .A1(n_743), .A2(n_160), .B(n_154), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_781), .Y(n_894) );
INVx2_ASAP7_75t_SL g895 ( .A(n_840), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_829), .Y(n_896) );
O2A1O1Ixp33_ASAP7_75t_L g897 ( .A1(n_733), .A2(n_45), .B(n_42), .C(n_44), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_829), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_840), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_785), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_737), .A2(n_48), .B1(n_45), .B2(n_47), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_741), .B(n_717), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_770), .A2(n_165), .B(n_164), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_797), .A2(n_49), .B1(n_47), .B2(n_48), .Y(n_904) );
INVx5_ASAP7_75t_L g905 ( .A(n_709), .Y(n_905) );
AOI21xp5_ASAP7_75t_L g906 ( .A1(n_787), .A2(n_167), .B(n_166), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_795), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_742), .B(n_53), .Y(n_908) );
OAI21x1_ASAP7_75t_L g909 ( .A1(n_842), .A2(n_169), .B(n_168), .Y(n_909) );
OAI211xp5_ASAP7_75t_L g910 ( .A1(n_777), .A2(n_54), .B(n_55), .C(n_56), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_835), .Y(n_911) );
OAI21x1_ASAP7_75t_L g912 ( .A1(n_822), .A2(n_173), .B(n_171), .Y(n_912) );
AO32x2_ASAP7_75t_L g913 ( .A1(n_788), .A2(n_54), .A3(n_55), .B1(n_56), .B2(n_57), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_820), .Y(n_914) );
OA21x2_ASAP7_75t_L g915 ( .A1(n_826), .A2(n_177), .B(n_175), .Y(n_915) );
AOI21xp33_ASAP7_75t_L g916 ( .A1(n_739), .A2(n_57), .B(n_58), .Y(n_916) );
AO31x2_ASAP7_75t_L g917 ( .A1(n_803), .A2(n_58), .A3(n_59), .B(n_60), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g918 ( .A1(n_794), .A2(n_185), .B(n_184), .Y(n_918) );
INVx2_ASAP7_75t_SL g919 ( .A(n_709), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_755), .B(n_59), .Y(n_920) );
AND2x4_ASAP7_75t_L g921 ( .A(n_711), .B(n_60), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_798), .A2(n_190), .B(n_187), .Y(n_922) );
BUFx8_ASAP7_75t_SL g923 ( .A(n_769), .Y(n_923) );
BUFx2_ASAP7_75t_L g924 ( .A(n_797), .Y(n_924) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_745), .A2(n_62), .B1(n_63), .B2(n_64), .C(n_65), .Y(n_925) );
O2A1O1Ixp33_ASAP7_75t_SL g926 ( .A1(n_735), .A2(n_235), .B(n_340), .C(n_339), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_828), .B(n_62), .Y(n_927) );
BUFx8_ASAP7_75t_SL g928 ( .A(n_783), .Y(n_928) );
O2A1O1Ixp33_ASAP7_75t_SL g929 ( .A1(n_754), .A2(n_234), .B(n_337), .C(n_336), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_764), .A2(n_63), .B1(n_65), .B2(n_66), .Y(n_930) );
O2A1O1Ixp33_ASAP7_75t_SL g931 ( .A1(n_771), .A2(n_236), .B(n_335), .C(n_333), .Y(n_931) );
NOR2xp67_ASAP7_75t_L g932 ( .A(n_768), .B(n_67), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_797), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_736), .Y(n_934) );
AOI32xp33_ASAP7_75t_L g935 ( .A1(n_763), .A2(n_67), .A3(n_68), .B1(n_69), .B2(n_70), .Y(n_935) );
OAI21x1_ASAP7_75t_L g936 ( .A1(n_765), .A2(n_193), .B(n_192), .Y(n_936) );
O2A1O1Ixp5_ASAP7_75t_L g937 ( .A1(n_791), .A2(n_238), .B(n_332), .C(n_328), .Y(n_937) );
A2O1A1Ixp33_ASAP7_75t_L g938 ( .A1(n_727), .A2(n_71), .B(n_72), .C(n_73), .Y(n_938) );
O2A1O1Ixp33_ASAP7_75t_SL g939 ( .A1(n_809), .A2(n_746), .B(n_827), .C(n_791), .Y(n_939) );
OAI22x1_ASAP7_75t_L g940 ( .A1(n_813), .A2(n_72), .B1(n_74), .B2(n_76), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_756), .B(n_76), .Y(n_941) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_728), .A2(n_196), .B(n_195), .Y(n_942) );
AOI21xp5_ASAP7_75t_L g943 ( .A1(n_728), .A2(n_198), .B(n_197), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_832), .A2(n_77), .B1(n_78), .B2(n_79), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_843), .A2(n_78), .B1(n_79), .B2(n_81), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_711), .B(n_81), .Y(n_946) );
A2O1A1Ixp33_ASAP7_75t_L g947 ( .A1(n_819), .A2(n_82), .B(n_84), .C(n_85), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_767), .A2(n_204), .B(n_199), .Y(n_948) );
A2O1A1Ixp33_ASAP7_75t_L g949 ( .A1(n_762), .A2(n_82), .B(n_84), .C(n_86), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_722), .A2(n_757), .B1(n_753), .B2(n_760), .Y(n_950) );
OAI21xp5_ASAP7_75t_L g951 ( .A1(n_806), .A2(n_209), .B(n_205), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_774), .B(n_87), .Y(n_952) );
AOI21xp5_ASAP7_75t_L g953 ( .A1(n_834), .A2(n_254), .B(n_326), .Y(n_953) );
O2A1O1Ixp33_ASAP7_75t_L g954 ( .A1(n_831), .A2(n_87), .B(n_88), .C(n_90), .Y(n_954) );
AO31x2_ASAP7_75t_L g955 ( .A1(n_778), .A2(n_814), .A3(n_838), .B(n_738), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_817), .Y(n_956) );
BUFx3_ASAP7_75t_L g957 ( .A(n_711), .Y(n_957) );
AND2x4_ASAP7_75t_L g958 ( .A(n_753), .B(n_90), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_780), .B(n_91), .Y(n_959) );
BUFx6f_ASAP7_75t_L g960 ( .A(n_753), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_789), .A2(n_256), .B(n_324), .Y(n_961) );
O2A1O1Ixp33_ASAP7_75t_L g962 ( .A1(n_793), .A2(n_92), .B(n_93), .C(n_94), .Y(n_962) );
OR2x2_ASAP7_75t_L g963 ( .A(n_815), .B(n_92), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_748), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_964) );
AO31x2_ASAP7_75t_L g965 ( .A1(n_784), .A2(n_95), .A3(n_97), .B(n_98), .Y(n_965) );
BUFx3_ASAP7_75t_L g966 ( .A(n_825), .Y(n_966) );
NAND2xp5_ASAP7_75t_SL g967 ( .A(n_757), .B(n_97), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_759), .A2(n_99), .B1(n_100), .B2(n_103), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_757), .A2(n_99), .B1(n_100), .B2(n_105), .Y(n_969) );
AOI21xp5_ASAP7_75t_L g970 ( .A1(n_830), .A2(n_261), .B(n_322), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_782), .B(n_107), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_800), .A2(n_107), .B1(n_108), .B2(n_109), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_800), .A2(n_108), .B1(n_109), .B2(n_110), .Y(n_973) );
AOI21xp5_ASAP7_75t_L g974 ( .A1(n_776), .A2(n_265), .B(n_321), .Y(n_974) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_818), .Y(n_975) );
AOI221x1_ASAP7_75t_L g976 ( .A1(n_744), .A2(n_110), .B1(n_111), .B2(n_112), .C(n_113), .Y(n_976) );
BUFx6f_ASAP7_75t_L g977 ( .A(n_808), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_821), .Y(n_978) );
CKINVDCx11_ASAP7_75t_R g979 ( .A(n_808), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_796), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g981 ( .A1(n_779), .A2(n_257), .B(n_313), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_779), .A2(n_111), .B1(n_112), .B2(n_113), .Y(n_982) );
OAI21x1_ASAP7_75t_L g983 ( .A1(n_824), .A2(n_267), .B(n_310), .Y(n_983) );
OAI22x1_ASAP7_75t_L g984 ( .A1(n_810), .A2(n_114), .B1(n_115), .B2(n_118), .Y(n_984) );
AOI21xp5_ASAP7_75t_L g985 ( .A1(n_810), .A2(n_268), .B(n_309), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_812), .B(n_114), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g987 ( .A(n_773), .B(n_119), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_836), .B(n_119), .Y(n_988) );
A2O1A1Ixp33_ASAP7_75t_L g989 ( .A1(n_710), .A2(n_120), .B(n_121), .C(n_122), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g990 ( .A(n_732), .B(n_120), .Y(n_990) );
NAND2xp5_ASAP7_75t_SL g991 ( .A(n_709), .B(n_121), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_772), .Y(n_992) );
A2O1A1Ixp33_ASAP7_75t_L g993 ( .A1(n_710), .A2(n_122), .B(n_123), .C(n_124), .Y(n_993) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_836), .Y(n_994) );
INVx5_ASAP7_75t_L g995 ( .A(n_709), .Y(n_995) );
AOI221xp5_ASAP7_75t_SL g996 ( .A1(n_726), .A2(n_124), .B1(n_125), .B2(n_126), .C(n_127), .Y(n_996) );
A2O1A1Ixp33_ASAP7_75t_L g997 ( .A1(n_710), .A2(n_125), .B(n_126), .C(n_127), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_720), .Y(n_998) );
INVxp67_ASAP7_75t_L g999 ( .A(n_836), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_836), .B(n_128), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_884), .B(n_129), .Y(n_1001) );
OAI21xp5_ASAP7_75t_L g1002 ( .A1(n_846), .A2(n_130), .B(n_131), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_889), .B(n_130), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_956), .B(n_131), .Y(n_1004) );
AO31x2_ASAP7_75t_L g1005 ( .A1(n_866), .A2(n_210), .A3(n_212), .B(n_216), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_848), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_867), .B(n_218), .Y(n_1007) );
O2A1O1Ixp33_ASAP7_75t_L g1008 ( .A1(n_850), .A2(n_220), .B(n_222), .C(n_224), .Y(n_1008) );
NAND2x1p5_ASAP7_75t_L g1009 ( .A(n_905), .B(n_305), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_994), .B(n_237), .Y(n_1010) );
AND2x4_ASAP7_75t_L g1011 ( .A(n_924), .B(n_239), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_914), .Y(n_1012) );
A2O1A1Ixp33_ASAP7_75t_L g1013 ( .A1(n_891), .A2(n_243), .B(n_245), .C(n_249), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_914), .Y(n_1014) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_871), .Y(n_1015) );
AOI21xp5_ASAP7_75t_L g1016 ( .A1(n_939), .A2(n_250), .B(n_252), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_999), .B(n_253), .Y(n_1017) );
INVx4_ASAP7_75t_SL g1018 ( .A(n_847), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_894), .Y(n_1019) );
AOI222xp33_ASAP7_75t_L g1020 ( .A1(n_908), .A2(n_271), .B1(n_274), .B2(n_280), .C1(n_281), .C2(n_284), .Y(n_1020) );
OAI21xp5_ASAP7_75t_L g1021 ( .A1(n_851), .A2(n_286), .B(n_287), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_873), .A2(n_289), .B(n_291), .Y(n_1022) );
BUFx12f_ASAP7_75t_L g1023 ( .A(n_895), .Y(n_1023) );
AOI222xp33_ASAP7_75t_L g1024 ( .A1(n_858), .A2(n_883), .B1(n_940), .B2(n_920), .C1(n_890), .C2(n_944), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_905), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_998), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_988), .B(n_293), .Y(n_1027) );
INVx2_ASAP7_75t_L g1028 ( .A(n_900), .Y(n_1028) );
NOR2xp67_ASAP7_75t_L g1029 ( .A(n_995), .B(n_302), .Y(n_1029) );
OA21x2_ASAP7_75t_L g1030 ( .A1(n_893), .A2(n_300), .B(n_301), .Y(n_1030) );
AND2x4_ASAP7_75t_L g1031 ( .A(n_995), .B(n_933), .Y(n_1031) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_897), .A2(n_862), .B(n_880), .C(n_962), .Y(n_1032) );
BUFx3_ASAP7_75t_L g1033 ( .A(n_979), .Y(n_1033) );
AOI211xp5_ASAP7_75t_L g1034 ( .A1(n_868), .A2(n_863), .B(n_904), .C(n_910), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_860), .A2(n_896), .B1(n_898), .B2(n_899), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_892), .B(n_952), .Y(n_1036) );
O2A1O1Ixp33_ASAP7_75t_SL g1037 ( .A1(n_989), .A2(n_993), .B(n_997), .C(n_938), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_907), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_869), .Y(n_1039) );
AOI222xp33_ASAP7_75t_L g1040 ( .A1(n_925), .A2(n_930), .B1(n_855), .B2(n_901), .C1(n_984), .C2(n_975), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_860), .B(n_1000), .Y(n_1041) );
INVxp33_ASAP7_75t_L g1042 ( .A(n_928), .Y(n_1042) );
A2O1A1Ixp33_ASAP7_75t_L g1043 ( .A1(n_954), .A2(n_870), .B(n_932), .C(n_882), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_963), .B(n_849), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_861), .B(n_966), .Y(n_1045) );
O2A1O1Ixp33_ASAP7_75t_L g1046 ( .A1(n_947), .A2(n_949), .B(n_927), .C(n_959), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_992), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_859), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_934), .Y(n_1049) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_923), .Y(n_1050) );
AOI21xp5_ASAP7_75t_L g1051 ( .A1(n_885), .A2(n_865), .B(n_942), .Y(n_1051) );
OA21x2_ASAP7_75t_L g1052 ( .A1(n_943), .A2(n_937), .B(n_936), .Y(n_1052) );
INVx4_ASAP7_75t_L g1053 ( .A(n_995), .Y(n_1053) );
INVx3_ASAP7_75t_L g1054 ( .A(n_957), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_921), .A2(n_887), .B1(n_878), .B2(n_986), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_877), .B(n_978), .Y(n_1056) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_856), .B(n_872), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_977), .Y(n_1058) );
OA21x2_ASAP7_75t_L g1059 ( .A1(n_912), .A2(n_983), .B(n_857), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_921), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_877), .B(n_911), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_877), .B(n_996), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_845), .B(n_935), .Y(n_1063) );
OA21x2_ASAP7_75t_L g1064 ( .A1(n_874), .A2(n_976), .B(n_951), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_986), .A2(n_888), .B1(n_958), .B2(n_945), .Y(n_1065) );
OAI21xp5_ASAP7_75t_L g1066 ( .A1(n_906), .A2(n_918), .B(n_922), .Y(n_1066) );
OAI21x1_ASAP7_75t_L g1067 ( .A1(n_909), .A2(n_948), .B(n_970), .Y(n_1067) );
AO31x2_ASAP7_75t_L g1068 ( .A1(n_961), .A2(n_985), .A3(n_981), .B(n_953), .Y(n_1068) );
A2O1A1Ixp33_ASAP7_75t_L g1069 ( .A1(n_886), .A2(n_987), .B(n_982), .C(n_916), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_965), .Y(n_1070) );
A2O1A1Ixp33_ASAP7_75t_L g1071 ( .A1(n_971), .A2(n_980), .B(n_974), .C(n_946), .Y(n_1071) );
INVx3_ASAP7_75t_SL g1072 ( .A(n_919), .Y(n_1072) );
OAI21xp5_ASAP7_75t_L g1073 ( .A1(n_903), .A2(n_967), .B(n_852), .Y(n_1073) );
OAI21xp5_ASAP7_75t_L g1074 ( .A1(n_968), .A2(n_991), .B(n_973), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_977), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_917), .Y(n_1076) );
BUFx4f_ASAP7_75t_L g1077 ( .A(n_958), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_917), .Y(n_1078) );
BUFx6f_ASAP7_75t_L g1079 ( .A(n_960), .Y(n_1079) );
OAI21xp5_ASAP7_75t_SL g1080 ( .A1(n_972), .A2(n_964), .B(n_969), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_917), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_913), .Y(n_1082) );
AOI21xp5_ASAP7_75t_L g1083 ( .A1(n_926), .A2(n_931), .B(n_929), .Y(n_1083) );
OA21x2_ASAP7_75t_L g1084 ( .A1(n_853), .A2(n_864), .B(n_875), .Y(n_1084) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_960), .B(n_881), .Y(n_1085) );
INVx3_ASAP7_75t_L g1086 ( .A(n_960), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_864), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_950), .A2(n_913), .B1(n_876), .B2(n_915), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_913), .A2(n_876), .B1(n_955), .B2(n_875), .Y(n_1089) );
BUFx6f_ASAP7_75t_L g1090 ( .A(n_876), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_955), .B(n_629), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_955), .Y(n_1092) );
CKINVDCx6p67_ASAP7_75t_R g1093 ( .A(n_847), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_889), .B(n_731), .Y(n_1094) );
OA21x2_ASAP7_75t_L g1095 ( .A1(n_846), .A2(n_743), .B(n_854), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_867), .B(n_629), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_850), .A2(n_732), .B1(n_742), .B2(n_737), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_848), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_884), .B(n_593), .Y(n_1099) );
BUFx6f_ASAP7_75t_L g1100 ( .A(n_905), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_889), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_848), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_871), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_848), .Y(n_1104) );
CKINVDCx11_ASAP7_75t_R g1105 ( .A(n_847), .Y(n_1105) );
INVxp67_ASAP7_75t_L g1106 ( .A(n_867), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1107 ( .A(n_867), .B(n_629), .Y(n_1107) );
A2O1A1Ixp33_ASAP7_75t_L g1108 ( .A1(n_941), .A2(n_850), .B(n_990), .C(n_891), .Y(n_1108) );
AOI21xp5_ASAP7_75t_L g1109 ( .A1(n_846), .A2(n_879), .B(n_866), .Y(n_1109) );
AO21x2_ASAP7_75t_L g1110 ( .A1(n_846), .A2(n_743), .B(n_866), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_884), .B(n_593), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_884), .A2(n_721), .B1(n_713), .B2(n_921), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_850), .A2(n_732), .B1(n_742), .B2(n_737), .Y(n_1113) );
AOI21xp5_ASAP7_75t_L g1114 ( .A1(n_846), .A2(n_879), .B(n_866), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_889), .Y(n_1115) );
AO31x2_ASAP7_75t_L g1116 ( .A1(n_866), .A2(n_943), .A3(n_942), .B(n_873), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_884), .B(n_593), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_884), .B(n_593), .Y(n_1118) );
OR2x6_ASAP7_75t_L g1119 ( .A(n_872), .B(n_704), .Y(n_1119) );
AOI21xp33_ASAP7_75t_L g1120 ( .A1(n_902), .A2(n_727), .B(n_941), .Y(n_1120) );
A2O1A1Ixp33_ASAP7_75t_L g1121 ( .A1(n_941), .A2(n_850), .B(n_990), .C(n_891), .Y(n_1121) );
AOI21xp5_ASAP7_75t_L g1122 ( .A1(n_846), .A2(n_879), .B(n_866), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_889), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_850), .A2(n_732), .B1(n_742), .B2(n_737), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_956), .B(n_654), .Y(n_1125) );
OA21x2_ASAP7_75t_L g1126 ( .A1(n_846), .A2(n_743), .B(n_854), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_848), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_848), .Y(n_1128) );
A2O1A1Ixp33_ASAP7_75t_L g1129 ( .A1(n_941), .A2(n_850), .B(n_990), .C(n_891), .Y(n_1129) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_902), .A2(n_704), .B1(n_732), .B2(n_674), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_889), .Y(n_1131) );
AND2x4_ASAP7_75t_L g1132 ( .A(n_889), .B(n_731), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g1133 ( .A1(n_860), .A2(n_704), .B1(n_696), .B2(n_693), .Y(n_1133) );
OA21x2_ASAP7_75t_L g1134 ( .A1(n_846), .A2(n_743), .B(n_854), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_884), .A2(n_721), .B1(n_713), .B2(n_921), .Y(n_1135) );
AO21x2_ASAP7_75t_L g1136 ( .A1(n_846), .A2(n_743), .B(n_866), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_889), .Y(n_1137) );
BUFx2_ASAP7_75t_L g1138 ( .A(n_871), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_867), .B(n_629), .Y(n_1139) );
NOR2xp33_ASAP7_75t_L g1140 ( .A(n_902), .B(n_742), .Y(n_1140) );
A2O1A1Ixp33_ASAP7_75t_L g1141 ( .A1(n_941), .A2(n_850), .B(n_990), .C(n_891), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1012), .B(n_1014), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1024), .A2(n_1040), .B1(n_1133), .B2(n_1120), .Y(n_1143) );
BUFx4f_ASAP7_75t_SL g1144 ( .A(n_1093), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1006), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1019), .B(n_1028), .Y(n_1146) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1084), .Y(n_1147) );
INVx3_ASAP7_75t_L g1148 ( .A(n_1100), .Y(n_1148) );
OAI21xp5_ASAP7_75t_L g1149 ( .A1(n_1108), .A2(n_1129), .B(n_1121), .Y(n_1149) );
AOI22xp5_ASAP7_75t_L g1150 ( .A1(n_1140), .A2(n_1024), .B1(n_1125), .B2(n_1130), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_1097), .A2(n_1124), .B1(n_1113), .B2(n_1130), .C(n_1141), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1026), .B(n_1098), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_1040), .A2(n_1119), .B1(n_1044), .B2(n_1135), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_1119), .A2(n_1135), .B1(n_1112), .B2(n_1063), .Y(n_1154) );
OAI222xp33_ASAP7_75t_L g1155 ( .A1(n_1119), .A2(n_1112), .B1(n_1011), .B2(n_1065), .C1(n_1055), .C2(n_1091), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1092), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1096), .B(n_1107), .Y(n_1157) );
INVxp67_ASAP7_75t_L g1158 ( .A(n_1139), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1015), .B(n_1138), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1102), .B(n_1104), .Y(n_1160) );
AOI21xp5_ASAP7_75t_SL g1161 ( .A1(n_1011), .A2(n_1002), .B(n_1055), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1162 ( .A(n_1036), .B(n_1041), .Y(n_1162) );
OAI21xp5_ASAP7_75t_L g1163 ( .A1(n_1032), .A2(n_1043), .B(n_1069), .Y(n_1163) );
OA21x2_ASAP7_75t_L g1164 ( .A1(n_1062), .A2(n_1089), .B(n_1078), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g1165 ( .A1(n_1099), .A2(n_1111), .B1(n_1117), .B2(n_1118), .C(n_1035), .Y(n_1165) );
OA21x2_ASAP7_75t_L g1166 ( .A1(n_1076), .A2(n_1081), .B(n_1070), .Y(n_1166) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1086), .B(n_1058), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1038), .B(n_1039), .Y(n_1168) );
OR2x6_ASAP7_75t_L g1169 ( .A(n_1065), .B(n_1009), .Y(n_1169) );
AO31x2_ASAP7_75t_L g1170 ( .A1(n_1088), .A2(n_1061), .A3(n_1056), .B(n_1082), .Y(n_1170) );
OAI21xp5_ASAP7_75t_L g1171 ( .A1(n_1046), .A2(n_1080), .B(n_1074), .Y(n_1171) );
AO21x2_ASAP7_75t_L g1172 ( .A1(n_1088), .A2(n_1051), .B(n_1136), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1127), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1047), .B(n_1101), .Y(n_1174) );
OA21x2_ASAP7_75t_L g1175 ( .A1(n_1087), .A2(n_1071), .B(n_1016), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_1106), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1128), .Y(n_1177) );
AO21x2_ASAP7_75t_L g1178 ( .A1(n_1110), .A2(n_1136), .B(n_1002), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1115), .B(n_1123), .Y(n_1179) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_1100), .Y(n_1180) );
OAI21xp5_ASAP7_75t_L g1181 ( .A1(n_1080), .A2(n_1074), .B(n_1034), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1131), .B(n_1137), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1049), .Y(n_1183) );
OR2x6_ASAP7_75t_L g1184 ( .A(n_1053), .B(n_1100), .Y(n_1184) );
OAI211xp5_ASAP7_75t_L g1185 ( .A1(n_1034), .A2(n_1020), .B(n_1057), .C(n_1001), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_1048), .A2(n_1090), .B1(n_1020), .B2(n_1077), .Y(n_1186) );
BUFx3_ASAP7_75t_L g1187 ( .A(n_1072), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1094), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1094), .Y(n_1189) );
INVx3_ASAP7_75t_L g1190 ( .A(n_1053), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1132), .Y(n_1191) );
OAI21x1_ASAP7_75t_L g1192 ( .A1(n_1067), .A2(n_1083), .B(n_1126), .Y(n_1192) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1045), .B(n_1010), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1004), .B(n_1003), .Y(n_1194) );
OAI21x1_ASAP7_75t_L g1195 ( .A1(n_1095), .A2(n_1134), .B(n_1126), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1060), .B(n_1027), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_1105), .Y(n_1197) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_1025), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1017), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1007), .Y(n_1200) );
AOI22xp33_ASAP7_75t_SL g1201 ( .A1(n_1033), .A2(n_1090), .B1(n_1021), .B2(n_1050), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1031), .B(n_1054), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_1031), .Y(n_1203) );
AO21x2_ASAP7_75t_L g1204 ( .A1(n_1110), .A2(n_1073), .B(n_1066), .Y(n_1204) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1079), .Y(n_1205) );
INVx3_ASAP7_75t_L g1206 ( .A(n_1079), .Y(n_1206) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1086), .Y(n_1207) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1005), .Y(n_1208) );
BUFx3_ASAP7_75t_L g1209 ( .A(n_1023), .Y(n_1209) );
INVx4_ASAP7_75t_L g1210 ( .A(n_1054), .Y(n_1210) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1005), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1090), .Y(n_1212) );
OAI21xp5_ASAP7_75t_L g1213 ( .A1(n_1013), .A2(n_1073), .B(n_1037), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1214 ( .A(n_1075), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1085), .B(n_1021), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1029), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1029), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1042), .B(n_1085), .Y(n_1218) );
INVx2_ASAP7_75t_SL g1219 ( .A(n_1018), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1064), .B(n_1116), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1008), .Y(n_1221) );
BUFx3_ASAP7_75t_L g1222 ( .A(n_1059), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1116), .B(n_1030), .Y(n_1223) );
INVx4_ASAP7_75t_L g1224 ( .A(n_1052), .Y(n_1224) );
AND2x4_ASAP7_75t_L g1225 ( .A(n_1022), .B(n_1068), .Y(n_1225) );
HB1xp67_ASAP7_75t_L g1226 ( .A(n_1068), .Y(n_1226) );
OR2x6_ASAP7_75t_L g1227 ( .A(n_1011), .B(n_1112), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1096), .B(n_1107), .Y(n_1228) );
AO21x2_ASAP7_75t_L g1229 ( .A1(n_1109), .A2(n_1122), .B(n_1114), .Y(n_1229) );
INVx5_ASAP7_75t_SL g1230 ( .A(n_1093), .Y(n_1230) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1012), .Y(n_1231) );
HB1xp67_ASAP7_75t_L g1232 ( .A(n_1103), .Y(n_1232) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1012), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1012), .B(n_1014), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1235 ( .A(n_1103), .Y(n_1235) );
INVx1_ASAP7_75t_SL g1236 ( .A(n_1015), .Y(n_1236) );
OAI21xp5_ASAP7_75t_L g1237 ( .A1(n_1108), .A2(n_1129), .B(n_1121), .Y(n_1237) );
HB1xp67_ASAP7_75t_L g1238 ( .A(n_1103), .Y(n_1238) );
INVx2_ASAP7_75t_SL g1239 ( .A(n_1100), .Y(n_1239) );
NOR2xp33_ASAP7_75t_L g1240 ( .A(n_1133), .B(n_749), .Y(n_1240) );
BUFx3_ASAP7_75t_L g1241 ( .A(n_1100), .Y(n_1241) );
INVx2_ASAP7_75t_SL g1242 ( .A(n_1100), .Y(n_1242) );
OA21x2_ASAP7_75t_L g1243 ( .A1(n_1109), .A2(n_1122), .B(n_1114), .Y(n_1243) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1012), .Y(n_1244) );
AND2x4_ASAP7_75t_L g1245 ( .A(n_1169), .B(n_1147), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_1143), .A2(n_1151), .B1(n_1181), .B2(n_1240), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1166), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1227), .B(n_1171), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1143), .B(n_1179), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1142), .B(n_1234), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1231), .B(n_1244), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1227), .B(n_1231), .Y(n_1252) );
INVx3_ASAP7_75t_L g1253 ( .A(n_1169), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1182), .B(n_1150), .Y(n_1254) );
INVx3_ASAP7_75t_L g1255 ( .A(n_1169), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1233), .B(n_1244), .Y(n_1256) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_1233), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1227), .B(n_1157), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1174), .B(n_1168), .Y(n_1259) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_1232), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_1240), .A2(n_1153), .B1(n_1227), .B2(n_1186), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1174), .B(n_1168), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_1153), .A2(n_1186), .B1(n_1154), .B2(n_1237), .Y(n_1263) );
NOR2xp67_ASAP7_75t_L g1264 ( .A(n_1210), .B(n_1190), .Y(n_1264) );
HB1xp67_ASAP7_75t_L g1265 ( .A(n_1235), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1146), .B(n_1163), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1146), .B(n_1220), .Y(n_1267) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_1238), .Y(n_1268) );
INVx3_ASAP7_75t_L g1269 ( .A(n_1169), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1228), .B(n_1154), .Y(n_1270) );
INVxp67_ASAP7_75t_SL g1271 ( .A(n_1196), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1220), .B(n_1164), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1158), .B(n_1145), .Y(n_1273) );
NOR2xp67_ASAP7_75t_L g1274 ( .A(n_1210), .B(n_1190), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1166), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1164), .B(n_1156), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1149), .B(n_1183), .Y(n_1277) );
AND2x4_ASAP7_75t_L g1278 ( .A(n_1212), .B(n_1216), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1173), .B(n_1177), .Y(n_1279) );
BUFx2_ASAP7_75t_L g1280 ( .A(n_1210), .Y(n_1280) );
OAI21xp5_ASAP7_75t_L g1281 ( .A1(n_1185), .A2(n_1155), .B(n_1194), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1166), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1170), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1170), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1170), .B(n_1159), .Y(n_1285) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1170), .B(n_1193), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1162), .B(n_1152), .Y(n_1287) );
HB1xp67_ASAP7_75t_L g1288 ( .A(n_1198), .Y(n_1288) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_1162), .A2(n_1165), .B1(n_1196), .B2(n_1199), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1226), .Y(n_1290) );
AND2x4_ASAP7_75t_L g1291 ( .A(n_1217), .B(n_1205), .Y(n_1291) );
INVx1_ASAP7_75t_SL g1292 ( .A(n_1187), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1236), .B(n_1160), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1176), .B(n_1200), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1204), .B(n_1178), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1229), .Y(n_1296) );
HB1xp67_ASAP7_75t_L g1297 ( .A(n_1180), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1218), .B(n_1161), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1229), .Y(n_1299) );
OR2x6_ASAP7_75t_SL g1300 ( .A(n_1197), .B(n_1161), .Y(n_1300) );
BUFx3_ASAP7_75t_L g1301 ( .A(n_1241), .Y(n_1301) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1203), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1214), .B(n_1184), .Y(n_1303) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1184), .B(n_1215), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1184), .B(n_1202), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1172), .B(n_1243), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1286), .B(n_1201), .Y(n_1307) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1286), .B(n_1208), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1285), .B(n_1211), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1267), .B(n_1223), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1267), .B(n_1223), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1272), .B(n_1211), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1272), .B(n_1222), .Y(n_1313) );
NAND3xp33_ASAP7_75t_L g1314 ( .A(n_1246), .B(n_1221), .C(n_1213), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1249), .B(n_1225), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_1257), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1247), .Y(n_1317) );
INVx2_ASAP7_75t_SL g1318 ( .A(n_1280), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1250), .B(n_1195), .Y(n_1319) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_1280), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1295), .B(n_1195), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1250), .B(n_1225), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1285), .B(n_1225), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1259), .B(n_1224), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1275), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1295), .B(n_1224), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1270), .B(n_1191), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1282), .Y(n_1328) );
INVx1_ASAP7_75t_SL g1329 ( .A(n_1301), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1259), .B(n_1224), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1270), .B(n_1188), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1251), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1251), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1256), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1277), .B(n_1189), .Y(n_1335) );
INVx2_ASAP7_75t_SL g1336 ( .A(n_1303), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1306), .B(n_1192), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1256), .Y(n_1338) );
BUFx2_ASAP7_75t_L g1339 ( .A(n_1300), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1262), .B(n_1175), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1262), .B(n_1175), .Y(n_1341) );
BUFx3_ASAP7_75t_L g1342 ( .A(n_1301), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1289), .B(n_1167), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1319), .B(n_1276), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1332), .B(n_1279), .Y(n_1345) );
INVx1_ASAP7_75t_SL g1346 ( .A(n_1329), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1317), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1319), .B(n_1276), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1315), .B(n_1258), .Y(n_1349) );
NAND2xp33_ASAP7_75t_SL g1350 ( .A(n_1339), .B(n_1219), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1340), .B(n_1283), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1341), .B(n_1284), .Y(n_1352) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_1315), .B(n_1258), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1317), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1310), .B(n_1248), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1332), .B(n_1279), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1333), .B(n_1248), .Y(n_1357) );
INVx1_ASAP7_75t_SL g1358 ( .A(n_1329), .Y(n_1358) );
INVx2_ASAP7_75t_L g1359 ( .A(n_1325), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1333), .B(n_1260), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1334), .B(n_1265), .Y(n_1361) );
HB1xp67_ASAP7_75t_L g1362 ( .A(n_1316), .Y(n_1362) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1334), .B(n_1252), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1310), .B(n_1245), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1311), .B(n_1296), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1311), .B(n_1296), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1338), .B(n_1268), .Y(n_1367) );
INVx2_ASAP7_75t_L g1368 ( .A(n_1328), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1327), .B(n_1288), .Y(n_1369) );
NAND2x1p5_ASAP7_75t_L g1370 ( .A(n_1320), .B(n_1264), .Y(n_1370) );
AND3x2_ASAP7_75t_L g1371 ( .A(n_1339), .B(n_1230), .C(n_1281), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1324), .B(n_1299), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1324), .B(n_1299), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1330), .B(n_1290), .Y(n_1374) );
HB1xp67_ASAP7_75t_L g1375 ( .A(n_1316), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1330), .B(n_1290), .Y(n_1376) );
BUFx3_ASAP7_75t_L g1377 ( .A(n_1320), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1331), .B(n_1293), .Y(n_1378) );
AND2x4_ASAP7_75t_L g1379 ( .A(n_1321), .B(n_1253), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1351), .B(n_1312), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1359), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1382 ( .A(n_1369), .B(n_1309), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1359), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1351), .B(n_1312), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1344), .B(n_1326), .Y(n_1385) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1368), .Y(n_1386) );
OR2x6_ASAP7_75t_L g1387 ( .A(n_1370), .B(n_1318), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1344), .B(n_1326), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1347), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1348), .B(n_1326), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1352), .B(n_1335), .Y(n_1391) );
OR2x2_ASAP7_75t_L g1392 ( .A(n_1378), .B(n_1309), .Y(n_1392) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1347), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1360), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1354), .Y(n_1395) );
BUFx2_ASAP7_75t_L g1396 ( .A(n_1350), .Y(n_1396) );
INVx2_ASAP7_75t_SL g1397 ( .A(n_1377), .Y(n_1397) );
NOR2xp33_ASAP7_75t_L g1398 ( .A(n_1346), .B(n_1292), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1365), .B(n_1366), .Y(n_1399) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1348), .B(n_1308), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1365), .B(n_1313), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1366), .B(n_1313), .Y(n_1402) );
OR2x2_ASAP7_75t_L g1403 ( .A(n_1362), .B(n_1308), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1372), .B(n_1337), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1372), .B(n_1337), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1358), .B(n_1219), .Y(n_1406) );
NOR2xp33_ASAP7_75t_L g1407 ( .A(n_1361), .B(n_1209), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1373), .B(n_1337), .Y(n_1408) );
NAND3xp33_ASAP7_75t_L g1409 ( .A(n_1396), .B(n_1375), .C(n_1314), .Y(n_1409) );
OAI22x1_ASAP7_75t_L g1410 ( .A1(n_1396), .A2(n_1370), .B1(n_1318), .B2(n_1379), .Y(n_1410) );
OAI22xp33_ASAP7_75t_R g1411 ( .A1(n_1407), .A2(n_1298), .B1(n_1293), .B2(n_1271), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1394), .B(n_1355), .Y(n_1412) );
NAND2x1_ASAP7_75t_SL g1413 ( .A(n_1385), .B(n_1379), .Y(n_1413) );
INVxp67_ASAP7_75t_L g1414 ( .A(n_1398), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1404), .B(n_1364), .Y(n_1415) );
INVxp67_ASAP7_75t_L g1416 ( .A(n_1406), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1403), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1392), .Y(n_1418) );
NAND2xp5_ASAP7_75t_SL g1419 ( .A(n_1397), .B(n_1370), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1399), .B(n_1374), .Y(n_1420) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_1382), .A2(n_1379), .B1(n_1314), .B2(n_1263), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_1387), .A2(n_1300), .B1(n_1261), .B2(n_1318), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g1423 ( .A1(n_1387), .A2(n_1298), .B1(n_1307), .B2(n_1377), .Y(n_1423) );
AOI211xp5_ASAP7_75t_SL g1424 ( .A1(n_1400), .A2(n_1144), .B(n_1274), .C(n_1264), .Y(n_1424) );
OAI322xp33_ASAP7_75t_L g1425 ( .A1(n_1382), .A2(n_1367), .A3(n_1353), .B1(n_1349), .B2(n_1356), .C1(n_1345), .C2(n_1357), .Y(n_1425) );
AOI21xp33_ASAP7_75t_SL g1426 ( .A1(n_1387), .A2(n_1371), .B(n_1307), .Y(n_1426) );
AOI22xp5_ASAP7_75t_L g1427 ( .A1(n_1405), .A2(n_1374), .B1(n_1376), .B2(n_1322), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1417), .Y(n_1428) );
INVx2_ASAP7_75t_L g1429 ( .A(n_1413), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1421), .B(n_1408), .Y(n_1430) );
O2A1O1Ixp5_ASAP7_75t_SL g1431 ( .A1(n_1414), .A2(n_1395), .B(n_1393), .C(n_1389), .Y(n_1431) );
O2A1O1Ixp33_ASAP7_75t_SL g1432 ( .A1(n_1424), .A2(n_1384), .B(n_1380), .C(n_1391), .Y(n_1432) );
AOI321xp33_ASAP7_75t_L g1433 ( .A1(n_1422), .A2(n_1343), .A3(n_1322), .B1(n_1266), .B2(n_1390), .C(n_1388), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1418), .Y(n_1434) );
AOI21xp33_ASAP7_75t_L g1435 ( .A1(n_1409), .A2(n_1294), .B(n_1273), .Y(n_1435) );
AOI32xp33_ASAP7_75t_L g1436 ( .A1(n_1424), .A2(n_1388), .A3(n_1402), .B1(n_1401), .B2(n_1408), .Y(n_1436) );
NAND2xp5_ASAP7_75t_SL g1437 ( .A(n_1410), .B(n_1274), .Y(n_1437) );
O2A1O1Ixp33_ASAP7_75t_L g1438 ( .A1(n_1426), .A2(n_1343), .B(n_1302), .C(n_1287), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_1411), .A2(n_1266), .B1(n_1254), .B2(n_1323), .Y(n_1439) );
OAI21xp33_ASAP7_75t_L g1440 ( .A1(n_1436), .A2(n_1423), .B(n_1416), .Y(n_1440) );
NAND4xp25_ASAP7_75t_SL g1441 ( .A(n_1439), .B(n_1427), .C(n_1412), .D(n_1420), .Y(n_1441) );
AOI211xp5_ASAP7_75t_L g1442 ( .A1(n_1432), .A2(n_1423), .B(n_1419), .C(n_1425), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1434), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1444 ( .A(n_1430), .B(n_1415), .Y(n_1444) );
NOR2x1_ASAP7_75t_L g1445 ( .A(n_1437), .B(n_1184), .Y(n_1445) );
OAI221xp5_ASAP7_75t_L g1446 ( .A1(n_1433), .A2(n_1269), .B1(n_1253), .B2(n_1255), .C(n_1336), .Y(n_1446) );
AOI211xp5_ASAP7_75t_L g1447 ( .A1(n_1441), .A2(n_1438), .B(n_1435), .C(n_1429), .Y(n_1447) );
NAND3xp33_ASAP7_75t_L g1448 ( .A(n_1442), .B(n_1431), .C(n_1428), .Y(n_1448) );
AOI221xp5_ASAP7_75t_L g1449 ( .A1(n_1440), .A2(n_1429), .B1(n_1381), .B2(n_1383), .C(n_1386), .Y(n_1449) );
BUFx12f_ASAP7_75t_L g1450 ( .A(n_1445), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1451 ( .A(n_1444), .B(n_1363), .Y(n_1451) );
BUFx6f_ASAP7_75t_L g1452 ( .A(n_1450), .Y(n_1452) );
NOR3xp33_ASAP7_75t_L g1453 ( .A(n_1448), .B(n_1446), .C(n_1443), .Y(n_1453) );
NOR5xp2_ASAP7_75t_L g1454 ( .A(n_1449), .B(n_1297), .C(n_1386), .D(n_1383), .E(n_1381), .Y(n_1454) );
OAI22xp5_ASAP7_75t_SL g1455 ( .A1(n_1452), .A2(n_1447), .B1(n_1451), .B2(n_1342), .Y(n_1455) );
AOI22xp5_ASAP7_75t_L g1456 ( .A1(n_1455), .A2(n_1453), .B1(n_1454), .B2(n_1269), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1457 ( .A1(n_1456), .A2(n_1305), .B1(n_1255), .B2(n_1304), .Y(n_1457) );
AOI21xp33_ASAP7_75t_L g1458 ( .A1(n_1457), .A2(n_1242), .B(n_1239), .Y(n_1458) );
OAI211xp5_ASAP7_75t_L g1459 ( .A1(n_1458), .A2(n_1148), .B(n_1206), .C(n_1207), .Y(n_1459) );
INVxp67_ASAP7_75t_L g1460 ( .A(n_1459), .Y(n_1460) );
AOI21xp5_ASAP7_75t_L g1461 ( .A1(n_1460), .A2(n_1291), .B(n_1278), .Y(n_1461) );
endmodule