module fake_jpeg_18391_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_51),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_77),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_61),
.B1(n_59),
.B2(n_45),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_49),
.B1(n_40),
.B2(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_62),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_92),
.Y(n_102)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_44),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_60),
.B(n_55),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_102),
.C(n_100),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_58),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_47),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_41),
.B1(n_39),
.B2(n_7),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_36),
.B1(n_10),
.B2(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_4),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_6),
.B1(n_16),
.B2(n_17),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_35),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_117),
.C(n_112),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_120),
.B(n_121),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_122),
.B1(n_126),
.B2(n_116),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_100),
.C(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_18),
.B(n_20),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_22),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_23),
.Y(n_136)
);


endmodule