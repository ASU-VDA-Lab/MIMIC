module fake_jpeg_6352_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_47),
.Y(n_62)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g89 ( 
.A(n_65),
.Y(n_89)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_28),
.B1(n_36),
.B2(n_30),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_28),
.B1(n_19),
.B2(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_80),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_74),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_28),
.B1(n_41),
.B2(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_30),
.B1(n_89),
.B2(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_84),
.Y(n_124)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_86),
.Y(n_126)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_92),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_23),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_33),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_34),
.C(n_26),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_36),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_28),
.B1(n_46),
.B2(n_19),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_19),
.B1(n_67),
.B2(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_21),
.Y(n_117)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_110),
.B1(n_125),
.B2(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_98),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_88),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_46),
.B1(n_53),
.B2(n_56),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_33),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_34),
.B(n_90),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_42),
.B1(n_39),
.B2(n_56),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_83),
.B1(n_75),
.B2(n_84),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_42),
.B1(n_26),
.B2(n_22),
.Y(n_125)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_127),
.A2(n_113),
.B1(n_95),
.B2(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_132),
.A2(n_32),
.B1(n_74),
.B2(n_35),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_133),
.A2(n_128),
.B1(n_27),
.B2(n_31),
.Y(n_183)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_137),
.A2(n_13),
.B(n_16),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_148),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_94),
.B1(n_88),
.B2(n_17),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_45),
.B(n_82),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_149),
.B(n_124),
.Y(n_177)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_72),
.B1(n_37),
.B2(n_44),
.Y(n_144)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_150),
.B1(n_154),
.B2(n_18),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_157),
.B1(n_126),
.B2(n_100),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_70),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_35),
.B(n_25),
.Y(n_149)
);

AO22x2_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_18),
.B1(n_29),
.B2(n_73),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_40),
.C(n_37),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_37),
.C(n_44),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_102),
.A2(n_20),
.B1(n_31),
.B2(n_27),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_124),
.B(n_20),
.C(n_17),
.Y(n_169)
);

AO22x2_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_18),
.B1(n_29),
.B2(n_73),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_70),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_79),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_75),
.B1(n_79),
.B2(n_77),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_21),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_108),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_120),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_159),
.A2(n_177),
.B(n_179),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_162),
.B1(n_169),
.B2(n_189),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_105),
.B1(n_126),
.B2(n_100),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_127),
.B1(n_77),
.B2(n_101),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_167),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_105),
.A3(n_121),
.B1(n_116),
.B2(n_108),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_74),
.B1(n_38),
.B2(n_2),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_187),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_122),
.B(n_106),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_181),
.B(n_44),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_106),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_38),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_101),
.B(n_20),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_31),
.B1(n_29),
.B2(n_40),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_155),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_74),
.B1(n_32),
.B2(n_12),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_154),
.B1(n_153),
.B2(n_137),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_138),
.B(n_32),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_147),
.C(n_140),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_194),
.B(n_196),
.Y(n_234)
);

AO21x2_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_144),
.B(n_150),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_168),
.B1(n_182),
.B2(n_181),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_206),
.C(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_152),
.B1(n_154),
.B2(n_150),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_140),
.B(n_158),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_211),
.B(n_217),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_154),
.C(n_146),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_150),
.B1(n_129),
.B2(n_151),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_209),
.B1(n_169),
.B2(n_188),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_151),
.B1(n_135),
.B2(n_145),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_174),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_212),
.B(n_218),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_40),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_221),
.B1(n_211),
.B2(n_163),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_0),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_179),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_167),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_166),
.B(n_38),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_213),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_15),
.A3(n_6),
.B1(n_7),
.B2(n_14),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_169),
.B(n_185),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_227),
.B(n_228),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_224),
.A2(n_170),
.B1(n_1),
.B2(n_2),
.Y(n_266)
);

OAI22x1_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_159),
.B1(n_175),
.B2(n_169),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_210),
.B1(n_207),
.B2(n_193),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_214),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_230),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_229),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_161),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_245),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_206),
.C(n_197),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_238),
.B(n_210),
.CI(n_216),
.CON(n_264),
.SN(n_264)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_241),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_200),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_159),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_202),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_203),
.A2(n_165),
.B1(n_170),
.B2(n_2),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_217),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_254),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_225),
.B(n_201),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_237),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_220),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_205),
.C(n_198),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_262),
.C(n_233),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_198),
.C(n_204),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_224),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_270),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_193),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_238),
.B1(n_248),
.B2(n_224),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_269),
.A2(n_244),
.B1(n_224),
.B2(n_246),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_276),
.C(n_286),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_242),
.C(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_260),
.B(n_252),
.Y(n_294)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_283),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_223),
.B1(n_227),
.B2(n_232),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_285),
.B1(n_257),
.B2(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_235),
.B1(n_242),
.B2(n_5),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_10),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_264),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_257),
.B(n_256),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_292),
.B(n_294),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_251),
.B(n_259),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_262),
.C(n_254),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_300),
.C(n_3),
.Y(n_308)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_6),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_250),
.C(n_255),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_264),
.B(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_284),
.B1(n_286),
.B2(n_272),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_302),
.B1(n_295),
.B2(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_284),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_306),
.B(n_307),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_10),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_7),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_315),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_310),
.B(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_6),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_4),
.Y(n_315)
);

INVx11_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_5),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_317),
.B(n_11),
.CI(n_13),
.CON(n_328),
.SN(n_328)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_288),
.B1(n_289),
.B2(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_320),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_295),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_300),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_322),
.A2(n_323),
.B(n_5),
.Y(n_325)
);

O2A1O1Ixp33_ASAP7_75t_SL g323 ( 
.A1(n_303),
.A2(n_304),
.B(n_314),
.C(n_4),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_326),
.B(n_327),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_324),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_329),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_11),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_11),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_321),
.C(n_316),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_332),
.A2(n_328),
.B(n_326),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_323),
.B(n_330),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_333),
.C(n_15),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_14),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_14),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_5),
.Y(n_340)
);


endmodule