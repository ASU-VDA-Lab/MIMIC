module fake_netlist_6_2054_n_1741 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1741);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1741;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_835;
wire n_242;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx2_ASAP7_75t_L g154 ( 
.A(n_23),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_37),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_49),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_56),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_59),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_35),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_49),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_39),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_86),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_2),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_33),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_52),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_90),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_36),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_28),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_58),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_59),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_31),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_43),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_95),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_45),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_30),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_98),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_89),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_33),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_74),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_63),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_55),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_17),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_35),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_120),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_96),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_56),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_72),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_27),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_54),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_133),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_116),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_118),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_24),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_51),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_43),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_24),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_62),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_79),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_51),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_91),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_145),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_30),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_88),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_100),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_135),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_143),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_3),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_66),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_4),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g228 ( 
.A(n_150),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_42),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_126),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_81),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_65),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_97),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_12),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_117),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_32),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_53),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_38),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_36),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_69),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_5),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_99),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_94),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_14),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_111),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_140),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_14),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_137),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_7),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_54),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_19),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_2),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_109),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_70),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_136),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_47),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_113),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_21),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_52),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_123),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_32),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_141),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_39),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_46),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_134),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_26),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_75),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_44),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_18),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_4),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_60),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_58),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_21),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_124),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_53),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_55),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_61),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_26),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_138),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_27),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_29),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_45),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_67),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_146),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_29),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_131),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_12),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_125),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_129),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_107),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_18),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_0),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_1),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_15),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_130),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_23),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_31),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_115),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_57),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_180),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_267),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_156),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_224),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_198),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_256),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_198),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_163),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_198),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_164),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_256),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_198),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_198),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_198),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_198),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_198),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_167),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_155),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_155),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_155),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_169),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_155),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_155),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_154),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_170),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_181),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_290),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_184),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_177),
.B(n_0),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_155),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_185),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_290),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_189),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_192),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_154),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_192),
.B(n_1),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_194),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_195),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_273),
.B(n_3),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_271),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_201),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_157),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_204),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_157),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_205),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_304),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_239),
.B(n_5),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_227),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_206),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_227),
.B(n_6),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_212),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_179),
.B(n_6),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_227),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_253),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_213),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_179),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_216),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_253),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_217),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_202),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_220),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_221),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_202),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_177),
.B(n_8),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_232),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_326),
.A2(n_306),
.B(n_211),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_319),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_310),
.B(n_286),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_319),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_235),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_310),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_232),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_362),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_340),
.B(n_235),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_314),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_307),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_337),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_308),
.A2(n_304),
.B1(n_172),
.B2(n_187),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_316),
.A2(n_188),
.B(n_173),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

BUFx8_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_320),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_321),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_311),
.A2(n_160),
.B1(n_215),
.B2(n_208),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_331),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_359),
.B(n_364),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_313),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_340),
.B(n_286),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_318),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_263),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_350),
.A2(n_306),
.B(n_211),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_344),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_359),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_344),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_377),
.B(n_240),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

BUFx8_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_365),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_309),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_381),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_410),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_315),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_357),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_389),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_380),
.B(n_240),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_389),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_317),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_410),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_324),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_422),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_380),
.B(n_240),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_328),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_395),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g474 ( 
.A(n_392),
.B(n_351),
.C(n_347),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_332),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_368),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_395),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_347),
.B1(n_351),
.B2(n_343),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_411),
.B(n_333),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_412),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_396),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_414),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

BUFx4f_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_411),
.B(n_334),
.Y(n_487)
);

XOR2x2_ASAP7_75t_L g488 ( 
.A(n_408),
.B(n_358),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_R g489 ( 
.A(n_426),
.B(n_440),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_411),
.B(n_335),
.Y(n_490)
);

BUFx4f_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_391),
.Y(n_492)
);

AND2x2_ASAP7_75t_SL g493 ( 
.A(n_380),
.B(n_173),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_411),
.B(n_338),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_440),
.B(n_341),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_411),
.B(n_345),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_411),
.B(n_348),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_389),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_440),
.B(n_352),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_440),
.B(n_354),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_438),
.B(n_356),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_388),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_391),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_394),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_389),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_389),
.B(n_360),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_380),
.A2(n_349),
.B1(n_353),
.B2(n_372),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_L g510 ( 
.A1(n_408),
.A2(n_165),
.B1(n_238),
.B2(n_258),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_366),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_396),
.B(n_263),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_391),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g517 ( 
.A(n_417),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_421),
.B(n_368),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_413),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_228),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_408),
.B(n_339),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_401),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_389),
.B(n_369),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_438),
.B(n_373),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_438),
.A2(n_349),
.B1(n_372),
.B2(n_353),
.Y(n_525)
);

OAI21xp33_ASAP7_75t_SL g526 ( 
.A1(n_435),
.A2(n_355),
.B(n_237),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_396),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_425),
.B(n_375),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_405),
.B(n_374),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_396),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_438),
.B(n_263),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_405),
.B(n_371),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_396),
.B(n_240),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

NOR2x1p5_ASAP7_75t_L g539 ( 
.A(n_435),
.B(n_289),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_401),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_438),
.B(n_418),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_429),
.B(n_196),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_432),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_391),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_415),
.Y(n_547)
);

CKINVDCx12_ASAP7_75t_R g548 ( 
.A(n_417),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_432),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_405),
.B(n_199),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_429),
.B(n_370),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_398),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_417),
.A2(n_358),
.B1(n_251),
.B2(n_218),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_420),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_378),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_437),
.B(n_370),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_429),
.B(n_394),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_378),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_429),
.B(n_231),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_429),
.B(n_244),
.Y(n_562)
);

BUFx6f_ASAP7_75t_SL g563 ( 
.A(n_429),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_437),
.A2(n_355),
.B1(n_249),
.B2(n_303),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_437),
.B(n_367),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_398),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_394),
.B(n_245),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_398),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_421),
.B(n_433),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_398),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_383),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_442),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_378),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_383),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_442),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_432),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_394),
.B(n_397),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_426),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_379),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_432),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_398),
.Y(n_584)
);

BUFx4f_ASAP7_75t_L g585 ( 
.A(n_383),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_441),
.B(n_199),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_394),
.B(n_247),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_394),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_397),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_421),
.B(n_158),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_L g591 ( 
.A(n_474),
.B(n_424),
.Y(n_591)
);

INVx8_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_447),
.B(n_397),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_557),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_557),
.Y(n_595)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_520),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_566),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_493),
.B(n_441),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_483),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_493),
.A2(n_383),
.B1(n_259),
.B2(n_208),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_560),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_493),
.A2(n_385),
.B1(n_260),
.B2(n_188),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_560),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_475),
.A2(n_272),
.B1(n_441),
.B2(n_421),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_457),
.B(n_422),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_520),
.Y(n_606)
);

BUFx6f_ASAP7_75t_SL g607 ( 
.A(n_478),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_575),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_511),
.B(n_441),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_483),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_575),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

BUFx5_ASAP7_75t_L g613 ( 
.A(n_573),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_543),
.A2(n_385),
.B(n_424),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_444),
.B(n_397),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_528),
.B(n_441),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_449),
.B(n_457),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_496),
.B(n_397),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_571),
.A2(n_491),
.B(n_585),
.C(n_486),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_456),
.B(n_441),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_582),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_459),
.A2(n_225),
.B1(n_269),
.B2(n_248),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_465),
.B(n_250),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_527),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_500),
.B(n_264),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_502),
.B(n_397),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_443),
.B(n_477),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_530),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_443),
.B(n_419),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_530),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_474),
.B(n_581),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_508),
.B(n_419),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_450),
.B(n_442),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_450),
.B(n_442),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_477),
.B(n_419),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_506),
.B(n_446),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_454),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_446),
.B(n_419),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_582),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_454),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_499),
.A2(n_297),
.B1(n_305),
.B2(n_281),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_451),
.B(n_458),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_555),
.B(n_385),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_451),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_525),
.B(n_266),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_499),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_458),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_469),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_507),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_509),
.B(n_291),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_545),
.A2(n_383),
.B1(n_241),
.B2(n_246),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_518),
.B(n_436),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_469),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_507),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_472),
.B(n_419),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_563),
.Y(n_656)
);

BUFx5_ASAP7_75t_L g657 ( 
.A(n_573),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_523),
.B(n_419),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_515),
.B(n_426),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_486),
.B(n_260),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_479),
.B(n_293),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_486),
.A2(n_409),
.B(n_436),
.C(n_284),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_472),
.B(n_398),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_481),
.B(n_398),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_515),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_481),
.Y(n_666)
);

BUFx8_ASAP7_75t_L g667 ( 
.A(n_449),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_566),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_518),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_526),
.B(n_159),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_524),
.B(n_296),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_482),
.Y(n_673)
);

AND2x2_ASAP7_75t_SL g674 ( 
.A(n_491),
.B(n_585),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_526),
.B(n_161),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_482),
.B(n_484),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_484),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_590),
.B(n_162),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_501),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_501),
.B(n_398),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_466),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_534),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_491),
.A2(n_233),
.B1(n_186),
.B2(n_200),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_534),
.B(n_399),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_540),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_540),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_487),
.B(n_199),
.Y(n_687)
);

INVxp33_ASAP7_75t_L g688 ( 
.A(n_521),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_513),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_513),
.B(n_436),
.Y(n_690)
);

INVxp33_ASAP7_75t_L g691 ( 
.A(n_521),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_480),
.B(n_199),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_576),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_545),
.A2(n_237),
.B1(n_241),
.B2(n_246),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_532),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_550),
.B(n_166),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_513),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_513),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_576),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_539),
.A2(n_228),
.B1(n_248),
.B2(n_233),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_544),
.B(n_168),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_549),
.A2(n_433),
.B(n_436),
.C(n_303),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_490),
.B(n_422),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_495),
.B(n_442),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_549),
.A2(n_259),
.B1(n_249),
.B2(n_261),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_552),
.B(n_399),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_585),
.B(n_442),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_552),
.B(n_399),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_570),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_588),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_399),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_532),
.B(n_442),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_588),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_532),
.B(n_442),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_577),
.B(n_399),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_579),
.A2(n_261),
.B1(n_278),
.B2(n_285),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_579),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_583),
.B(n_399),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_583),
.B(n_399),
.Y(n_720)
);

INVx8_ASAP7_75t_L g721 ( 
.A(n_520),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_589),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_L g723 ( 
.A(n_586),
.B(n_433),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_466),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_589),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_539),
.B(n_399),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_512),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_460),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_559),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_520),
.A2(n_214),
.B1(n_302),
.B2(n_295),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_497),
.B(n_442),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_498),
.B(n_240),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_452),
.B(n_399),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_452),
.B(n_403),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_532),
.B(n_240),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_510),
.B(n_209),
.C(n_191),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_561),
.B(n_171),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_562),
.B(n_174),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_452),
.B(n_403),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_452),
.B(n_403),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_489),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_564),
.B(n_178),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_512),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_563),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_558),
.B(n_186),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_514),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_531),
.B(n_175),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_529),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_563),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_580),
.A2(n_409),
.B(n_207),
.C(n_214),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_452),
.B(n_462),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_533),
.B(n_236),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_568),
.B(n_403),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_587),
.B(n_176),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_514),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_519),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_462),
.B(n_200),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_505),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_522),
.B(n_182),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_462),
.B(n_403),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_627),
.A2(n_503),
.B(n_453),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_683),
.A2(n_517),
.B(n_519),
.C(n_556),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_613),
.B(n_462),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_593),
.B(n_462),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_670),
.B(n_462),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_644),
.Y(n_766)
);

O2A1O1Ixp5_ASAP7_75t_L g767 ( 
.A1(n_593),
.A2(n_547),
.B(n_542),
.C(n_556),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_613),
.B(n_505),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_728),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_678),
.B(n_462),
.Y(n_770)
);

OAI21xp33_ASAP7_75t_L g771 ( 
.A1(n_678),
.A2(n_488),
.B(n_554),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_644),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_600),
.A2(n_554),
.B1(n_517),
.B2(n_269),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_600),
.A2(n_302),
.B1(n_207),
.B2(n_219),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_647),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_694),
.A2(n_488),
.B1(n_298),
.B2(n_278),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_605),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_706),
.A2(n_492),
.B(n_471),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_707),
.A2(n_453),
.B(n_448),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_648),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_741),
.B(n_748),
.C(n_759),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_648),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_612),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_707),
.A2(n_453),
.B(n_448),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_591),
.B(n_471),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_612),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_701),
.B(n_471),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_671),
.A2(n_537),
.B(n_538),
.C(n_542),
.Y(n_788)
);

INVx3_ASAP7_75t_SL g789 ( 
.A(n_681),
.Y(n_789)
);

AOI21x1_ASAP7_75t_L g790 ( 
.A1(n_633),
.A2(n_634),
.B(n_726),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_708),
.A2(n_470),
.B(n_448),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_701),
.B(n_492),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_669),
.B(n_548),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_671),
.A2(n_257),
.B(n_295),
.C(n_230),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_597),
.B(n_643),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_659),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_653),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_729),
.B(n_492),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_612),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_747),
.B(n_516),
.Y(n_800)
);

NOR2x2_ASAP7_75t_L g801 ( 
.A(n_659),
.B(n_548),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_617),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_612),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_747),
.B(n_516),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_665),
.B(n_522),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_675),
.A2(n_225),
.B(n_226),
.C(n_219),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_752),
.B(n_478),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_754),
.B(n_516),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_754),
.B(n_536),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_666),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_659),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_711),
.A2(n_553),
.B(n_470),
.Y(n_812)
);

O2A1O1Ixp5_ASAP7_75t_L g813 ( 
.A1(n_602),
.A2(n_547),
.B(n_537),
.C(n_538),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_716),
.A2(n_553),
.B(n_470),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_666),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_619),
.A2(n_409),
.B(n_536),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_668),
.B(n_536),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_667),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_660),
.A2(n_693),
.B1(n_699),
.B2(n_709),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_673),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_631),
.B(n_478),
.Y(n_821)
);

INVx6_ASAP7_75t_L g822 ( 
.A(n_656),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_719),
.A2(n_584),
.B(n_553),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_737),
.B(n_565),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_633),
.A2(n_455),
.B(n_445),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_724),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_720),
.A2(n_584),
.B(n_546),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_660),
.A2(n_738),
.B1(n_737),
.B2(n_599),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_693),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_673),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_699),
.B(n_478),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_614),
.A2(n_584),
.B(n_546),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_677),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_738),
.B(n_565),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_696),
.B(n_565),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_749),
.B(n_226),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_613),
.B(n_505),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_677),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_712),
.A2(n_505),
.B(n_546),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_709),
.B(n_445),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_712),
.A2(n_505),
.B(n_546),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_679),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_715),
.A2(n_546),
.B(n_572),
.Y(n_843)
);

AO21x1_ASAP7_75t_L g844 ( 
.A1(n_598),
.A2(n_255),
.B(n_257),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_652),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_662),
.A2(n_409),
.B(n_473),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_714),
.B(n_718),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_675),
.A2(n_292),
.B(n_298),
.C(n_294),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_714),
.B(n_455),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_679),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_652),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_613),
.B(n_569),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_696),
.A2(n_252),
.B(n_276),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_718),
.B(n_461),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_703),
.B(n_541),
.C(n_255),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_736),
.B(n_541),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_661),
.B(n_569),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_710),
.Y(n_858)
);

AOI21xp33_ASAP7_75t_L g859 ( 
.A1(n_650),
.A2(n_230),
.B(n_284),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_690),
.Y(n_860)
);

AO21x1_ASAP7_75t_L g861 ( 
.A1(n_609),
.A2(n_285),
.B(n_292),
.Y(n_861)
);

INVx11_ASAP7_75t_L g862 ( 
.A(n_667),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_592),
.Y(n_863)
);

O2A1O1Ixp5_ASAP7_75t_L g864 ( 
.A1(n_618),
.A2(n_463),
.B(n_461),
.C(n_464),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_632),
.B(n_463),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_715),
.A2(n_569),
.B(n_572),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_613),
.B(n_569),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_632),
.B(n_464),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_688),
.B(n_691),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_658),
.B(n_467),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_700),
.B(n_569),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_658),
.A2(n_467),
.B(n_468),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_753),
.A2(n_572),
.B(n_567),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_713),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_682),
.B(n_468),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_753),
.A2(n_758),
.B(n_635),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_592),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_685),
.B(n_473),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_722),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_629),
.A2(n_572),
.B(n_567),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_695),
.A2(n_572),
.B(n_567),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_744),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_742),
.A2(n_622),
.B(n_645),
.C(n_745),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_695),
.A2(n_567),
.B(n_476),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_694),
.A2(n_210),
.B(n_223),
.Y(n_885)
);

AO21x1_ASAP7_75t_L g886 ( 
.A1(n_616),
.A2(n_294),
.B(n_379),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_686),
.B(n_476),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_725),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_607),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_689),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_637),
.B(n_183),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_640),
.B(n_190),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_615),
.B(n_485),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_615),
.A2(n_485),
.B(n_504),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_626),
.B(n_494),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_690),
.A2(n_567),
.B(n_494),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_626),
.A2(n_504),
.B(n_535),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_613),
.B(n_578),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_646),
.B(n_193),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_636),
.B(n_535),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_723),
.A2(n_434),
.B(n_427),
.C(n_386),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_757),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_634),
.A2(n_567),
.B(n_574),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_610),
.B(n_236),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_594),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_757),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_735),
.A2(n_578),
.B(n_574),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_624),
.B(n_236),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_697),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_638),
.A2(n_535),
.B(n_382),
.Y(n_910)
);

BUFx4f_ASAP7_75t_L g911 ( 
.A(n_592),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_705),
.A2(n_717),
.B1(n_651),
.B2(n_674),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_642),
.A2(n_404),
.B(n_407),
.C(n_379),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_698),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_649),
.B(n_535),
.Y(n_915)
);

O2A1O1Ixp5_ASAP7_75t_L g916 ( 
.A1(n_750),
.A2(n_407),
.B(n_382),
.C(n_402),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_595),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_676),
.A2(n_404),
.B(n_407),
.C(n_382),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_657),
.B(n_674),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_654),
.B(n_197),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_704),
.A2(n_578),
.B(n_574),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_657),
.B(n_578),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_651),
.B(n_535),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_656),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_657),
.B(n_535),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_657),
.B(n_535),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_655),
.A2(n_386),
.B(n_402),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_744),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_731),
.A2(n_574),
.B(n_403),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_733),
.A2(n_403),
.B(n_416),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_628),
.A2(n_403),
.B1(n_416),
.B2(n_434),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_734),
.A2(n_403),
.B(n_416),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_630),
.A2(n_434),
.B(n_427),
.C(n_386),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_601),
.Y(n_934)
);

AND2x6_ASAP7_75t_L g935 ( 
.A(n_751),
.B(n_416),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_739),
.A2(n_416),
.B(n_434),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_657),
.B(n_416),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_596),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_596),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_740),
.A2(n_416),
.B(n_387),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_L g941 ( 
.A(n_657),
.B(n_416),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_596),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_760),
.A2(n_416),
.B(n_387),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_623),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_601),
.B(n_431),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_941),
.A2(n_620),
.B(n_606),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_763),
.A2(n_721),
.B(n_606),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_912),
.B(n_705),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_771),
.A2(n_692),
.B(n_604),
.C(n_732),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_SL g950 ( 
.A1(n_794),
.A2(n_687),
.B(n_672),
.C(n_625),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_SL g951 ( 
.A1(n_821),
.A2(n_702),
.B(n_611),
.C(n_621),
.Y(n_951)
);

OAI22xp33_ASAP7_75t_L g952 ( 
.A1(n_773),
.A2(n_777),
.B1(n_828),
.B2(n_802),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_793),
.B(n_607),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_786),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_826),
.B(n_730),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_912),
.B(n_717),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_796),
.B(n_606),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_776),
.A2(n_721),
.B1(n_611),
.B2(n_621),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_807),
.B(n_641),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_848),
.A2(n_603),
.B(n_639),
.C(n_608),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_845),
.B(n_608),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_766),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_772),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_781),
.A2(n_721),
.B1(n_639),
.B2(n_755),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_789),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_845),
.B(n_727),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_883),
.A2(n_684),
.B(n_664),
.C(n_680),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_775),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_789),
.Y(n_969)
);

NAND2x1p5_ASAP7_75t_L g970 ( 
.A(n_803),
.B(n_727),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_863),
.B(n_663),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_831),
.B(n_743),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_769),
.Y(n_973)
);

AO22x1_ASAP7_75t_L g974 ( 
.A1(n_793),
.A2(n_275),
.B1(n_229),
.B2(n_234),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_859),
.A2(n_756),
.B(n_746),
.C(n_288),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_SL g976 ( 
.A1(n_776),
.A2(n_811),
.B1(n_805),
.B2(n_818),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_889),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_769),
.B(n_746),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_795),
.B(n_756),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_SL g980 ( 
.A(n_863),
.B(n_203),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_L g981 ( 
.A(n_944),
.B(n_64),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_891),
.B(n_71),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_SL g983 ( 
.A1(n_835),
.A2(n_404),
.B(n_387),
.C(n_393),
.Y(n_983)
);

NOR2x1_ASAP7_75t_L g984 ( 
.A(n_882),
.B(n_393),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_SL g985 ( 
.A1(n_835),
.A2(n_406),
.B(n_393),
.C(n_400),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_904),
.B(n_236),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_767),
.A2(n_400),
.B(n_402),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_780),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_781),
.B(n_242),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_847),
.B(n_400),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_853),
.B(n_243),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_820),
.B(n_406),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_898),
.A2(n_430),
.B(n_428),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_898),
.A2(n_430),
.B(n_428),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_806),
.A2(n_406),
.B(n_427),
.C(n_431),
.Y(n_995)
);

AO22x1_ASAP7_75t_L g996 ( 
.A1(n_855),
.A2(n_254),
.B1(n_262),
.B2(n_265),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_774),
.A2(n_283),
.B1(n_270),
.B2(n_274),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_767),
.A2(n_813),
.B(n_864),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_831),
.B(n_299),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_782),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_922),
.A2(n_430),
.B(n_428),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_855),
.A2(n_431),
.B(n_430),
.C(n_428),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_858),
.B(n_431),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_928),
.B(n_924),
.Y(n_1004)
);

BUFx4f_ASAP7_75t_L g1005 ( 
.A(n_863),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_830),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_922),
.A2(n_423),
.B(n_82),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_869),
.B(n_268),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_863),
.B(n_80),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_761),
.A2(n_423),
.B(n_83),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_L g1011 ( 
.A(n_891),
.B(n_78),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_836),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_892),
.A2(n_899),
.B(n_920),
.C(n_762),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_SL g1014 ( 
.A1(n_856),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_L g1015 ( 
.A(n_892),
.B(n_301),
.C(n_300),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_860),
.B(n_287),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_808),
.A2(n_423),
.B(n_114),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_809),
.A2(n_423),
.B(n_119),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_838),
.B(n_282),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_842),
.B(n_152),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_801),
.Y(n_1021)
);

AND2x2_ASAP7_75t_SL g1022 ( 
.A(n_911),
.B(n_8),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_877),
.B(n_151),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_786),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_899),
.B(n_10),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_L g1026 ( 
.A(n_920),
.B(n_885),
.C(n_851),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_836),
.A2(n_908),
.B1(n_874),
.B2(n_879),
.C(n_888),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_797),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_902),
.B(n_10),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_860),
.B(n_11),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_824),
.A2(n_144),
.B(n_142),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_822),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_906),
.B(n_11),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_764),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_834),
.A2(n_837),
.B(n_768),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_923),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_1036)
);

AO32x2_ASAP7_75t_L g1037 ( 
.A1(n_819),
.A2(n_19),
.A3(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_890),
.B(n_20),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_768),
.A2(n_139),
.B(n_128),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_829),
.B(n_22),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_914),
.A2(n_25),
.B1(n_34),
.B2(n_38),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_810),
.B(n_40),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_786),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_815),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_837),
.A2(n_76),
.B(n_110),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_786),
.B(n_105),
.Y(n_1046)
);

BUFx12f_ASAP7_75t_L g1047 ( 
.A(n_822),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_813),
.A2(n_104),
.B(n_93),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_933),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_852),
.A2(n_92),
.B(n_87),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_862),
.Y(n_1051)
);

CKINVDCx16_ASAP7_75t_R g1052 ( 
.A(n_877),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_833),
.Y(n_1053)
);

AND2x6_ASAP7_75t_SL g1054 ( 
.A(n_871),
.B(n_44),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_770),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_SL g1056 ( 
.A(n_861),
.B(n_48),
.C(n_50),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_783),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_829),
.B(n_50),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_850),
.Y(n_1059)
);

AO32x2_ASAP7_75t_L g1060 ( 
.A1(n_803),
.A2(n_57),
.A3(n_77),
.B1(n_85),
.B2(n_882),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_917),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_871),
.A2(n_919),
.B1(n_857),
.B2(n_909),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_829),
.B(n_919),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_829),
.B(n_909),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_877),
.Y(n_1065)
);

INVxp67_ASAP7_75t_L g1066 ( 
.A(n_783),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_857),
.A2(n_792),
.B(n_787),
.C(n_876),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_877),
.B(n_938),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_799),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_SL g1070 ( 
.A1(n_911),
.A2(n_938),
.B1(n_939),
.B2(n_942),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_938),
.B(n_939),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_799),
.B(n_938),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_939),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_939),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_942),
.B(n_765),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_785),
.B(n_800),
.Y(n_1076)
);

OA22x2_ASAP7_75t_L g1077 ( 
.A1(n_765),
.A2(n_816),
.B1(n_934),
.B2(n_905),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_804),
.A2(n_788),
.B(n_900),
.C(n_910),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_852),
.A2(n_867),
.B(n_926),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_942),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_817),
.B(n_887),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_875),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_878),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_942),
.A2(n_886),
.B1(n_844),
.B2(n_915),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_945),
.Y(n_1085)
);

BUFx12f_ASAP7_75t_L g1086 ( 
.A(n_935),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1082),
.B(n_798),
.Y(n_1087)
);

BUFx8_ASAP7_75t_L g1088 ( 
.A(n_973),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1067),
.A2(n_893),
.B(n_895),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_1078),
.A2(n_1076),
.A3(n_967),
.B(n_1035),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_1010),
.A2(n_901),
.A3(n_832),
.B(n_865),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1013),
.A2(n_790),
.B(n_897),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1025),
.A2(n_918),
.B(n_913),
.C(n_896),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1079),
.A2(n_778),
.B(n_825),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_946),
.A2(n_870),
.B(n_868),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1027),
.B(n_925),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_957),
.B(n_867),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1083),
.B(n_849),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_991),
.A2(n_935),
.B1(n_945),
.B2(n_937),
.Y(n_1099)
);

AOI211x1_ASAP7_75t_L g1100 ( 
.A1(n_952),
.A2(n_846),
.B(n_927),
.C(n_943),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_989),
.A2(n_916),
.B(n_937),
.C(n_872),
.Y(n_1101)
);

AO31x2_ASAP7_75t_L g1102 ( 
.A1(n_949),
.A2(n_1017),
.A3(n_1018),
.B(n_956),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_957),
.B(n_841),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_977),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_962),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_948),
.A2(n_823),
.A3(n_791),
.B(n_812),
.Y(n_1106)
);

BUFx10_ASAP7_75t_L g1107 ( 
.A(n_953),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_948),
.A2(n_956),
.A3(n_1063),
.B(n_958),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_947),
.A2(n_779),
.B(n_784),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_963),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_978),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_1046),
.A2(n_840),
.B(n_854),
.C(n_839),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_982),
.A2(n_843),
.B(n_866),
.C(n_921),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_1015),
.B(n_931),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1029),
.Y(n_1115)
);

AO21x1_ASAP7_75t_L g1116 ( 
.A1(n_1048),
.A2(n_894),
.B(n_884),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_972),
.A2(n_814),
.B(n_827),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_958),
.A2(n_873),
.A3(n_880),
.B(n_929),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1062),
.A2(n_940),
.B(n_936),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1051),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1008),
.A2(n_935),
.B1(n_907),
.B2(n_932),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_979),
.B(n_930),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_1047),
.B(n_881),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_988),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1065),
.Y(n_1125)
);

INVx3_ASAP7_75t_SL g1126 ( 
.A(n_965),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1006),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_950),
.A2(n_903),
.B(n_864),
.Y(n_1128)
);

INVx3_ASAP7_75t_SL g1129 ( 
.A(n_969),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_959),
.A2(n_916),
.B(n_935),
.C(n_1036),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_975),
.A2(n_1020),
.A3(n_1036),
.B(n_994),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1011),
.A2(n_935),
.B(n_1026),
.C(n_1048),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_986),
.B(n_1022),
.Y(n_1133)
);

BUFx8_ASAP7_75t_SL g1134 ( 
.A(n_1032),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1012),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1014),
.B(n_996),
.C(n_1041),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_976),
.A2(n_955),
.B1(n_1016),
.B2(n_1021),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1077),
.A2(n_964),
.B(n_1030),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_998),
.A2(n_1081),
.B(n_951),
.Y(n_1139)
);

OAI22x1_ASAP7_75t_L g1140 ( 
.A1(n_1033),
.A2(n_1058),
.B1(n_1040),
.B2(n_999),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1068),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_SL g1142 ( 
.A1(n_1020),
.A2(n_983),
.B(n_985),
.C(n_1042),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_961),
.A2(n_1084),
.B(n_960),
.Y(n_1143)
);

NOR2x1_ASAP7_75t_SL g1144 ( 
.A(n_1086),
.B(n_971),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1019),
.B(n_1038),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_957),
.B(n_1009),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_981),
.A2(n_980),
.B1(n_997),
.B2(n_1019),
.Y(n_1147)
);

AOI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_997),
.A2(n_1044),
.B(n_1059),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_998),
.A2(n_990),
.B(n_1007),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_990),
.A2(n_1064),
.B(n_966),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1075),
.A2(n_1009),
.B1(n_1023),
.B2(n_1052),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1023),
.A2(n_1004),
.B1(n_1068),
.B2(n_1071),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_974),
.A2(n_1055),
.B1(n_1034),
.B2(n_1049),
.C(n_1056),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_987),
.A2(n_1001),
.B(n_993),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_1073),
.B(n_1074),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_987),
.A2(n_970),
.B(n_992),
.Y(n_1157)
);

AO32x2_ASAP7_75t_L g1158 ( 
.A1(n_1037),
.A2(n_1060),
.A3(n_1073),
.B1(n_1054),
.B2(n_992),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_966),
.A2(n_1003),
.B(n_1085),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_SL g1160 ( 
.A(n_1005),
.B(n_1004),
.Y(n_1160)
);

AO21x2_ASAP7_75t_L g1161 ( 
.A1(n_1031),
.A2(n_1039),
.B(n_1050),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_968),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1000),
.A2(n_1028),
.B(n_1053),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1002),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1045),
.A2(n_1005),
.B(n_995),
.C(n_1066),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_SL g1166 ( 
.A(n_1070),
.B(n_1080),
.C(n_1069),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1057),
.B(n_1043),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1074),
.B(n_1072),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_954),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_984),
.A2(n_971),
.B(n_970),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_971),
.A2(n_954),
.B(n_1024),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1024),
.Y(n_1172)
);

OAI22x1_ASAP7_75t_L g1173 ( 
.A1(n_1037),
.A2(n_1025),
.B1(n_554),
.B2(n_521),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1037),
.A2(n_1025),
.B(n_771),
.C(n_1013),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1060),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_1060),
.A2(n_771),
.B1(n_392),
.B2(n_474),
.C(n_510),
.Y(n_1176)
);

AO32x2_ASAP7_75t_L g1177 ( 
.A1(n_1036),
.A2(n_976),
.A3(n_774),
.B1(n_773),
.B2(n_602),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_965),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1013),
.A2(n_771),
.B(n_1025),
.C(n_678),
.Y(n_1179)
);

AOI31xp67_ASAP7_75t_L g1180 ( 
.A1(n_1077),
.A2(n_620),
.A3(n_1062),
.B(n_609),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1061),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1079),
.A2(n_778),
.B(n_816),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1061),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1082),
.B(n_741),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1013),
.A2(n_771),
.B(n_1025),
.C(n_678),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1067),
.A2(n_941),
.B(n_763),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1061),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1067),
.A2(n_941),
.B(n_763),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1013),
.A2(n_771),
.B(n_1025),
.C(n_678),
.Y(n_1189)
);

BUFx5_ASAP7_75t_L g1190 ( 
.A(n_1086),
.Y(n_1190)
);

NOR2x1_ASAP7_75t_L g1191 ( 
.A(n_965),
.B(n_969),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1079),
.A2(n_778),
.B(n_816),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1022),
.A2(n_548),
.B1(n_517),
.B2(n_521),
.Y(n_1193)
);

AOI221x1_ASAP7_75t_L g1194 ( 
.A1(n_1025),
.A2(n_771),
.B1(n_1048),
.B2(n_1036),
.C(n_392),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1079),
.A2(n_778),
.B(n_816),
.Y(n_1195)
);

AO21x1_ASAP7_75t_L g1196 ( 
.A1(n_1013),
.A2(n_1025),
.B(n_1048),
.Y(n_1196)
);

CKINVDCx16_ASAP7_75t_R g1197 ( 
.A(n_977),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1013),
.A2(n_828),
.B(n_1062),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_SL g1199 ( 
.A(n_1047),
.B(n_728),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1025),
.A2(n_771),
.B1(n_311),
.B2(n_307),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_998),
.A2(n_1048),
.B(n_1067),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1067),
.A2(n_941),
.B(n_763),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1067),
.A2(n_886),
.A3(n_844),
.B(n_1078),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1013),
.A2(n_771),
.B(n_1025),
.C(n_678),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1082),
.B(n_741),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1061),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_978),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_948),
.A2(n_912),
.B1(n_828),
.B2(n_956),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1013),
.A2(n_771),
.B(n_1025),
.C(n_678),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1082),
.B(n_741),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1061),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1061),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1067),
.A2(n_886),
.A3(n_844),
.B(n_1078),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_973),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1082),
.B(n_741),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1067),
.A2(n_941),
.B(n_763),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_973),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_SL g1218 ( 
.A1(n_947),
.A2(n_1049),
.B(n_1013),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1013),
.A2(n_828),
.B(n_1062),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_973),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1067),
.A2(n_941),
.B(n_763),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1047),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_957),
.B(n_1068),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1067),
.A2(n_941),
.B(n_763),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1176),
.A2(n_1173),
.B1(n_1136),
.B2(n_1196),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1198),
.A2(n_1219),
.B1(n_1193),
.B2(n_1140),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1207),
.A2(n_1179),
.B1(n_1189),
.B2(n_1209),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1175),
.A2(n_1133),
.B1(n_1208),
.B2(n_1111),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1104),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1185),
.A2(n_1204),
.B1(n_1200),
.B2(n_1137),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1088),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1153),
.A2(n_1145),
.B1(n_1147),
.B2(n_1218),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_SL g1233 ( 
.A1(n_1201),
.A2(n_1158),
.B1(n_1160),
.B2(n_1115),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1105),
.Y(n_1234)
);

INVx6_ASAP7_75t_L g1235 ( 
.A(n_1088),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1110),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1151),
.A2(n_1146),
.B1(n_1152),
.B2(n_1166),
.Y(n_1237)
);

CKINVDCx6p67_ASAP7_75t_R g1238 ( 
.A(n_1126),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1096),
.A2(n_1210),
.B1(n_1184),
.B2(n_1205),
.Y(n_1239)
);

BUFx4_ASAP7_75t_R g1240 ( 
.A(n_1134),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1194),
.A2(n_1215),
.B1(n_1087),
.B2(n_1098),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1197),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1214),
.A2(n_1174),
.B1(n_1132),
.B2(n_1220),
.Y(n_1243)
);

BUFx4_ASAP7_75t_SL g1244 ( 
.A(n_1120),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1156),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1097),
.B(n_1223),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1217),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1222),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1222),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1114),
.A2(n_1103),
.B1(n_1138),
.B2(n_1148),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1103),
.A2(n_1107),
.B1(n_1135),
.B2(n_1164),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1092),
.A2(n_1183),
.B1(n_1212),
.B2(n_1211),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1099),
.A2(n_1187),
.B1(n_1181),
.B2(n_1127),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1158),
.A2(n_1177),
.B1(n_1186),
.B2(n_1221),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1206),
.A2(n_1122),
.B1(n_1162),
.B2(n_1167),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1129),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1163),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1172),
.Y(n_1258)
);

CKINVDCx11_ASAP7_75t_R g1259 ( 
.A(n_1222),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1125),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1178),
.Y(n_1261)
);

OAI22x1_ASAP7_75t_SL g1262 ( 
.A1(n_1199),
.A2(n_1141),
.B1(n_1191),
.B2(n_1190),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1125),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1169),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1141),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1100),
.A2(n_1168),
.B1(n_1170),
.B2(n_1121),
.Y(n_1266)
);

CKINVDCx6p67_ASAP7_75t_R g1267 ( 
.A(n_1190),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1143),
.A2(n_1161),
.B1(n_1190),
.B2(n_1139),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1155),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1158),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1190),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1165),
.A2(n_1093),
.B1(n_1216),
.B2(n_1202),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1157),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1171),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1108),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1089),
.A2(n_1150),
.B1(n_1159),
.B2(n_1116),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1123),
.B(n_1188),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1144),
.B(n_1177),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1090),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1177),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1224),
.A2(n_1149),
.B1(n_1119),
.B2(n_1095),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1154),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1130),
.A2(n_1113),
.B1(n_1101),
.B2(n_1128),
.Y(n_1283)
);

CKINVDCx6p67_ASAP7_75t_R g1284 ( 
.A(n_1142),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1203),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1117),
.A2(n_1195),
.B1(n_1182),
.B2(n_1192),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1109),
.A2(n_1094),
.B1(n_1102),
.B2(n_1180),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1203),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1102),
.A2(n_1131),
.B1(n_1213),
.B2(n_1112),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1213),
.B(n_1131),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1131),
.A2(n_1118),
.B1(n_1091),
.B2(n_1106),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1106),
.A2(n_771),
.B1(n_1176),
.B2(n_1025),
.Y(n_1292)
);

INVx8_ASAP7_75t_L g1293 ( 
.A(n_1106),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1091),
.A2(n_771),
.B1(n_1176),
.B2(n_1025),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1091),
.B(n_1207),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1136),
.A2(n_771),
.B1(n_1025),
.B2(n_1176),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1193),
.A2(n_517),
.B1(n_1025),
.B2(n_1022),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1176),
.A2(n_956),
.B1(n_948),
.B2(n_1194),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1176),
.A2(n_956),
.B1(n_948),
.B2(n_1194),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1120),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1193),
.A2(n_517),
.B1(n_1025),
.B2(n_1022),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1223),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1124),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1124),
.Y(n_1304)
);

BUFx4f_ASAP7_75t_L g1305 ( 
.A(n_1222),
.Y(n_1305)
);

BUFx8_ASAP7_75t_L g1306 ( 
.A(n_1222),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1156),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1136),
.A2(n_771),
.B1(n_1025),
.B2(n_1176),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1136),
.A2(n_771),
.B1(n_1025),
.B2(n_1176),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1200),
.A2(n_771),
.B1(n_395),
.B2(n_311),
.Y(n_1310)
);

BUFx4f_ASAP7_75t_SL g1311 ( 
.A(n_1104),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1104),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1120),
.Y(n_1313)
);

INVx3_ASAP7_75t_SL g1314 ( 
.A(n_1120),
.Y(n_1314)
);

BUFx10_ASAP7_75t_L g1315 ( 
.A(n_1120),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1088),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1207),
.A2(n_1179),
.B1(n_1189),
.B2(n_1185),
.Y(n_1317)
);

BUFx2_ASAP7_75t_SL g1318 ( 
.A(n_1104),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1120),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1156),
.Y(n_1320)
);

OAI21xp33_ASAP7_75t_L g1321 ( 
.A1(n_1179),
.A2(n_771),
.B(n_1025),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1133),
.B(n_1115),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1156),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1207),
.A2(n_1179),
.B1(n_1189),
.B2(n_1185),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1193),
.A2(n_517),
.B1(n_1025),
.B2(n_1022),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1104),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1133),
.B(n_1115),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1176),
.A2(n_771),
.B1(n_1025),
.B2(n_1173),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1133),
.B(n_1115),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1176),
.A2(n_956),
.B1(n_948),
.B2(n_1194),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1193),
.A2(n_517),
.B1(n_1025),
.B2(n_1022),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1207),
.A2(n_1179),
.B1(n_1189),
.B2(n_1185),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1193),
.A2(n_517),
.B1(n_1025),
.B2(n_1022),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1214),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1124),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1124),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1088),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1089),
.A2(n_1188),
.B(n_1186),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1120),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1104),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1285),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1283),
.A2(n_1291),
.A3(n_1272),
.B(n_1288),
.Y(n_1342)
);

AOI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1321),
.A2(n_1308),
.B(n_1296),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1279),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1267),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1322),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1295),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1273),
.B(n_1278),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1275),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1290),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1270),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1327),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1270),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1280),
.B(n_1233),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1273),
.B(n_1282),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1233),
.B(n_1254),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1254),
.B(n_1225),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1273),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1228),
.B(n_1292),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1234),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1228),
.B(n_1292),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1293),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1236),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1294),
.B(n_1226),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1329),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1241),
.B(n_1298),
.Y(n_1366)
);

CKINVDCx12_ASAP7_75t_R g1367 ( 
.A(n_1240),
.Y(n_1367)
);

BUFx2_ASAP7_75t_SL g1368 ( 
.A(n_1274),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_R g1369 ( 
.A(n_1312),
.B(n_1326),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1294),
.B(n_1226),
.Y(n_1370)
);

INVxp33_ASAP7_75t_L g1371 ( 
.A(n_1229),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1310),
.B(n_1311),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1257),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1266),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1253),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1338),
.B(n_1277),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1284),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1252),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1287),
.A2(n_1286),
.B(n_1289),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1227),
.A2(n_1324),
.A3(n_1317),
.B(n_1332),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1252),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1250),
.B(n_1328),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1287),
.A2(n_1286),
.B(n_1289),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1271),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1230),
.A2(n_1309),
.B(n_1232),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1311),
.B(n_1334),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1265),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1243),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1244),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1335),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1255),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1328),
.B(n_1336),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1302),
.B(n_1268),
.Y(n_1393)
);

AOI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1303),
.A2(n_1304),
.B(n_1263),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1281),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1281),
.Y(n_1396)
);

AO21x2_ASAP7_75t_L g1397 ( 
.A1(n_1298),
.A2(n_1330),
.B(n_1299),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1302),
.B(n_1237),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1232),
.B(n_1246),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1276),
.A2(n_1251),
.B(n_1258),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1299),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1264),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1330),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1241),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1239),
.A2(n_1248),
.B(n_1323),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1297),
.A2(n_1301),
.B(n_1333),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1269),
.A2(n_1301),
.B(n_1297),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1262),
.A2(n_1337),
.B(n_1316),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1325),
.B(n_1333),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1269),
.Y(n_1410)
);

CKINVDCx16_ASAP7_75t_R g1411 ( 
.A(n_1247),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1260),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1340),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1235),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1248),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1348),
.B(n_1325),
.Y(n_1416)
);

AND2x4_ASAP7_75t_SL g1417 ( 
.A(n_1355),
.B(n_1315),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1384),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1410),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1348),
.B(n_1331),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1385),
.A2(n_1331),
.B(n_1305),
.C(n_1231),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1348),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1410),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1346),
.B(n_1318),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1379),
.A2(n_1235),
.B(n_1305),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1373),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1406),
.A2(n_1235),
.B1(n_1238),
.B2(n_1320),
.Y(n_1427)
);

AOI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1343),
.A2(n_1307),
.B1(n_1245),
.B2(n_1320),
.C(n_1314),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1394),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1379),
.A2(n_1242),
.B(n_1306),
.Y(n_1430)
);

NAND3xp33_ASAP7_75t_L g1431 ( 
.A(n_1385),
.B(n_1256),
.C(n_1306),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1352),
.B(n_1314),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1348),
.B(n_1315),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1356),
.B(n_1259),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1347),
.B(n_1395),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1356),
.B(n_1307),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1365),
.B(n_1261),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_SL g1438 ( 
.A(n_1368),
.B(n_1300),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1362),
.B(n_1244),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1392),
.B(n_1249),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1368),
.B(n_1313),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1345),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1347),
.B(n_1319),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1343),
.A2(n_1339),
.B1(n_1406),
.B2(n_1366),
.C(n_1388),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1392),
.B(n_1390),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1386),
.B(n_1372),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1345),
.Y(n_1447)
);

AO32x2_ASAP7_75t_L g1448 ( 
.A1(n_1414),
.A2(n_1397),
.A3(n_1404),
.B1(n_1345),
.B2(n_1366),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1355),
.B(n_1396),
.Y(n_1449)
);

OAI211xp5_ASAP7_75t_L g1450 ( 
.A1(n_1409),
.A2(n_1388),
.B(n_1374),
.C(n_1404),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1351),
.B(n_1353),
.Y(n_1451)
);

AOI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1409),
.A2(n_1364),
.B1(n_1370),
.B2(n_1382),
.C(n_1391),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1374),
.A2(n_1382),
.B1(n_1370),
.B2(n_1364),
.Y(n_1453)
);

AOI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1391),
.A2(n_1403),
.B1(n_1401),
.B2(n_1361),
.C(n_1359),
.Y(n_1454)
);

BUFx4f_ASAP7_75t_SL g1455 ( 
.A(n_1413),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1396),
.B(n_1354),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1371),
.B(n_1367),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1407),
.A2(n_1398),
.B1(n_1361),
.B2(n_1359),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1354),
.B(n_1355),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1402),
.B(n_1380),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1355),
.B(n_1342),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1357),
.A2(n_1380),
.B(n_1401),
.C(n_1403),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1342),
.B(n_1395),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1357),
.A2(n_1380),
.B(n_1375),
.C(n_1399),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1377),
.A2(n_1414),
.B1(n_1402),
.B2(n_1398),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1377),
.A2(n_1414),
.B1(n_1398),
.B2(n_1408),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1379),
.A2(n_1383),
.B(n_1400),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1342),
.B(n_1360),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1400),
.A2(n_1375),
.B(n_1376),
.Y(n_1469)
);

AND2x2_ASAP7_75t_SL g1470 ( 
.A(n_1393),
.B(n_1399),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1367),
.B(n_1411),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1342),
.B(n_1363),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1384),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1394),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1342),
.B(n_1363),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1444),
.A2(n_1407),
.B1(n_1397),
.B2(n_1398),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1460),
.B(n_1342),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1450),
.A2(n_1407),
.B1(n_1397),
.B2(n_1380),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1448),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1461),
.B(n_1383),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1461),
.B(n_1383),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1427),
.B(n_1407),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1463),
.B(n_1435),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1426),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1467),
.B(n_1344),
.Y(n_1485)
);

NOR2xp67_ASAP7_75t_L g1486 ( 
.A(n_1429),
.B(n_1358),
.Y(n_1486)
);

INVx3_ASAP7_75t_SL g1487 ( 
.A(n_1442),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1467),
.B(n_1468),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1458),
.A2(n_1378),
.B1(n_1381),
.B2(n_1384),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1418),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1474),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1462),
.B(n_1350),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1468),
.B(n_1344),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1472),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1475),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1445),
.B(n_1349),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1440),
.B(n_1387),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1422),
.B(n_1376),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1419),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1423),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1448),
.B(n_1350),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1448),
.B(n_1341),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1451),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1485),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1484),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1484),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1485),
.Y(n_1508)
);

OAI33xp33_ASAP7_75t_L g1509 ( 
.A1(n_1489),
.A2(n_1453),
.A3(n_1466),
.B1(n_1465),
.B2(n_1424),
.B3(n_1443),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1448),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1481),
.B(n_1430),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1481),
.B(n_1430),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1478),
.B(n_1421),
.C(n_1452),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1482),
.A2(n_1434),
.B1(n_1397),
.B2(n_1431),
.Y(n_1515)
);

AOI322xp5_ASAP7_75t_L g1516 ( 
.A1(n_1489),
.A2(n_1454),
.A3(n_1421),
.B1(n_1464),
.B2(n_1434),
.C1(n_1462),
.C2(n_1446),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1497),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1498),
.B(n_1425),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1488),
.B(n_1470),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1479),
.B(n_1464),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1488),
.B(n_1470),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1491),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1479),
.A2(n_1469),
.B(n_1425),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_SL g1524 ( 
.A(n_1478),
.B(n_1428),
.C(n_1443),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1491),
.Y(n_1525)
);

AND3x1_ASAP7_75t_L g1526 ( 
.A(n_1476),
.B(n_1471),
.C(n_1441),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1479),
.B(n_1449),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1483),
.B(n_1456),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1482),
.A2(n_1378),
.B1(n_1381),
.B2(n_1456),
.C(n_1416),
.Y(n_1529)
);

AOI222xp33_ASAP7_75t_L g1530 ( 
.A1(n_1492),
.A2(n_1455),
.B1(n_1457),
.B2(n_1420),
.C1(n_1416),
.C2(n_1438),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1488),
.B(n_1459),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1495),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1476),
.A2(n_1432),
.B1(n_1437),
.B2(n_1436),
.C(n_1408),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_SL g1534 ( 
.A(n_1492),
.B(n_1376),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1493),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1522),
.B(n_1494),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1506),
.B(n_1502),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1522),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1502),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1505),
.Y(n_1541)
);

AND2x2_ASAP7_75t_SL g1542 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1526),
.B(n_1418),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1527),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1525),
.B(n_1494),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1525),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1535),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1507),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1528),
.B(n_1501),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1535),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1510),
.B(n_1503),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1532),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1507),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1528),
.B(n_1501),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1532),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1520),
.B(n_1510),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1514),
.A2(n_1420),
.B1(n_1436),
.B2(n_1497),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1519),
.B(n_1503),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1504),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1519),
.B(n_1501),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1520),
.B(n_1483),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1519),
.B(n_1493),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1504),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1518),
.B(n_1498),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1520),
.B(n_1500),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1532),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1521),
.B(n_1511),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1521),
.B(n_1511),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1538),
.Y(n_1569)
);

NOR2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1556),
.B(n_1524),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1543),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1542),
.B(n_1521),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1561),
.B(n_1527),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1544),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1542),
.B(n_1531),
.Y(n_1575)
);

AOI211xp5_ASAP7_75t_L g1576 ( 
.A1(n_1543),
.A2(n_1533),
.B(n_1514),
.C(n_1524),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1561),
.B(n_1565),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1538),
.Y(n_1578)
);

OAI32xp33_ASAP7_75t_L g1579 ( 
.A1(n_1556),
.A2(n_1533),
.A3(n_1517),
.B1(n_1527),
.B2(n_1477),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1546),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1551),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

NOR3x1_ASAP7_75t_L g1583 ( 
.A(n_1565),
.B(n_1499),
.C(n_1509),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1557),
.B(n_1529),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1536),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1542),
.B(n_1531),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1557),
.B(n_1529),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1542),
.B(n_1516),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1551),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1567),
.B(n_1531),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1516),
.Y(n_1591)
);

NAND2x1p5_ASAP7_75t_L g1592 ( 
.A(n_1564),
.B(n_1523),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1536),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1562),
.B(n_1515),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1544),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1564),
.A2(n_1515),
.B1(n_1509),
.B2(n_1530),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1545),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1551),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1568),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1567),
.B(n_1518),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1564),
.B(n_1411),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1549),
.B(n_1504),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1545),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1547),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1549),
.B(n_1504),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1547),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1550),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1568),
.B(n_1511),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1550),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1570),
.B(n_1562),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1569),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1599),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1569),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1588),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1578),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1591),
.B(n_1562),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1604),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1574),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1572),
.B(n_1568),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1604),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1576),
.A2(n_1530),
.B1(n_1518),
.B2(n_1512),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1580),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1574),
.B(n_1560),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1582),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1599),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1572),
.B(n_1575),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1575),
.B(n_1560),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1595),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1595),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1590),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1584),
.B(n_1558),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1606),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1587),
.B(n_1558),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1573),
.B(n_1593),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1583),
.B(n_1558),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1590),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1596),
.A2(n_1601),
.B1(n_1571),
.B2(n_1594),
.Y(n_1641)
);

AND3x2_ASAP7_75t_L g1642 ( 
.A(n_1586),
.B(n_1439),
.C(n_1600),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1597),
.B(n_1559),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1607),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1607),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1620),
.Y(n_1646)
);

XNOR2xp5_ASAP7_75t_L g1647 ( 
.A(n_1641),
.B(n_1618),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_1586),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1628),
.A2(n_1523),
.B1(n_1600),
.B2(n_1518),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1628),
.A2(n_1523),
.B1(n_1600),
.B2(n_1518),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1612),
.B(n_1581),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1620),
.B(n_1439),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1634),
.A2(n_1579),
.B(n_1517),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1637),
.B(n_1581),
.Y(n_1654)
);

AOI211xp5_ASAP7_75t_L g1655 ( 
.A1(n_1639),
.A2(n_1579),
.B(n_1473),
.C(n_1418),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1623),
.A2(n_1512),
.B(n_1513),
.C(n_1585),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1631),
.A2(n_1523),
.B1(n_1592),
.B2(n_1609),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1621),
.B(n_1585),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1630),
.A2(n_1534),
.B(n_1603),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1621),
.A2(n_1603),
.B1(n_1610),
.B2(n_1609),
.C(n_1589),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1630),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1625),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1613),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1629),
.B(n_1564),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1642),
.A2(n_1523),
.B1(n_1513),
.B2(n_1512),
.Y(n_1665)
);

AOI222xp33_ASAP7_75t_L g1666 ( 
.A1(n_1629),
.A2(n_1534),
.B1(n_1589),
.B2(n_1598),
.C1(n_1513),
.C2(n_1537),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1617),
.B(n_1598),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1613),
.Y(n_1668)
);

OAI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1614),
.A2(n_1592),
.B(n_1602),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1619),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_1389),
.Y(n_1671)
);

AOI222xp33_ASAP7_75t_L g1672 ( 
.A1(n_1656),
.A2(n_1614),
.B1(n_1627),
.B2(n_1640),
.C1(n_1632),
.C2(n_1626),
.Y(n_1672)
);

BUFx2_ASAP7_75t_SL g1673 ( 
.A(n_1646),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1646),
.B(n_1627),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1662),
.Y(n_1675)
);

NOR4xp25_ASAP7_75t_SL g1676 ( 
.A(n_1669),
.B(n_1660),
.C(n_1668),
.D(n_1670),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1661),
.B(n_1632),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1663),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1652),
.B(n_1640),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1648),
.B(n_1638),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1667),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1654),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1651),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1658),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1652),
.B(n_1625),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1664),
.Y(n_1686)
);

OAI21xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1666),
.A2(n_1633),
.B(n_1638),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1653),
.B(n_1624),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1655),
.A2(n_1635),
.B(n_1615),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1673),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1671),
.B(n_1659),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_SL g1692 ( 
.A(n_1671),
.B(n_1657),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1674),
.Y(n_1693)
);

OAI32xp33_ASAP7_75t_L g1694 ( 
.A1(n_1687),
.A2(n_1688),
.A3(n_1676),
.B1(n_1680),
.B2(n_1675),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1674),
.B(n_1688),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1686),
.B(n_1633),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1689),
.A2(n_1665),
.B(n_1650),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1680),
.A2(n_1645),
.B1(n_1636),
.B2(n_1644),
.Y(n_1698)
);

OAI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1683),
.A2(n_1649),
.B1(n_1677),
.B2(n_1682),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1684),
.A2(n_1644),
.B1(n_1622),
.B2(n_1619),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1685),
.Y(n_1701)
);

XNOR2xp5_ASAP7_75t_L g1702 ( 
.A(n_1690),
.B(n_1679),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1701),
.B(n_1681),
.Y(n_1703)
);

NAND4xp25_ASAP7_75t_L g1704 ( 
.A(n_1691),
.B(n_1672),
.C(n_1678),
.D(n_1685),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1695),
.A2(n_1611),
.B1(n_1592),
.B2(n_1622),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1693),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1699),
.A2(n_1611),
.B1(n_1523),
.B2(n_1418),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1696),
.B(n_1537),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1700),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1692),
.B(n_1697),
.Y(n_1710)
);

AOI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1694),
.B(n_1698),
.C(n_1369),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1706),
.Y(n_1712)
);

OAI321xp33_ASAP7_75t_L g1713 ( 
.A1(n_1707),
.A2(n_1704),
.A3(n_1709),
.B1(n_1705),
.B2(n_1703),
.C(n_1698),
.Y(n_1713)
);

OAI211xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1707),
.A2(n_1700),
.B(n_1643),
.C(n_1608),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1702),
.A2(n_1643),
.B1(n_1608),
.B2(n_1605),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1712),
.Y(n_1716)
);

AOI211xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1713),
.A2(n_1708),
.B(n_1377),
.C(n_1439),
.Y(n_1717)
);

NOR4xp75_ASAP7_75t_L g1718 ( 
.A(n_1715),
.B(n_1377),
.C(n_1405),
.D(n_1537),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_SL g1719 ( 
.A(n_1711),
.B(n_1714),
.C(n_1345),
.Y(n_1719)
);

AOI211xp5_ASAP7_75t_SL g1720 ( 
.A1(n_1713),
.A2(n_1605),
.B(n_1602),
.C(n_1412),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1711),
.A2(n_1473),
.B1(n_1564),
.B2(n_1490),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1716),
.Y(n_1722)
);

XNOR2xp5_ASAP7_75t_L g1723 ( 
.A(n_1721),
.B(n_1417),
.Y(n_1723)
);

BUFx12f_ASAP7_75t_L g1724 ( 
.A(n_1717),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1719),
.Y(n_1725)
);

NAND4xp75_ASAP7_75t_L g1726 ( 
.A(n_1720),
.B(n_1540),
.C(n_1433),
.D(n_1486),
.Y(n_1726)
);

AOI31xp33_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1718),
.A3(n_1387),
.B(n_1415),
.Y(n_1727)
);

OR3x2_ASAP7_75t_L g1728 ( 
.A(n_1722),
.B(n_1412),
.C(n_1496),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1723),
.A2(n_1473),
.B1(n_1563),
.B2(n_1559),
.C(n_1405),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1728),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1730),
.Y(n_1731)
);

OA22x2_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1724),
.B1(n_1727),
.B2(n_1726),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1724),
.B1(n_1729),
.B2(n_1559),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1473),
.B1(n_1563),
.B2(n_1559),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1734),
.A2(n_1563),
.B1(n_1447),
.B2(n_1442),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1734),
.A2(n_1563),
.B(n_1566),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1735),
.B(n_1736),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1735),
.B(n_1552),
.Y(n_1738)
);

OAI31xp33_ASAP7_75t_L g1739 ( 
.A1(n_1737),
.A2(n_1738),
.A3(n_1566),
.B(n_1555),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1539),
.B1(n_1553),
.B2(n_1541),
.C(n_1548),
.Y(n_1740)
);

AOI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1487),
.B(n_1415),
.C(n_1555),
.Y(n_1741)
);


endmodule