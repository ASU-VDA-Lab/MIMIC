module fake_netlist_6_4765_n_90 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_90);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_90;

wire n_52;
wire n_46;
wire n_88;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_86;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_16),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_4),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_22),
.B(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_12),
.B(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_5),
.B(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_1),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_23),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_32),
.B(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_36),
.B1(n_34),
.B2(n_30),
.Y(n_50)
);

OAI21x1_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_32),
.B(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_24),
.B(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_38),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_42),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx2_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_55),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_50),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

AOI221xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_29),
.B1(n_33),
.B2(n_48),
.C(n_57),
.Y(n_71)
);

NOR2x1_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_68),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND4xp25_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_65),
.C(n_68),
.D(n_34),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_36),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_83),
.Y(n_84)
);

NAND4xp75_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_76),
.C(n_38),
.D(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_81),
.B1(n_82),
.B2(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_33),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_86),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_63),
.Y(n_90)
);


endmodule