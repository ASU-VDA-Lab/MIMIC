module fake_jpeg_30172_n_150 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_32),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_79),
.Y(n_85)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_58),
.C(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_3),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_89),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_60),
.B1(n_59),
.B2(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_88),
.B1(n_65),
.B2(n_55),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_60),
.B1(n_69),
.B2(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_95),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_62),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_85),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_65),
.B1(n_55),
.B2(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_101),
.B1(n_107),
.B2(n_8),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_70),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_71),
.B1(n_67),
.B2(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_4),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_7),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_5),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_46),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_122),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_105),
.B1(n_94),
.B2(n_109),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_121)
);

BUFx12f_ASAP7_75t_SL g122 ( 
.A(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_29),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_22),
.B(n_27),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_117),
.B(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_48),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_33),
.A3(n_35),
.B1(n_37),
.B2(n_41),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_135),
.B1(n_110),
.B2(n_119),
.C(n_47),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_43),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_140),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_139),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_130),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_126),
.B(n_142),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_130),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_127),
.B(n_137),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_145),
.Y(n_150)
);


endmodule