module fake_jpeg_11715_n_428 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_428);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_428;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_3),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_53),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_70),
.Y(n_103)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_63),
.Y(n_115)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_21),
.B(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_15),
.B(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_84),
.Y(n_107)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_15),
.B(n_11),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_18),
.Y(n_96)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_96),
.B(n_25),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_47),
.A2(n_23),
.B1(n_24),
.B2(n_16),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_85),
.B1(n_64),
.B2(n_77),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_46),
.A2(n_32),
.B1(n_17),
.B2(n_24),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_111),
.A2(n_126),
.B1(n_32),
.B2(n_75),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g118 ( 
.A(n_72),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_118),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_122),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_42),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_43),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_56),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_33),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_23),
.B1(n_61),
.B2(n_66),
.Y(n_151)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_99),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_147),
.B(n_166),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_205)
);

CKINVDCx12_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_33),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_153),
.B(n_183),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_186),
.B1(n_124),
.B2(n_139),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_163),
.B1(n_176),
.B2(n_181),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

CKINVDCx12_ASAP7_75t_R g158 ( 
.A(n_115),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_160),
.Y(n_220)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_83),
.B1(n_81),
.B2(n_78),
.Y(n_163)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_105),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_26),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_106),
.B(n_116),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_98),
.A2(n_67),
.B1(n_59),
.B2(n_58),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_172),
.A2(n_139),
.B1(n_135),
.B2(n_110),
.Y(n_222)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_103),
.A2(n_19),
.B1(n_25),
.B2(n_17),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_40),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_184),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_179),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_182),
.Y(n_196)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_19),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_101),
.B(n_40),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_18),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_187),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_111),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_10),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_102),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_126),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_126),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_8),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_106),
.C(n_133),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_195),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_128),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_210),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_0),
.B(n_4),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_208),
.A2(n_171),
.B(n_161),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_121),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_123),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_229),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_167),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_223),
.B1(n_165),
.B2(n_181),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_172),
.A2(n_133),
.B1(n_141),
.B2(n_135),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_164),
.B(n_124),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_138),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_154),
.A2(n_138),
.B1(n_123),
.B2(n_92),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_160),
.B1(n_169),
.B2(n_150),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_232),
.B(n_192),
.Y(n_293)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_148),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_241),
.Y(n_272)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_238),
.B(n_242),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_200),
.A2(n_145),
.B1(n_149),
.B2(n_162),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_221),
.B(n_222),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_244),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_156),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_204),
.Y(n_242)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_186),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_196),
.B(n_186),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_245),
.B(n_251),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_252),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_229),
.B1(n_205),
.B2(n_193),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_249),
.B1(n_253),
.B2(n_220),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_205),
.A2(n_186),
.B1(n_141),
.B2(n_92),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_210),
.B(n_195),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_175),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_159),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_257),
.Y(n_285)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_261),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_170),
.Y(n_257)
);

NOR2x1_ASAP7_75t_R g274 ( 
.A(n_258),
.B(n_208),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_260),
.Y(n_290)
);

AND2x6_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_119),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_263),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_193),
.B(n_173),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_195),
.B(n_0),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_6),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_277),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_210),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_269),
.B(n_241),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_219),
.B(n_212),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_271),
.B(n_245),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_193),
.B(n_194),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_274),
.B(n_264),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_276),
.A2(n_233),
.B1(n_247),
.B2(n_263),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_295),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_235),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_283),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_248),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_231),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_286),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_231),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_213),
.C(n_202),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_294),
.C(n_256),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_249),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_246),
.B(n_213),
.C(n_194),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_248),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_310),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_316),
.C(n_293),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_309),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_248),
.B(n_244),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_266),
.B(n_259),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_302),
.B(n_282),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_274),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_321),
.B1(n_270),
.B2(n_278),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_261),
.Y(n_307)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_267),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_277),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_312),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_262),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_285),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_314),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_269),
.B(n_240),
.C(n_251),
.Y(n_316)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_322),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_318),
.A2(n_319),
.B(n_287),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_271),
.A2(n_265),
.B(n_275),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_276),
.A2(n_260),
.B1(n_253),
.B2(n_243),
.Y(n_321)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_301),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_325),
.B(n_305),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_300),
.B(n_290),
.Y(n_326)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_291),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_333),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_341),
.C(n_344),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_287),
.B(n_295),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_330),
.A2(n_322),
.B(n_317),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_302),
.B(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_337),
.A2(n_297),
.B1(n_278),
.B2(n_268),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_296),
.A2(n_308),
.B1(n_320),
.B2(n_304),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_340),
.A2(n_309),
.B1(n_312),
.B2(n_315),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_289),
.C(n_272),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_300),
.B(n_272),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_303),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_255),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_345),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_275),
.C(n_282),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_320),
.B(n_280),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_307),
.Y(n_347)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_361),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_328),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_366),
.Y(n_370)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_336),
.A2(n_321),
.B1(n_316),
.B2(n_319),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_355),
.A2(n_365),
.B(n_336),
.Y(n_367)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_356),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_358),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_299),
.C(n_303),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_364),
.C(n_325),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_362),
.A2(n_330),
.B1(n_332),
.B2(n_331),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_299),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_335),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_297),
.C(n_305),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_324),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_369),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_355),
.A2(n_326),
.B(n_344),
.Y(n_368)
);

AO221x1_ASAP7_75t_L g389 ( 
.A1(n_368),
.A2(n_365),
.B1(n_357),
.B2(n_364),
.C(n_361),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_352),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_360),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_335),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_377),
.C(n_380),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_379),
.A2(n_382),
.B1(n_354),
.B2(n_358),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_338),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_353),
.A2(n_332),
.B1(n_331),
.B2(n_324),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_388),
.Y(n_396)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_376),
.A2(n_323),
.A3(n_334),
.B1(n_342),
.B2(n_346),
.C1(n_356),
.C2(n_337),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_387),
.A2(n_393),
.B1(n_371),
.B2(n_220),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_357),
.C(n_359),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_389),
.A2(n_390),
.B1(n_392),
.B2(n_394),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_349),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_370),
.A2(n_347),
.B(n_339),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_374),
.Y(n_395)
);

OAI321xp33_ASAP7_75t_L g392 ( 
.A1(n_372),
.A2(n_339),
.A3(n_322),
.B1(n_317),
.B2(n_288),
.C(n_279),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g393 ( 
.A(n_367),
.B(n_288),
.CI(n_279),
.CON(n_393),
.SN(n_393)
);

NOR3xp33_ASAP7_75t_SL g394 ( 
.A(n_381),
.B(n_374),
.C(n_369),
.Y(n_394)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_378),
.C(n_380),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_401),
.Y(n_405)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_400),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_378),
.C(n_371),
.Y(n_401)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_402),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_215),
.C(n_217),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_404),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_385),
.A2(n_216),
.B1(n_215),
.B2(n_221),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_399),
.B(n_384),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_406),
.A2(n_398),
.B(n_403),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_396),
.A2(n_391),
.B1(n_393),
.B2(n_394),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_412),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_393),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_397),
.C(n_401),
.Y(n_413)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_413),
.Y(n_420)
);

NOR2x1_ASAP7_75t_SL g418 ( 
.A(n_415),
.B(n_416),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_395),
.C(n_216),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_179),
.Y(n_417)
);

AOI322xp5_ASAP7_75t_L g419 ( 
.A1(n_417),
.A2(n_178),
.A3(n_409),
.B1(n_179),
.B2(n_410),
.C1(n_407),
.C2(n_157),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_419),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_420),
.A2(n_414),
.B(n_411),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_421),
.B(n_418),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_422),
.Y(n_424)
);

MAJx2_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_178),
.C(n_114),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_8),
.C(n_6),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_7),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_7),
.Y(n_428)
);


endmodule