module fake_jpeg_12411_n_390 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_0),
.B(n_2),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_43),
.B(n_64),
.C(n_4),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_44),
.B(n_48),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_13),
.B(n_12),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_61),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_68),
.Y(n_115)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_11),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_16),
.B(n_3),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_76),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_3),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_82),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_4),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_22),
.B1(n_34),
.B2(n_41),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_96),
.B1(n_129),
.B2(n_59),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_15),
.B1(n_34),
.B2(n_28),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_86),
.A2(n_90),
.B(n_103),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_22),
.B1(n_28),
.B2(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_87),
.A2(n_100),
.B1(n_102),
.B2(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_69),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_15),
.B1(n_37),
.B2(n_35),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_71),
.B1(n_15),
.B2(n_45),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_40),
.B1(n_32),
.B2(n_27),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_38),
.B1(n_33),
.B2(n_40),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_110),
.B1(n_123),
.B2(n_130),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_32),
.B1(n_27),
.B2(n_38),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_56),
.A2(n_37),
.B1(n_35),
.B2(n_23),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_82),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_65),
.A2(n_23),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_23),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_4),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_133),
.B(n_152),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_143),
.Y(n_181)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_66),
.B1(n_80),
.B2(n_77),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_180),
.B1(n_93),
.B2(n_132),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_141),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_139),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_148),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_78),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_142),
.B(n_149),
.C(n_164),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_74),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_116),
.Y(n_144)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_146),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_128),
.B1(n_126),
.B2(n_84),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_157),
.B(n_159),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_101),
.B(n_67),
.Y(n_149)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_82),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_63),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_53),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_172),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_111),
.A2(n_82),
.B1(n_73),
.B2(n_57),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_118),
.B(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_169),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_73),
.B(n_54),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_162),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_87),
.A2(n_73),
.B(n_61),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_163),
.A2(n_171),
.B(n_177),
.C(n_170),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_7),
.B(n_8),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_119),
.A2(n_75),
.B1(n_9),
.B2(n_10),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_89),
.B1(n_121),
.B2(n_127),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_112),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_107),
.C(n_106),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_7),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_170),
.B(n_177),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_122),
.B(n_107),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_9),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_10),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_98),
.B(n_117),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_91),
.B(n_10),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_117),
.B(n_49),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_89),
.A2(n_49),
.B1(n_121),
.B2(n_127),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_183),
.A2(n_167),
.B1(n_144),
.B2(n_176),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_93),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_184),
.B(n_213),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_186),
.A2(n_191),
.B1(n_195),
.B2(n_220),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_133),
.A2(n_132),
.B1(n_153),
.B2(n_173),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_135),
.B1(n_171),
.B2(n_134),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_197),
.B(n_201),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_159),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_198),
.A2(n_219),
.B(n_208),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_152),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_137),
.A2(n_152),
.B1(n_172),
.B2(n_174),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_214),
.B1(n_182),
.B2(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_142),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_161),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_136),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_160),
.B1(n_139),
.B2(n_163),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_175),
.B1(n_139),
.B2(n_179),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_168),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_176),
.C(n_167),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_226),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_151),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_224),
.B(n_234),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_144),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_237),
.B1(n_255),
.B2(n_194),
.Y(n_266)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_232),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_167),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_176),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_206),
.B1(n_209),
.B2(n_207),
.Y(n_264)
);

XNOR2x2_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_216),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_244),
.B(n_251),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_195),
.B1(n_208),
.B2(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_239),
.B(n_246),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_252),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_254),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_201),
.B(n_193),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_238),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_198),
.B(n_183),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_200),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_205),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_205),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_203),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_254),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_190),
.B(n_199),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_186),
.A2(n_184),
.B1(n_206),
.B2(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_258),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_264),
.A2(n_276),
.B1(n_283),
.B2(n_284),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_237),
.A2(n_194),
.B1(n_207),
.B2(n_196),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_266),
.B1(n_272),
.B2(n_244),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_196),
.B(n_217),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_267),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_217),
.C(n_218),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_273),
.C(n_253),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_233),
.A2(n_194),
.B1(n_217),
.B2(n_188),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_188),
.B1(n_218),
.B2(n_235),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_224),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_242),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_223),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_233),
.A2(n_218),
.B1(n_255),
.B2(n_225),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_240),
.B1(n_226),
.B2(n_232),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_236),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_261),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_291),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_234),
.Y(n_290)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

BUFx12_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_294),
.A2(n_305),
.B1(n_262),
.B2(n_271),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

BUFx12_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_298),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_261),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_243),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_311),
.C(n_312),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_263),
.Y(n_300)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_227),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_288),
.C(n_274),
.Y(n_315)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_288),
.A2(n_245),
.B(n_231),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_309),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_259),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_236),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_238),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_229),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_265),
.B1(n_272),
.B2(n_287),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_314),
.A2(n_325),
.B1(n_302),
.B2(n_269),
.Y(n_349)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_284),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_326),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_276),
.B1(n_274),
.B2(n_259),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_324),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_322),
.B(n_230),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_303),
.A2(n_268),
.B1(n_280),
.B2(n_262),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_260),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_260),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_297),
.C(n_311),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_350),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_335),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_338),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_328),
.B(n_301),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_256),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_346),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_290),
.C(n_303),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_343),
.C(n_344),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_290),
.C(n_313),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_313),
.C(n_306),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_316),
.A2(n_302),
.B(n_271),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_332),
.B(n_269),
.Y(n_347)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_347),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_325),
.Y(n_348)
);

INVx11_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_321),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_340),
.A2(n_316),
.B(n_333),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_354),
.B(n_358),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_345),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_326),
.C(n_329),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_340),
.A2(n_314),
.B1(n_317),
.B2(n_315),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_361),
.A2(n_336),
.B1(n_346),
.B2(n_344),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_322),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_334),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_357),
.B(n_341),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_366),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_342),
.C(n_337),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_368),
.C(n_369),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_350),
.C(n_320),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_363),
.B(n_327),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g378 ( 
.A1(n_370),
.A2(n_356),
.B(n_358),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_361),
.A2(n_295),
.B1(n_279),
.B2(n_248),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_372),
.A2(n_354),
.B(n_355),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_369),
.A2(n_362),
.B1(n_353),
.B2(n_355),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_375),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_367),
.A2(n_362),
.B1(n_353),
.B2(n_351),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_376),
.A2(n_378),
.B(n_379),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_377),
.A2(n_371),
.B(n_360),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_380),
.B(n_381),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_377),
.Y(n_382)
);

AOI322xp5_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_291),
.A3(n_296),
.B1(n_351),
.B2(n_360),
.C1(n_370),
.C2(n_359),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_385),
.B(n_383),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_386),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_359),
.C(n_279),
.Y(n_387)
);

O2A1O1Ixp33_ASAP7_75t_SL g389 ( 
.A1(n_388),
.A2(n_387),
.B(n_291),
.C(n_296),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_257),
.Y(n_390)
);


endmodule