module fake_jpeg_13133_n_101 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_0),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_34),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_39),
.B1(n_31),
.B2(n_37),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_29),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_39),
.B1(n_31),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_58),
.B1(n_50),
.B2(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_1),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_68),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_70),
.B(n_19),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_1),
.C(n_2),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_69),
.C(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_5),
.B(n_8),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_10),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_9),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_12),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_83),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_21),
.C(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_20),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_23),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_89),
.B1(n_91),
.B2(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_79),
.B1(n_76),
.B2(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_76),
.B1(n_88),
.B2(n_61),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_78),
.B(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_96),
.B(n_95),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_26),
.Y(n_101)
);


endmodule