module fake_jpeg_10390_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_51),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_28),
.B1(n_20),
.B2(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_53),
.B1(n_33),
.B2(n_26),
.Y(n_93)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_65),
.Y(n_82)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_20),
.B1(n_28),
.B2(n_22),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_18),
.B1(n_25),
.B2(n_33),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_20),
.B1(n_23),
.B2(n_31),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_18),
.B(n_25),
.Y(n_107)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_92),
.Y(n_125)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_31),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_91),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_37),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_89),
.B1(n_50),
.B2(n_101),
.Y(n_131)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_96),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_39),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_26),
.B(n_33),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_27),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_102),
.B1(n_61),
.B2(n_49),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_46),
.B1(n_27),
.B2(n_31),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_54),
.B(n_30),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_86),
.Y(n_122)
);

NAND2x1_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_88),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_107),
.B(n_124),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_115),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_120),
.B1(n_97),
.B2(n_89),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_98),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_81),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_76),
.C(n_72),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_85),
.C(n_36),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_85),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_77),
.A2(n_76),
.B1(n_70),
.B2(n_99),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_14),
.C(n_13),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_10),
.Y(n_156)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_50),
.A3(n_61),
.B1(n_49),
.B2(n_36),
.Y(n_124)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_78),
.B1(n_94),
.B2(n_90),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_30),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_50),
.B1(n_100),
.B2(n_78),
.Y(n_141)
);

XOR2x1_ASAP7_75t_L g197 ( 
.A(n_133),
.B(n_29),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_136),
.B(n_142),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_138),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_115),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_110),
.C(n_29),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_116),
.B1(n_117),
.B2(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_148),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_79),
.B1(n_71),
.B2(n_92),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_64),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_32),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_152),
.B(n_159),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_32),
.B1(n_19),
.B2(n_34),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_32),
.B1(n_19),
.B2(n_34),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_32),
.B1(n_34),
.B2(n_44),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_44),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_24),
.B1(n_17),
.B2(n_29),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_117),
.B(n_114),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_74),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_104),
.B(n_0),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_74),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_181),
.C(n_183),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_113),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_187),
.Y(n_203)
);

OAI22x1_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_151),
.B1(n_133),
.B2(n_162),
.Y(n_213)
);

XOR2x2_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_116),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_175),
.B(n_197),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_147),
.A2(n_126),
.B1(n_109),
.B2(n_127),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_195),
.B1(n_159),
.B2(n_150),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_182),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_199),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_111),
.C(n_122),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_111),
.A3(n_130),
.B1(n_24),
.B2(n_17),
.Y(n_188)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_109),
.B1(n_74),
.B2(n_24),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_154),
.B1(n_153),
.B2(n_136),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_141),
.A2(n_17),
.B1(n_29),
.B2(n_11),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_201),
.A2(n_205),
.B1(n_212),
.B2(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_209),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_206),
.B(n_214),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_145),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_216),
.C(n_219),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_144),
.B1(n_157),
.B2(n_148),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_224),
.B1(n_172),
.B2(n_191),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_178),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_134),
.B1(n_142),
.B2(n_133),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_178),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_134),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_162),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_194),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_227),
.C(n_189),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_135),
.B1(n_129),
.B2(n_123),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_172),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_225),
.B(n_228),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_135),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_174),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_241),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_213),
.A2(n_190),
.B1(n_189),
.B2(n_175),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_234),
.B1(n_245),
.B2(n_249),
.Y(n_261)
);

BUFx4f_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_190),
.B1(n_229),
.B2(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_244),
.C(n_252),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_187),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_251),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_185),
.CI(n_188),
.CON(n_241),
.SN(n_241)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_253),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_185),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_208),
.A2(n_166),
.B1(n_177),
.B2(n_192),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_177),
.B1(n_168),
.B2(n_139),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_220),
.B(n_203),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_29),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_223),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_129),
.B1(n_123),
.B2(n_29),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_216),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_207),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_262),
.C(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_210),
.B1(n_226),
.B2(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_226),
.B(n_203),
.C(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_242),
.A2(n_231),
.B(n_235),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_260),
.A2(n_241),
.B(n_233),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_14),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_14),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_13),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_247),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_12),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.C(n_275),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_11),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_243),
.A2(n_12),
.B1(n_1),
.B2(n_3),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_254),
.B1(n_234),
.B2(n_249),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_12),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_277),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_281),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_252),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_288),
.C(n_291),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_290),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_233),
.C(n_1),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_0),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_273),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_270),
.B1(n_260),
.B2(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_261),
.B1(n_265),
.B2(n_267),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_280),
.B1(n_290),
.B2(n_278),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_271),
.B1(n_275),
.B2(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_288),
.C(n_282),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_280),
.B(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_279),
.A2(n_256),
.B1(n_4),
.B2(n_5),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_3),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_6),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_3),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_4),
.B(n_5),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_293),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_297),
.C(n_299),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_301),
.B(n_304),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_295),
.B(n_297),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_4),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_314),
.B(n_310),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_6),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_317),
.B(n_7),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_7),
.B(n_8),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_325),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_324),
.B(n_314),
.C(n_316),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_323),
.B(n_293),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_298),
.C(n_294),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_296),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_318),
.B1(n_309),
.B2(n_298),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_332),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_330),
.B(n_322),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_334),
.A2(n_335),
.B(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_336),
.B(n_323),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_328),
.Y(n_340)
);

OAI321xp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_8),
.A3(n_9),
.B1(n_327),
.B2(n_321),
.C(n_335),
.Y(n_341)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_8),
.CI(n_9),
.CON(n_342),
.SN(n_342)
);


endmodule