module real_aes_1270_n_14 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_14);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_14;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_34;
wire n_19;
wire n_40;
wire n_25;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_0), .Y(n_24) );
NOR3xp33_ASAP7_75t_SL g22 ( .A(n_1), .B(n_4), .C(n_23), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_2), .Y(n_23) );
NAND3xp33_ASAP7_75t_SL g26 ( .A(n_3), .B(n_27), .C(n_28), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_5), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_7), .Y(n_27) );
NAND2xp33_ASAP7_75t_SL g16 ( .A(n_8), .B(n_17), .Y(n_16) );
NAND2xp33_ASAP7_75t_SL g31 ( .A(n_8), .B(n_32), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g37 ( .A(n_8), .B(n_18), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g40 ( .A(n_8), .Y(n_40) );
AOI22xp33_ASAP7_75t_SL g34 ( .A1(n_9), .A2(n_13), .B1(n_35), .B2(n_38), .Y(n_34) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_10), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_11), .Y(n_25) );
NAND2xp33_ASAP7_75t_SL g33 ( .A(n_11), .B(n_20), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g28 ( .A(n_12), .B(n_29), .Y(n_28) );
OAI221xp5_ASAP7_75t_R g14 ( .A1(n_15), .A2(n_16), .B1(n_30), .B2(n_31), .C(n_34), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_19), .B(n_26), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g19 ( .A(n_20), .B(n_25), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_21), .Y(n_20) );
NAND2xp33_ASAP7_75t_SL g21 ( .A(n_22), .B(n_24), .Y(n_21) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_26), .B(n_33), .Y(n_32) );
NAND2xp33_ASAP7_75t_SL g39 ( .A(n_32), .B(n_40), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g35 ( .A(n_36), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_37), .Y(n_36) );
INVx1_ASAP7_75t_SL g38 ( .A(n_39), .Y(n_38) );
endmodule