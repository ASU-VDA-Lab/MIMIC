module fake_jpeg_18537_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_20),
.Y(n_54)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_1),
.CON(n_42),
.SN(n_42)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_30),
.CON(n_56),
.SN(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_40),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_34),
.B1(n_25),
.B2(n_26),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_32),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_40),
.C(n_37),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_75),
.C(n_31),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_45),
.B1(n_22),
.B2(n_31),
.Y(n_106)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_76),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_28),
.B1(n_36),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_57),
.B1(n_22),
.B2(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_19),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_29),
.B(n_24),
.C(n_30),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_55),
.B(n_58),
.C(n_33),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_40),
.C(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_81),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_27),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_49),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_57),
.B1(n_51),
.B2(n_55),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_93),
.B(n_80),
.Y(n_112)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

CKINVDCx10_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_31),
.B(n_18),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_100),
.B1(n_108),
.B2(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_68),
.B1(n_64),
.B2(n_61),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_113),
.B1(n_115),
.B2(n_1),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_125),
.B1(n_104),
.B2(n_94),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_85),
.B(n_102),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_60),
.B1(n_66),
.B2(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_66),
.B1(n_74),
.B2(n_59),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_81),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_81),
.B(n_63),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_2),
.B(n_4),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_90),
.C(n_103),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_101),
.B(n_97),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_67),
.C(n_18),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_129),
.Y(n_142)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_134),
.B(n_143),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_97),
.A3(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_136),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_131),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_154),
.B1(n_115),
.B2(n_111),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_140),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_98),
.B(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_98),
.B1(n_96),
.B2(n_84),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_153),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_30),
.B1(n_18),
.B2(n_99),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_151),
.B(n_121),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_15),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_154)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_168),
.B1(n_140),
.B2(n_8),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_117),
.C(n_112),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_116),
.C(n_126),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_116),
.C(n_125),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_151),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_137),
.B1(n_134),
.B2(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_185),
.B1(n_167),
.B2(n_157),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_142),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_165),
.B(n_168),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_145),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_186),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_165),
.C(n_162),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_164),
.C(n_160),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g183 ( 
.A(n_172),
.B(n_154),
.C(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_140),
.B1(n_8),
.B2(n_9),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_159),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_198),
.C(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_164),
.B1(n_176),
.B2(n_175),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_180),
.B1(n_185),
.B2(n_171),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_155),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_201),
.Y(n_212)
);

NAND2xp67_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_192),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_161),
.C(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_140),
.B1(n_156),
.B2(n_155),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_208),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_188),
.B(n_12),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_211),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_189),
.B(n_193),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_197),
.B(n_198),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_13),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_200),
.C(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_218),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_192),
.B1(n_207),
.B2(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_221),
.A2(n_212),
.B1(n_217),
.B2(n_216),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.C(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_14),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_224),
.C(n_14),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_7),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_10),
.Y(n_229)
);


endmodule