module real_aes_12131_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_559;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_0), .A2(n_9), .B1(n_853), .B2(n_854), .C(n_856), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_0), .A2(n_9), .B1(n_460), .B2(n_869), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_1), .A2(n_258), .B1(n_359), .B2(n_446), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_1), .A2(n_258), .B1(n_511), .B2(n_582), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_2), .A2(n_16), .B1(n_574), .B2(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1109 ( .A(n_2), .Y(n_1109) );
INVx1_ASAP7_75t_L g573 ( .A(n_3), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_3), .A2(n_154), .B1(n_476), .B2(n_521), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_4), .A2(n_22), .B1(n_818), .B2(n_819), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_4), .A2(n_279), .B1(n_414), .B2(n_840), .Y(n_1022) );
INVx1_ASAP7_75t_L g1307 ( .A(n_5), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_6), .A2(n_13), .B1(n_526), .B2(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g605 ( .A(n_6), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_7), .A2(n_196), .B1(n_836), .B2(n_840), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_7), .A2(n_196), .B1(n_637), .B2(n_1148), .Y(n_1191) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_8), .Y(n_311) );
INVx1_ASAP7_75t_L g443 ( .A(n_8), .Y(n_443) );
INVx1_ASAP7_75t_L g1078 ( .A(n_10), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_11), .A2(n_273), .B1(n_813), .B2(n_816), .Y(n_812) );
INVx1_ASAP7_75t_L g844 ( .A(n_11), .Y(n_844) );
AOI22xp33_ASAP7_75t_SL g424 ( .A1(n_12), .A2(n_238), .B1(n_425), .B2(n_426), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_12), .A2(n_238), .B1(n_449), .B2(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g607 ( .A(n_13), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_14), .A2(n_50), .B1(n_912), .B2(n_914), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_14), .A2(n_50), .B1(n_732), .B2(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g884 ( .A(n_15), .Y(n_884) );
INVx1_ASAP7_75t_L g1107 ( .A(n_16), .Y(n_1107) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_17), .A2(n_48), .B1(n_636), .B2(n_638), .Y(n_635) );
INVxp67_ASAP7_75t_SL g687 ( .A(n_17), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_18), .A2(n_291), .B1(n_449), .B2(n_450), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_18), .A2(n_291), .B1(n_836), .B2(n_840), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_19), .A2(n_233), .B1(n_476), .B2(n_511), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_19), .A2(n_233), .B1(n_524), .B2(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1366 ( .A(n_20), .Y(n_1366) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_21), .Y(n_566) );
INVx1_ASAP7_75t_L g1009 ( .A(n_22), .Y(n_1009) );
CKINVDCx16_ASAP7_75t_R g1292 ( .A(n_23), .Y(n_1292) );
INVx1_ASAP7_75t_L g571 ( .A(n_24), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_24), .A2(n_293), .B1(n_516), .B2(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g329 ( .A(n_25), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_25), .A2(n_140), .B1(n_428), .B2(n_432), .Y(n_439) );
AO221x2_ASAP7_75t_L g1271 ( .A1(n_26), .A2(n_69), .B1(n_1242), .B2(n_1250), .C(n_1272), .Y(n_1271) );
XNOR2xp5_ASAP7_75t_L g972 ( .A(n_27), .B(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g1261 ( .A(n_27), .Y(n_1261) );
INVxp33_ASAP7_75t_L g1497 ( .A(n_28), .Y(n_1497) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_28), .A2(n_266), .B1(n_734), .B2(n_1123), .Y(n_1530) );
INVx2_ASAP7_75t_L g333 ( .A(n_29), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_30), .A2(n_259), .B1(n_836), .B2(n_840), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_30), .A2(n_259), .B1(n_450), .B2(n_869), .Y(n_874) );
INVxp33_ASAP7_75t_SL g625 ( .A(n_31), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_31), .A2(n_190), .B1(n_658), .B2(n_660), .Y(n_657) );
INVx1_ASAP7_75t_L g1273 ( .A(n_32), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_33), .A2(n_188), .B1(n_425), .B2(n_1201), .Y(n_1200) );
INVxp67_ASAP7_75t_SL g1226 ( .A(n_33), .Y(n_1226) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_34), .A2(n_103), .B1(n_780), .B2(n_781), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_34), .A2(n_103), .B1(n_649), .B2(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g494 ( .A(n_35), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_35), .A2(n_242), .B1(n_432), .B2(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g379 ( .A(n_36), .Y(n_379) );
BUFx2_ASAP7_75t_L g421 ( .A(n_36), .Y(n_421) );
INVx1_ASAP7_75t_L g668 ( .A(n_36), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_37), .A2(n_217), .B1(n_948), .B2(n_1209), .Y(n_1208) );
OAI211xp5_ASAP7_75t_SL g1212 ( .A1(n_37), .A2(n_489), .B(n_1213), .C(n_1216), .Y(n_1212) );
INVx1_ASAP7_75t_L g1364 ( .A(n_38), .Y(n_1364) );
AOI22xp33_ASAP7_75t_SL g949 ( .A1(n_39), .A2(n_121), .B1(n_449), .B2(n_950), .Y(n_949) );
INVxp67_ASAP7_75t_L g959 ( .A(n_39), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_40), .A2(n_275), .B1(n_630), .B2(n_633), .Y(n_629) );
INVxp67_ASAP7_75t_SL g682 ( .A(n_40), .Y(n_682) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_41), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_41), .A2(n_171), .B1(n_395), .B2(n_398), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_42), .A2(n_243), .B1(n_383), .B2(n_709), .Y(n_1084) );
AOI22xp33_ASAP7_75t_SL g1090 ( .A1(n_42), .A2(n_243), .B1(n_574), .B2(n_731), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_43), .A2(n_253), .B1(n_649), .B2(n_651), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_43), .A2(n_253), .B1(n_658), .B2(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g762 ( .A(n_44), .Y(n_762) );
INVx1_ASAP7_75t_L g887 ( .A(n_45), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_45), .A2(n_113), .B1(n_476), .B2(n_905), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_46), .A2(n_223), .B1(n_713), .B2(n_715), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_46), .A2(n_223), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g1247 ( .A(n_47), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_47), .B(n_1257), .Y(n_1260) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_48), .Y(n_688) );
INVx1_ASAP7_75t_L g889 ( .A(n_49), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_49), .A2(n_168), .B1(n_398), .B2(n_744), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_51), .A2(n_202), .B1(n_428), .B2(n_476), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_51), .A2(n_202), .B1(n_359), .B2(n_947), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_52), .A2(n_62), .B1(n_516), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_52), .A2(n_62), .B1(n_592), .B2(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g1020 ( .A(n_53), .Y(n_1020) );
INVxp67_ASAP7_75t_L g1134 ( .A(n_54), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_54), .A2(n_139), .B1(n_649), .B2(n_651), .Y(n_1152) );
CKINVDCx16_ASAP7_75t_R g1251 ( .A(n_55), .Y(n_1251) );
INVx1_ASAP7_75t_L g1506 ( .A(n_56), .Y(n_1506) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_56), .A2(n_206), .B1(n_709), .B2(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_L g1360 ( .A(n_57), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_58), .A2(n_60), .B1(n_633), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_58), .A2(n_60), .B1(n_601), .B2(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g346 ( .A(n_59), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_59), .A2(n_272), .B1(n_426), .B2(n_438), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g1075 ( .A1(n_61), .A2(n_558), .B(n_822), .C(n_1076), .Y(n_1075) );
AOI22xp33_ASAP7_75t_SL g1088 ( .A1(n_61), .A2(n_240), .B1(n_383), .B2(n_663), .Y(n_1088) );
XNOR2xp5_ASAP7_75t_L g1155 ( .A(n_63), .B(n_1156), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_64), .A2(n_271), .B1(n_476), .B2(n_709), .Y(n_1514) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_64), .A2(n_271), .B1(n_734), .B2(n_948), .Y(n_1520) );
INVx1_ASAP7_75t_L g767 ( .A(n_65), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_65), .A2(n_236), .B1(n_480), .B2(n_603), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_66), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_67), .A2(n_203), .B1(n_718), .B2(n_1082), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_67), .A2(n_203), .B1(n_1092), .B2(n_1094), .Y(n_1091) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_68), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_70), .A2(n_261), .B1(n_947), .B2(n_948), .Y(n_946) );
INVxp33_ASAP7_75t_L g961 ( .A(n_70), .Y(n_961) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_71), .A2(n_278), .B1(n_709), .B2(n_710), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_71), .A2(n_278), .B1(n_731), .B2(n_732), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_72), .A2(n_248), .B1(n_476), .B2(n_511), .Y(n_1202) );
INVx1_ASAP7_75t_L g1223 ( .A(n_72), .Y(n_1223) );
INVx1_ASAP7_75t_L g700 ( .A(n_73), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_73), .A2(n_216), .B1(n_709), .B2(n_721), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_74), .A2(n_101), .B1(n_813), .B2(n_818), .Y(n_1033) );
INVx1_ASAP7_75t_L g1050 ( .A(n_74), .Y(n_1050) );
INVx1_ASAP7_75t_L g1122 ( .A(n_75), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_75), .A2(n_97), .B1(n_383), .B2(n_795), .Y(n_1144) );
OAI22xp33_ASAP7_75t_L g1039 ( .A1(n_76), .A2(n_274), .B1(n_816), .B2(n_819), .Y(n_1039) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_76), .A2(n_274), .B1(n_713), .B2(n_1047), .C(n_1049), .Y(n_1046) );
INVx1_ASAP7_75t_L g1284 ( .A(n_77), .Y(n_1284) );
CKINVDCx16_ASAP7_75t_R g1289 ( .A(n_78), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_79), .A2(n_280), .B1(n_359), .B2(n_446), .Y(n_594) );
INVx1_ASAP7_75t_L g600 ( .A(n_79), .Y(n_600) );
INVx1_ASAP7_75t_L g1019 ( .A(n_80), .Y(n_1019) );
XOR2x2_ASAP7_75t_L g612 ( .A(n_81), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g1119 ( .A(n_82), .Y(n_1119) );
INVx1_ASAP7_75t_L g1164 ( .A(n_83), .Y(n_1164) );
INVx1_ASAP7_75t_L g985 ( .A(n_84), .Y(n_985) );
INVx1_ASAP7_75t_L g1167 ( .A(n_85), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_85), .A2(n_142), .B1(n_516), .B2(n_903), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_86), .A2(n_268), .B1(n_713), .B2(n_1512), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_86), .A2(n_268), .B1(n_1522), .B2(n_1523), .Y(n_1521) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_87), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_87), .A2(n_165), .B1(n_638), .B2(n_649), .Y(n_922) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_88), .A2(n_289), .B1(n_425), .B2(n_426), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_88), .A2(n_289), .B1(n_526), .B2(n_527), .Y(n_525) );
OAI211xp5_ASAP7_75t_L g820 ( .A1(n_89), .A2(n_558), .B(n_821), .C(n_824), .Y(n_820) );
INVx1_ASAP7_75t_L g847 ( .A(n_89), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g809 ( .A(n_90), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g1308 ( .A(n_90), .Y(n_1308) );
INVxp67_ASAP7_75t_SL g770 ( .A(n_91), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_91), .A2(n_151), .B1(n_524), .B2(n_798), .Y(n_804) );
INVx1_ASAP7_75t_L g419 ( .A(n_92), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_92), .A2(n_100), .B1(n_449), .B2(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g1495 ( .A(n_93), .Y(n_1495) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_94), .A2(n_173), .B1(n_428), .B2(n_432), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_94), .A2(n_173), .B1(n_359), .B2(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_95), .A2(n_117), .B1(n_364), .B2(n_369), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_95), .A2(n_117), .B1(n_395), .B2(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g989 ( .A(n_96), .Y(n_989) );
OAI211xp5_ASAP7_75t_SL g1023 ( .A1(n_96), .A2(n_489), .B(n_1024), .C(n_1026), .Y(n_1023) );
INVxp33_ASAP7_75t_SL g1116 ( .A(n_97), .Y(n_1116) );
INVxp33_ASAP7_75t_SL g882 ( .A(n_98), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_98), .A2(n_186), .B1(n_516), .B2(n_903), .Y(n_902) );
AO22x2_ASAP7_75t_L g468 ( .A1(n_99), .A2(n_469), .B1(n_536), .B2(n_537), .Y(n_468) );
INVxp67_ASAP7_75t_L g536 ( .A(n_99), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g1264 ( .A1(n_99), .A2(n_152), .B1(n_1265), .B2(n_1268), .Y(n_1264) );
INVx1_ASAP7_75t_L g411 ( .A(n_100), .Y(n_411) );
INVx1_ASAP7_75t_L g1065 ( .A(n_101), .Y(n_1065) );
INVx1_ASAP7_75t_L g934 ( .A(n_102), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_102), .A2(n_108), .B1(n_603), .B2(n_744), .Y(n_956) );
INVx1_ASAP7_75t_L g377 ( .A(n_104), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_105), .Y(n_859) );
INVx1_ASAP7_75t_L g1218 ( .A(n_106), .Y(n_1218) );
INVx1_ASAP7_75t_L g1229 ( .A(n_107), .Y(n_1229) );
INVx1_ASAP7_75t_L g935 ( .A(n_108), .Y(n_935) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_109), .A2(n_160), .B1(n_785), .B2(n_787), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_109), .A2(n_160), .B1(n_630), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1043 ( .A(n_110), .Y(n_1043) );
INVx1_ASAP7_75t_L g979 ( .A(n_111), .Y(n_979) );
INVxp67_ASAP7_75t_SL g1131 ( .A(n_112), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_112), .A2(n_146), .B1(n_524), .B2(n_633), .Y(n_1151) );
INVxp33_ASAP7_75t_SL g881 ( .A(n_113), .Y(n_881) );
INVx1_ASAP7_75t_L g1013 ( .A(n_114), .Y(n_1013) );
INVx1_ASAP7_75t_L g577 ( .A(n_115), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_115), .A2(n_210), .B1(n_480), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_116), .A2(n_163), .B1(n_526), .B2(n_592), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_116), .A2(n_163), .B1(n_836), .B2(n_840), .Y(n_1211) );
INVx1_ASAP7_75t_L g472 ( .A(n_118), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_118), .A2(n_252), .B1(n_449), .B2(n_460), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_119), .A2(n_231), .B1(n_511), .B2(n_512), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_119), .A2(n_231), .B1(n_457), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1258 ( .A(n_120), .Y(n_1258) );
INVxp33_ASAP7_75t_L g958 ( .A(n_121), .Y(n_958) );
AO221x2_ASAP7_75t_L g1305 ( .A1(n_122), .A2(n_201), .B1(n_1250), .B2(n_1291), .C(n_1306), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g857 ( .A(n_123), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_124), .A2(n_256), .B1(n_425), .B2(n_426), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_124), .A2(n_256), .B1(n_590), .B2(n_592), .Y(n_589) );
INVx1_ASAP7_75t_L g988 ( .A(n_125), .Y(n_988) );
OAI22xp33_ASAP7_75t_SL g1027 ( .A1(n_125), .A2(n_169), .B1(n_312), .B2(n_836), .Y(n_1027) );
AO22x2_ASAP7_75t_L g924 ( .A1(n_126), .A2(n_925), .B1(n_962), .B2(n_963), .Y(n_924) );
INVx1_ASAP7_75t_L g962 ( .A(n_126), .Y(n_962) );
INVx1_ASAP7_75t_L g703 ( .A(n_127), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_127), .A2(n_156), .B1(n_603), .B2(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g303 ( .A(n_128), .Y(n_303) );
INVx1_ASAP7_75t_L g403 ( .A(n_129), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_129), .A2(n_229), .B1(n_446), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_130), .A2(n_193), .B1(n_1101), .B2(n_1103), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_130), .A2(n_193), .B1(n_836), .B2(n_840), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_131), .A2(n_232), .B1(n_719), .B2(n_780), .C(n_1042), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_131), .A2(n_232), .B1(n_449), .B2(n_460), .Y(n_1055) );
INVx1_ASAP7_75t_L g1038 ( .A(n_132), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_133), .A2(n_217), .B1(n_312), .B2(n_414), .Y(n_1219) );
OAI22xp33_ASAP7_75t_L g1228 ( .A1(n_133), .A2(n_248), .B1(n_813), .B2(n_818), .Y(n_1228) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_134), .A2(n_192), .B1(n_1242), .B2(n_1250), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_135), .A2(n_167), .B1(n_818), .B2(n_819), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g842 ( .A1(n_135), .A2(n_273), .B1(n_713), .B2(n_715), .C(n_843), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_136), .Y(n_487) );
XNOR2xp5_ASAP7_75t_L g1070 ( .A(n_137), .B(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g937 ( .A(n_138), .Y(n_937) );
INVxp67_ASAP7_75t_L g1135 ( .A(n_139), .Y(n_1135) );
INVx1_ASAP7_75t_L g362 ( .A(n_140), .Y(n_362) );
INVxp33_ASAP7_75t_SL g773 ( .A(n_141), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_141), .A2(n_166), .B1(n_806), .B2(n_807), .Y(n_805) );
INVxp67_ASAP7_75t_SL g1166 ( .A(n_142), .Y(n_1166) );
INVxp67_ASAP7_75t_SL g1126 ( .A(n_143), .Y(n_1126) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_143), .A2(n_296), .B1(n_398), .B2(n_744), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_144), .A2(n_285), .B1(n_633), .B2(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_SL g742 ( .A(n_144), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_145), .A2(n_149), .B1(n_460), .B2(n_869), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_145), .A2(n_149), .B1(n_425), .B2(n_426), .Y(n_951) );
INVxp67_ASAP7_75t_SL g1129 ( .A(n_146), .Y(n_1129) );
INVx1_ASAP7_75t_L g1274 ( .A(n_147), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1535 ( .A1(n_147), .A2(n_1536), .B1(n_1540), .B2(n_1543), .Y(n_1535) );
CKINVDCx14_ASAP7_75t_R g1030 ( .A(n_148), .Y(n_1030) );
INVx1_ASAP7_75t_L g1037 ( .A(n_150), .Y(n_1037) );
INVxp33_ASAP7_75t_L g776 ( .A(n_151), .Y(n_776) );
INVxp33_ASAP7_75t_SL g928 ( .A(n_153), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_153), .A2(n_175), .B1(n_428), .B2(n_582), .Y(n_944) );
INVx1_ASAP7_75t_L g570 ( .A(n_154), .Y(n_570) );
INVxp33_ASAP7_75t_SL g695 ( .A(n_155), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_155), .A2(n_215), .B1(n_718), .B2(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g702 ( .A(n_156), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_157), .A2(n_269), .B1(n_818), .B2(n_819), .Y(n_1074) );
INVxp33_ASAP7_75t_SL g1110 ( .A(n_157), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_158), .A2(n_170), .B1(n_425), .B2(n_1197), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_158), .A2(n_170), .B1(n_527), .B2(n_637), .Y(n_1205) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_159), .A2(n_212), .B1(n_813), .B2(n_818), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_159), .A2(n_247), .B1(n_521), .B2(n_914), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_161), .A2(n_240), .B1(n_813), .B2(n_816), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_161), .A2(n_269), .B1(n_660), .B2(n_718), .Y(n_1087) );
INVxp33_ASAP7_75t_SL g760 ( .A(n_162), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_162), .A2(n_245), .B1(n_790), .B2(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g982 ( .A(n_164), .Y(n_982) );
INVxp33_ASAP7_75t_L g896 ( .A(n_165), .Y(n_896) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_166), .Y(n_774) );
INVx1_ASAP7_75t_L g834 ( .A(n_167), .Y(n_834) );
INVx1_ASAP7_75t_L g888 ( .A(n_168), .Y(n_888) );
INVx1_ASAP7_75t_L g992 ( .A(n_169), .Y(n_992) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_171), .Y(n_622) );
INVxp67_ASAP7_75t_SL g1502 ( .A(n_172), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_172), .A2(n_228), .B1(n_718), .B2(n_1047), .Y(n_1516) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_174), .A2(n_182), .B1(n_1265), .B2(n_1268), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_175), .Y(n_931) );
INVxp33_ASAP7_75t_SL g938 ( .A(n_176), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g943 ( .A1(n_176), .A2(n_197), .B1(n_425), .B2(n_426), .Y(n_943) );
INVxp33_ASAP7_75t_SL g1117 ( .A(n_177), .Y(n_1117) );
AOI22xp33_ASAP7_75t_SL g1142 ( .A1(n_177), .A2(n_276), .B1(n_853), .B2(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g697 ( .A(n_178), .Y(n_697) );
INVx1_ASAP7_75t_L g1008 ( .A(n_179), .Y(n_1008) );
OAI22xp33_ASAP7_75t_L g1015 ( .A1(n_179), .A2(n_195), .B1(n_813), .B2(n_816), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_180), .A2(n_270), .B1(n_511), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_180), .A2(n_270), .B1(n_359), .B2(n_446), .Y(n_588) );
INVx1_ASAP7_75t_L g624 ( .A(n_181), .Y(n_624) );
XNOR2xp5_ASAP7_75t_L g1112 ( .A(n_182), .B(n_1113), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1300 ( .A1(n_183), .A2(n_239), .B1(n_1291), .B2(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1490 ( .A(n_184), .Y(n_1490) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_185), .Y(n_305) );
AND3x2_ASAP7_75t_L g1243 ( .A(n_185), .B(n_303), .C(n_1244), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_185), .B(n_303), .Y(n_1255) );
INVxp33_ASAP7_75t_SL g885 ( .A(n_186), .Y(n_885) );
INVxp33_ASAP7_75t_SL g899 ( .A(n_187), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_187), .A2(n_254), .B1(n_732), .B2(n_917), .Y(n_921) );
INVx1_ASAP7_75t_L g1227 ( .A(n_188), .Y(n_1227) );
INVx1_ASAP7_75t_L g1163 ( .A(n_189), .Y(n_1163) );
INVxp33_ASAP7_75t_SL g617 ( .A(n_190), .Y(n_617) );
INVx2_ASAP7_75t_L g316 ( .A(n_191), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_194), .A2(n_263), .B1(n_660), .B2(n_853), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_194), .A2(n_263), .B1(n_650), .B2(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1012 ( .A(n_195), .Y(n_1012) );
INVxp33_ASAP7_75t_SL g929 ( .A(n_197), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g1295 ( .A1(n_198), .A2(n_205), .B1(n_1242), .B2(n_1250), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_199), .A2(n_213), .B1(n_795), .B2(n_1140), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_199), .A2(n_213), .B1(n_633), .B2(n_731), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_200), .A2(n_226), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_200), .A2(n_226), .B1(n_637), .B2(n_1148), .Y(n_1188) );
INVx1_ASAP7_75t_L g1244 ( .A(n_204), .Y(n_1244) );
INVxp33_ASAP7_75t_L g1501 ( .A(n_206), .Y(n_1501) );
INVxp67_ASAP7_75t_SL g1491 ( .A(n_207), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_207), .A2(n_249), .B1(n_460), .B2(n_1528), .Y(n_1527) );
CKINVDCx16_ASAP7_75t_R g1248 ( .A(n_208), .Y(n_1248) );
OAI211xp5_ASAP7_75t_L g1171 ( .A1(n_209), .A2(n_489), .B(n_1024), .C(n_1172), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_209), .A2(n_292), .B1(n_446), .B2(n_1186), .Y(n_1190) );
INVx1_ASAP7_75t_L g575 ( .A(n_210), .Y(n_575) );
INVx1_ASAP7_75t_L g1362 ( .A(n_211), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_212), .A2(n_292), .B1(n_312), .B2(n_414), .Y(n_1173) );
INVx1_ASAP7_75t_L g503 ( .A(n_214), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_214), .A2(n_260), .B1(n_516), .B2(n_517), .Y(n_515) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_215), .Y(n_698) );
INVxp33_ASAP7_75t_SL g694 ( .A(n_216), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_218), .Y(n_825) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_219), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_219), .A2(n_282), .B1(n_582), .B2(n_795), .Y(n_794) );
XNOR2xp5_ASAP7_75t_L g1541 ( .A(n_220), .B(n_1542), .Y(n_1541) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_221), .Y(n_341) );
INVx1_ASAP7_75t_L g1057 ( .A(n_222), .Y(n_1057) );
INVx1_ASAP7_75t_L g318 ( .A(n_224), .Y(n_318) );
INVx2_ASAP7_75t_L g393 ( .A(n_224), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g1034 ( .A1(n_225), .A2(n_558), .B(n_1035), .C(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1051 ( .A(n_225), .Y(n_1051) );
XNOR2xp5_ASAP7_75t_L g325 ( .A(n_227), .B(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_SL g1504 ( .A(n_228), .Y(n_1504) );
INVx1_ASAP7_75t_L g382 ( .A(n_229), .Y(n_382) );
INVx1_ASAP7_75t_L g475 ( .A(n_230), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_230), .A2(n_288), .B1(n_531), .B2(n_533), .Y(n_530) );
OAI211xp5_ASAP7_75t_L g540 ( .A1(n_230), .A2(n_489), .B(n_541), .C(n_546), .Y(n_540) );
XNOR2xp5_ASAP7_75t_L g562 ( .A(n_234), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g1045 ( .A(n_235), .Y(n_1045) );
INVx1_ASAP7_75t_L g766 ( .A(n_236), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g1294 ( .A1(n_237), .A2(n_265), .B1(n_1265), .B2(n_1268), .Y(n_1294) );
CKINVDCx20_ASAP7_75t_R g1493 ( .A(n_241), .Y(n_1493) );
INVx1_ASAP7_75t_L g498 ( .A(n_242), .Y(n_498) );
OAI211xp5_ASAP7_75t_L g552 ( .A1(n_242), .A2(n_553), .B(n_558), .C(n_559), .Y(n_552) );
AO22x2_ASAP7_75t_SL g689 ( .A1(n_244), .A2(n_690), .B1(n_691), .B2(n_750), .Y(n_689) );
CKINVDCx16_ASAP7_75t_R g690 ( .A(n_244), .Y(n_690) );
INVxp33_ASAP7_75t_L g763 ( .A(n_245), .Y(n_763) );
INVxp33_ASAP7_75t_SL g616 ( .A(n_246), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_246), .A2(n_281), .B1(n_601), .B2(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g1160 ( .A(n_247), .Y(n_1160) );
INVxp67_ASAP7_75t_SL g1498 ( .A(n_249), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_250), .Y(n_826) );
INVx1_ASAP7_75t_L g1285 ( .A(n_251), .Y(n_1285) );
INVx1_ASAP7_75t_L g473 ( .A(n_252), .Y(n_473) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_254), .Y(n_893) );
INVx1_ASAP7_75t_L g1077 ( .A(n_255), .Y(n_1077) );
XOR2x2_ASAP7_75t_L g877 ( .A(n_257), .B(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g495 ( .A(n_260), .Y(n_495) );
INVxp67_ASAP7_75t_SL g955 ( .A(n_261), .Y(n_955) );
INVx1_ASAP7_75t_L g977 ( .A(n_262), .Y(n_977) );
INVx1_ASAP7_75t_L g1217 ( .A(n_264), .Y(n_1217) );
INVxp67_ASAP7_75t_SL g1494 ( .A(n_266), .Y(n_1494) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_267), .Y(n_481) );
INVx1_ASAP7_75t_L g352 ( .A(n_272), .Y(n_352) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_275), .Y(n_685) );
INVxp67_ASAP7_75t_SL g1120 ( .A(n_276), .Y(n_1120) );
INVx2_ASAP7_75t_L g315 ( .A(n_277), .Y(n_315) );
INVx1_ASAP7_75t_L g994 ( .A(n_279), .Y(n_994) );
INVx1_ASAP7_75t_L g609 ( .A(n_280), .Y(n_609) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_281), .Y(n_619) );
INVxp33_ASAP7_75t_L g759 ( .A(n_282), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_283), .A2(n_294), .B1(n_737), .B2(n_738), .Y(n_736) );
INVxp33_ASAP7_75t_L g746 ( .A(n_283), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_284), .Y(n_830) );
INVxp33_ASAP7_75t_L g749 ( .A(n_285), .Y(n_749) );
BUFx3_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g356 ( .A(n_286), .Y(n_356) );
BUFx3_ASAP7_75t_L g340 ( .A(n_287), .Y(n_340) );
INVx1_ASAP7_75t_L g351 ( .A(n_287), .Y(n_351) );
INVx1_ASAP7_75t_L g486 ( .A(n_288), .Y(n_486) );
INVx1_ASAP7_75t_L g1058 ( .A(n_290), .Y(n_1058) );
INVx1_ASAP7_75t_L g567 ( .A(n_293), .Y(n_567) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_294), .Y(n_747) );
AO22x1_ASAP7_75t_L g754 ( .A1(n_295), .A2(n_755), .B1(n_756), .B2(n_808), .Y(n_754) );
INVxp67_ASAP7_75t_L g755 ( .A(n_295), .Y(n_755) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_296), .Y(n_1125) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_319), .B(n_1232), .Y(n_297) );
BUFx12f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_306), .Y(n_300) );
AND2x4_ASAP7_75t_L g1534 ( .A(n_301), .B(n_307), .Y(n_1534) );
NOR2xp33_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g1539 ( .A(n_302), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1546 ( .A(n_302), .B(n_304), .Y(n_1546) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_304), .B(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g420 ( .A(n_309), .B(n_421), .Y(n_420) );
OR2x6_ASAP7_75t_L g491 ( .A(n_309), .B(n_421), .Y(n_491) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g435 ( .A(n_310), .B(n_318), .Y(n_435) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_311), .B(n_406), .Y(n_1001) );
INVx8_ASAP7_75t_L g402 ( .A(n_312), .Y(n_402) );
OR2x6_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
OR2x6_ASAP7_75t_L g414 ( .A(n_313), .B(n_405), .Y(n_414) );
INVx2_ASAP7_75t_SL g846 ( .A(n_313), .Y(n_846) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_313), .Y(n_858) );
INVx2_ASAP7_75t_SL g999 ( .A(n_313), .Y(n_999) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_313), .Y(n_1044) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g387 ( .A(n_315), .Y(n_387) );
INVx1_ASAP7_75t_L g400 ( .A(n_315), .Y(n_400) );
INVx2_ASAP7_75t_L g408 ( .A(n_315), .Y(n_408) );
AND2x4_ASAP7_75t_L g418 ( .A(n_315), .B(n_388), .Y(n_418) );
AND2x2_ASAP7_75t_L g431 ( .A(n_315), .B(n_316), .Y(n_431) );
INVx2_ASAP7_75t_L g388 ( .A(n_316), .Y(n_388) );
INVx1_ASAP7_75t_L g397 ( .A(n_316), .Y(n_397) );
INVx1_ASAP7_75t_L g410 ( .A(n_316), .Y(n_410) );
INVx1_ASAP7_75t_L g545 ( .A(n_316), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_316), .B(n_408), .Y(n_839) );
AND2x4_ASAP7_75t_L g396 ( .A(n_317), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g398 ( .A(n_318), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g603 ( .A(n_318), .B(n_399), .Y(n_603) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B1(n_968), .B2(n_1231), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
XNOR2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_464), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI211xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_375), .B(n_380), .C(n_422), .Y(n_326) );
NAND4xp25_ASAP7_75t_L g327 ( .A(n_328), .B(n_345), .C(n_357), .D(n_372), .Y(n_327) );
AOI22xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_330), .B1(n_341), .B2(n_342), .Y(n_328) );
AOI22xp5_ASAP7_75t_SL g493 ( .A1(n_330), .A2(n_347), .B1(n_494), .B2(n_495), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_330), .A2(n_347), .B1(n_759), .B2(n_760), .Y(n_758) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
AND2x6_ASAP7_75t_L g353 ( .A(n_331), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g569 ( .A(n_331), .B(n_334), .Y(n_569) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g365 ( .A(n_332), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_333), .Y(n_344) );
INVx1_ASAP7_75t_L g349 ( .A(n_333), .Y(n_349) );
AND2x2_ASAP7_75t_L g454 ( .A(n_333), .B(n_377), .Y(n_454) );
INVx2_ASAP7_75t_L g463 ( .A(n_333), .Y(n_463) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_335), .Y(n_532) );
INVx2_ASAP7_75t_SL g632 ( .A(n_335), .Y(n_632) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_335), .Y(n_647) );
INVx2_ASAP7_75t_L g735 ( .A(n_335), .Y(n_735) );
INVx1_ASAP7_75t_L g1209 ( .A(n_335), .Y(n_1209) );
INVx6_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g342 ( .A(n_336), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g447 ( .A(n_336), .Y(n_447) );
BUFx2_ASAP7_75t_L g524 ( .A(n_336), .Y(n_524) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g350 ( .A(n_338), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g361 ( .A(n_338), .B(n_340), .Y(n_361) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g355 ( .A(n_340), .B(n_356), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_341), .A2(n_413), .B1(n_415), .B2(n_419), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_342), .A2(n_353), .B1(n_487), .B2(n_503), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_342), .A2(n_353), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_342), .A2(n_353), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_342), .A2(n_353), .B1(n_697), .B2(n_698), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_342), .A2(n_353), .B1(n_762), .B2(n_763), .Y(n_761) );
INVx4_ASAP7_75t_L g818 ( .A(n_342), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_342), .A2(n_353), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_342), .A2(n_353), .B1(n_937), .B2(n_938), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_342), .A2(n_353), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_342), .A2(n_353), .B1(n_1490), .B2(n_1504), .Y(n_1503) );
AND2x4_ASAP7_75t_L g500 ( .A(n_343), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_343), .B(n_501), .Y(n_576) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_352), .B2(n_353), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_347), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_347), .A2(n_373), .B1(n_569), .B2(n_616), .C(n_617), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_347), .A2(n_569), .B1(n_694), .B2(n_695), .Y(n_693) );
CKINVDCx6p67_ASAP7_75t_R g816 ( .A(n_347), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_347), .A2(n_569), .B1(n_881), .B2(n_882), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_347), .A2(n_569), .B1(n_928), .B2(n_929), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_347), .A2(n_569), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_347), .A2(n_353), .B1(n_1166), .B2(n_1167), .Y(n_1165) );
AOI22xp5_ASAP7_75t_L g1225 ( .A1(n_347), .A2(n_353), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_347), .A2(n_569), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
AND2x6_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AND2x2_ASAP7_75t_L g358 ( .A(n_348), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
INVx1_ASAP7_75t_L g814 ( .A(n_348), .Y(n_814) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x6_ASAP7_75t_L g370 ( .A(n_349), .B(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g449 ( .A(n_350), .Y(n_449) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_350), .Y(n_526) );
INVx2_ASAP7_75t_SL g591 ( .A(n_350), .Y(n_591) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_350), .Y(n_637) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_350), .Y(n_650) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_350), .Y(n_727) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_350), .Y(n_806) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_350), .Y(n_869) );
BUFx2_ASAP7_75t_L g919 ( .A(n_350), .Y(n_919) );
INVx1_ASAP7_75t_L g557 ( .A(n_351), .Y(n_557) );
INVx4_ASAP7_75t_L g819 ( .A(n_353), .Y(n_819) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_354), .Y(n_460) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_354), .Y(n_592) );
INVx1_ASAP7_75t_L g597 ( .A(n_354), .Y(n_597) );
INVx1_ASAP7_75t_L g652 ( .A(n_354), .Y(n_652) );
INVx1_ASAP7_75t_L g802 ( .A(n_354), .Y(n_802) );
INVx2_ASAP7_75t_L g993 ( .A(n_354), .Y(n_993) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_355), .Y(n_450) );
INVx1_ASAP7_75t_L g528 ( .A(n_355), .Y(n_528) );
INVx2_ASAP7_75t_L g641 ( .A(n_355), .Y(n_641) );
INVx1_ASAP7_75t_L g729 ( .A(n_355), .Y(n_729) );
INVx1_ASAP7_75t_L g556 ( .A(n_356), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_362), .B(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g1035 ( .A(n_358), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_359), .Y(n_497) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_359), .Y(n_701) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g373 ( .A(n_360), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g534 ( .A(n_360), .Y(n_534) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_360), .Y(n_634) );
INVx2_ASAP7_75t_L g799 ( .A(n_360), .Y(n_799) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_361), .Y(n_458) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI222xp33_ASAP7_75t_L g1018 ( .A1(n_365), .A2(n_370), .B1(n_798), .B2(n_1013), .C1(n_1019), .C2(n_1020), .Y(n_1018) );
AOI222xp33_ASAP7_75t_L g1222 ( .A1(n_365), .A2(n_370), .B1(n_1217), .B2(n_1218), .C1(n_1223), .C2(n_1224), .Y(n_1222) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g501 ( .A(n_367), .Y(n_501) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g496 ( .A1(n_370), .A2(n_478), .B1(n_481), .B2(n_497), .C1(n_498), .C2(n_499), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_370), .A2(n_478), .B1(n_481), .B2(n_500), .Y(n_559) );
AOI222xp33_ASAP7_75t_L g572 ( .A1(n_370), .A2(n_573), .B1(n_574), .B2(n_575), .C1(n_576), .C2(n_577), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g618 ( .A1(n_370), .A2(n_576), .B1(n_619), .B2(n_620), .C1(n_621), .C2(n_622), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_370), .A2(n_499), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_703), .Y(n_699) );
AOI222xp33_ASAP7_75t_L g764 ( .A1(n_370), .A2(n_457), .B1(n_576), .B2(n_765), .C1(n_766), .C2(n_767), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_370), .A2(n_500), .B1(n_825), .B2(n_826), .Y(n_824) );
AOI222xp33_ASAP7_75t_L g886 ( .A1(n_370), .A2(n_576), .B1(n_633), .B2(n_887), .C1(n_888), .C2(n_889), .Y(n_886) );
AOI222xp33_ASAP7_75t_L g930 ( .A1(n_370), .A2(n_576), .B1(n_931), .B2(n_932), .C1(n_934), .C2(n_935), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_370), .A2(n_500), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g1076 ( .A1(n_370), .A2(n_500), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
AOI222xp33_ASAP7_75t_L g1121 ( .A1(n_370), .A2(n_576), .B1(n_1122), .B2(n_1123), .C1(n_1125), .C2(n_1126), .Y(n_1121) );
AOI222xp33_ASAP7_75t_L g1159 ( .A1(n_370), .A2(n_576), .B1(n_1160), .B2(n_1161), .C1(n_1163), .C2(n_1164), .Y(n_1159) );
AOI222xp33_ASAP7_75t_L g1505 ( .A1(n_370), .A2(n_499), .B1(n_1493), .B2(n_1495), .C1(n_1506), .C2(n_1507), .Y(n_1505) );
NAND4xp25_ASAP7_75t_L g492 ( .A(n_372), .B(n_493), .C(n_496), .D(n_502), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g564 ( .A(n_372), .B(n_565), .C(n_568), .D(n_572), .Y(n_564) );
NAND4xp25_ASAP7_75t_SL g692 ( .A(n_372), .B(n_693), .C(n_696), .D(n_699), .Y(n_692) );
NAND4xp25_ASAP7_75t_SL g757 ( .A(n_372), .B(n_758), .C(n_761), .D(n_764), .Y(n_757) );
NAND4xp25_ASAP7_75t_L g1499 ( .A(n_372), .B(n_1500), .C(n_1503), .D(n_1505), .Y(n_1499) );
INVx5_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
CKINVDCx8_ASAP7_75t_R g558 ( .A(n_373), .Y(n_558) );
AOI211xp5_ASAP7_75t_L g563 ( .A1(n_375), .A2(n_564), .B(n_578), .C(n_598), .Y(n_563) );
OAI31xp33_ASAP7_75t_SL g811 ( .A1(n_375), .A2(n_812), .A3(n_817), .B(n_820), .Y(n_811) );
AOI211x1_ASAP7_75t_L g925 ( .A1(n_375), .A2(n_926), .B(n_939), .C(n_953), .Y(n_925) );
OAI31xp33_ASAP7_75t_L g1014 ( .A1(n_375), .A2(n_1015), .A3(n_1016), .B(n_1017), .Y(n_1014) );
OAI31xp33_ASAP7_75t_L g1032 ( .A1(n_375), .A2(n_1033), .A3(n_1034), .B(n_1039), .Y(n_1032) );
OAI31xp33_ASAP7_75t_L g1072 ( .A1(n_375), .A2(n_1073), .A3(n_1074), .B(n_1075), .Y(n_1072) );
OAI21xp5_ASAP7_75t_L g1157 ( .A1(n_375), .A2(n_1158), .B(n_1168), .Y(n_1157) );
OAI21xp5_ASAP7_75t_SL g1220 ( .A1(n_375), .A2(n_1221), .B(n_1228), .Y(n_1220) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
AND2x4_ASAP7_75t_L g505 ( .A(n_376), .B(n_378), .Y(n_505) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g462 ( .A(n_377), .B(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g434 ( .A(n_379), .Y(n_434) );
OR2x6_ASAP7_75t_L g1000 ( .A(n_379), .B(n_1001), .Y(n_1000) );
AOI31xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_401), .A3(n_412), .B(n_420), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_389), .C(n_394), .Y(n_381) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g914 ( .A(n_384), .Y(n_914) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_385), .Y(n_787) );
AOI222xp33_ASAP7_75t_L g1106 ( .A1(n_385), .A2(n_396), .B1(n_482), .B2(n_1077), .C1(n_1078), .C2(n_1107), .Y(n_1106) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_385), .Y(n_1140) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g389 ( .A(n_386), .B(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g432 ( .A(n_386), .Y(n_432) );
BUFx3_ASAP7_75t_L g477 ( .A(n_386), .Y(n_477) );
INVx1_ASAP7_75t_L g513 ( .A(n_386), .Y(n_513) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_386), .Y(n_582) );
BUFx2_ASAP7_75t_L g723 ( .A(n_386), .Y(n_723) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
CKINVDCx11_ASAP7_75t_R g489 ( .A(n_389), .Y(n_489) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_389), .A2(n_600), .B(n_601), .C(n_602), .Y(n_599) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_389), .A2(n_476), .B(n_682), .C(n_683), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g741 ( .A1(n_389), .A2(n_476), .B(n_742), .C(n_743), .Y(n_741) );
AOI211xp5_ASAP7_75t_L g769 ( .A1(n_389), .A2(n_601), .B(n_770), .C(n_771), .Y(n_769) );
AOI211xp5_ASAP7_75t_L g891 ( .A1(n_389), .A2(n_892), .B(n_893), .C(n_894), .Y(n_891) );
AOI211xp5_ASAP7_75t_L g954 ( .A1(n_389), .A2(n_601), .B(n_955), .C(n_956), .Y(n_954) );
AOI211xp5_ASAP7_75t_L g1130 ( .A1(n_389), .A2(n_512), .B(n_1131), .C(n_1132), .Y(n_1130) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g484 ( .A(n_391), .Y(n_484) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_392), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g406 ( .A(n_393), .Y(n_406) );
INVx1_ASAP7_75t_L g547 ( .A(n_395), .Y(n_547) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g480 ( .A(n_396), .Y(n_480) );
INVx2_ASAP7_75t_L g744 ( .A(n_396), .Y(n_744) );
AOI222xp33_ASAP7_75t_SL g829 ( .A1(n_396), .A2(n_482), .B1(n_825), .B2(n_826), .C1(n_830), .C2(n_831), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_396), .A2(n_548), .B1(n_1019), .B2(n_1020), .Y(n_1026) );
AOI222xp33_ASAP7_75t_L g1062 ( .A1(n_396), .A2(n_548), .B1(n_1037), .B2(n_1038), .C1(n_1058), .C2(n_1063), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_396), .A2(n_548), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
INVx1_ASAP7_75t_L g483 ( .A(n_399), .Y(n_483) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g544 ( .A(n_400), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_400), .B(n_545), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_404), .B2(n_411), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_402), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_402), .A2(n_488), .B1(n_566), .B2(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_402), .A2(n_488), .B1(n_624), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_402), .A2(n_413), .B1(n_697), .B2(n_749), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_402), .A2(n_413), .B1(n_762), .B2(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_402), .A2(n_488), .B1(n_833), .B2(n_834), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_402), .A2(n_413), .B1(n_884), .B2(n_899), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g960 ( .A1(n_402), .A2(n_413), .B1(n_937), .B2(n_961), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_402), .A2(n_488), .B1(n_1057), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_402), .A2(n_488), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
AOI22xp5_ASAP7_75t_L g1128 ( .A1(n_402), .A2(n_413), .B1(n_1119), .B2(n_1129), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1496 ( .A1(n_402), .A2(n_606), .B1(n_1497), .B2(n_1498), .Y(n_1496) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_404), .A2(n_415), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_404), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_604) );
AOI22xp5_ASAP7_75t_SL g686 ( .A1(n_404), .A2(n_606), .B1(n_687), .B2(n_688), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_404), .A2(n_415), .B1(n_746), .B2(n_747), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_404), .A2(n_606), .B1(n_773), .B2(n_774), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_404), .A2(n_606), .B1(n_896), .B2(n_897), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g957 ( .A1(n_404), .A2(n_606), .B1(n_958), .B2(n_959), .Y(n_957) );
AOI22xp5_ASAP7_75t_SL g1133 ( .A1(n_404), .A2(n_415), .B1(n_1134), .B2(n_1135), .Y(n_1133) );
AOI22xp33_ASAP7_75t_SL g1489 ( .A1(n_404), .A2(n_488), .B1(n_1490), .B2(n_1491), .Y(n_1489) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
AND2x4_ASAP7_75t_L g415 ( .A(n_405), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g606 ( .A(n_405), .B(n_416), .Y(n_606) );
INVx1_ASAP7_75t_L g837 ( .A(n_405), .Y(n_837) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_407), .Y(n_425) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_407), .Y(n_516) );
INVx1_ASAP7_75t_L g659 ( .A(n_407), .Y(n_659) );
BUFx2_ASAP7_75t_L g718 ( .A(n_407), .Y(n_718) );
BUFx2_ASAP7_75t_L g780 ( .A(n_407), .Y(n_780) );
INVx1_ASAP7_75t_L g791 ( .A(n_407), .Y(n_791) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx5_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx4_ASAP7_75t_L g488 ( .A(n_414), .Y(n_488) );
INVx5_ASAP7_75t_SL g840 ( .A(n_415), .Y(n_840) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_418), .Y(n_426) );
INVx3_ASAP7_75t_L g519 ( .A(n_418), .Y(n_519) );
INVx1_ASAP7_75t_L g674 ( .A(n_418), .Y(n_674) );
AOI31xp33_ASAP7_75t_L g953 ( .A1(n_420), .A2(n_954), .A3(n_957), .B(n_960), .Y(n_953) );
AND2x4_ASAP7_75t_L g461 ( .A(n_421), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g643 ( .A(n_421), .B(n_462), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g422 ( .A(n_423), .B(n_436), .C(n_444), .D(n_455), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .C(n_433), .Y(n_423) );
INVx2_ASAP7_75t_SL g716 ( .A(n_426), .Y(n_716) );
BUFx3_ASAP7_75t_L g719 ( .A(n_426), .Y(n_719) );
INVx2_ASAP7_75t_SL g1048 ( .A(n_426), .Y(n_1048) );
INVx4_ASAP7_75t_L g1083 ( .A(n_426), .Y(n_1083) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g511 ( .A(n_429), .Y(n_511) );
INVx2_ASAP7_75t_L g905 ( .A(n_429), .Y(n_905) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g521 ( .A(n_430), .Y(n_521) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g664 ( .A(n_431), .Y(n_664) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_432), .Y(n_1063) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_433), .B(n_509), .C(n_510), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_433), .B(n_580), .C(n_581), .Y(n_579) );
INVx2_ASAP7_75t_L g707 ( .A(n_433), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_433), .B(n_779), .C(n_784), .Y(n_778) );
BUFx3_ASAP7_75t_L g860 ( .A(n_433), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_433), .B(n_907), .C(n_911), .Y(n_906) );
AOI33xp33_ASAP7_75t_L g945 ( .A1(n_433), .A2(n_461), .A3(n_946), .B1(n_949), .B2(n_951), .B3(n_952), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g1137 ( .A(n_433), .B(n_1138), .C(n_1139), .Y(n_1137) );
NAND3xp33_ASAP7_75t_L g1175 ( .A(n_433), .B(n_1176), .C(n_1180), .Y(n_1175) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_433), .B(n_1196), .C(n_1198), .Y(n_1195) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AND2x2_ASAP7_75t_L g440 ( .A(n_434), .B(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g452 ( .A(n_434), .B(n_453), .Y(n_452) );
OR2x6_ASAP7_75t_L g654 ( .A(n_434), .B(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g679 ( .A(n_434), .B(n_435), .Y(n_679) );
OR2x2_ASAP7_75t_L g862 ( .A(n_434), .B(n_655), .Y(n_862) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .C(n_440), .Y(n_436) );
INVx2_ASAP7_75t_SL g714 ( .A(n_438), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_440), .B(n_515), .C(n_520), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_440), .B(n_584), .C(n_586), .Y(n_583) );
AOI33xp33_ASAP7_75t_L g940 ( .A1(n_440), .A2(n_451), .A3(n_941), .B1(n_942), .B2(n_943), .B3(n_944), .Y(n_940) );
INVx1_ASAP7_75t_L g1010 ( .A(n_440), .Y(n_1010) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x6_ASAP7_75t_L g666 ( .A(n_442), .B(n_667), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .C(n_451), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g947 ( .A(n_447), .Y(n_947) );
INVx2_ASAP7_75t_SL g1529 ( .A(n_449), .Y(n_1529) );
INVx1_ASAP7_75t_L g980 ( .A(n_450), .Y(n_980) );
INVx1_ASAP7_75t_L g1095 ( .A(n_450), .Y(n_1095) );
BUFx6f_ASAP7_75t_L g1148 ( .A(n_450), .Y(n_1148) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_451), .B(n_523), .C(n_525), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_451), .B(n_588), .C(n_589), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_451), .B(n_797), .C(n_800), .Y(n_796) );
NAND3xp33_ASAP7_75t_L g915 ( .A(n_451), .B(n_916), .C(n_918), .Y(n_915) );
NAND3xp33_ASAP7_75t_L g1184 ( .A(n_451), .B(n_1185), .C(n_1188), .Y(n_1184) );
NAND3xp33_ASAP7_75t_L g1203 ( .A(n_451), .B(n_1204), .C(n_1205), .Y(n_1203) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g655 ( .A(n_454), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_459), .C(n_461), .Y(n_455) );
BUFx2_ASAP7_75t_SL g620 ( .A(n_457), .Y(n_620) );
INVx1_ASAP7_75t_L g1124 ( .A(n_457), .Y(n_1124) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g574 ( .A(n_458), .Y(n_574) );
BUFx4f_ASAP7_75t_L g732 ( .A(n_458), .Y(n_732) );
INVx1_ASAP7_75t_L g933 ( .A(n_458), .Y(n_933) );
INVx1_ASAP7_75t_L g1162 ( .A(n_458), .Y(n_1162) );
INVx2_ASAP7_75t_SL g1187 ( .A(n_458), .Y(n_1187) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_461), .B(n_530), .C(n_535), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_461), .B(n_594), .C(n_595), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_461), .B(n_804), .C(n_805), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_461), .B(n_921), .C(n_922), .Y(n_920) );
INVx1_ASAP7_75t_L g995 ( .A(n_461), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g1189 ( .A(n_461), .B(n_1190), .C(n_1191), .Y(n_1189) );
NAND3xp33_ASAP7_75t_L g1206 ( .A(n_461), .B(n_1207), .C(n_1208), .Y(n_1206) );
AO22x2_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_752), .B1(n_966), .B2(n_967), .Y(n_464) );
INVx1_ASAP7_75t_L g966 ( .A(n_465), .Y(n_966) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_610), .Y(n_465) );
AO22x2_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_561), .B2(n_562), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI221x1_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_490), .B1(n_492), .B2(n_504), .C(n_506), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .C(n_485), .D(n_489), .Y(n_470) );
INVx1_ASAP7_75t_L g549 ( .A(n_471), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_478), .B2(n_479), .C1(n_481), .C2(n_482), .Y(n_474) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_476), .Y(n_892) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_478), .A2(n_481), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g1492 ( .A1(n_479), .A2(n_548), .B1(n_601), .B2(n_1493), .C1(n_1494), .C2(n_1495), .Y(n_1492) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
AND2x4_ASAP7_75t_L g548 ( .A(n_483), .B(n_484), .Y(n_548) );
INVx1_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
NAND3xp33_ASAP7_75t_SL g828 ( .A(n_489), .B(n_829), .C(n_832), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g1061 ( .A(n_489), .B(n_1062), .C(n_1064), .Y(n_1061) );
NAND3xp33_ASAP7_75t_L g1105 ( .A(n_489), .B(n_1106), .C(n_1108), .Y(n_1105) );
NAND4xp25_ASAP7_75t_L g1488 ( .A(n_489), .B(n_1489), .C(n_1492), .D(n_1496), .Y(n_1488) );
OAI31xp33_ASAP7_75t_L g538 ( .A1(n_490), .A2(n_539), .A3(n_540), .B(n_549), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_490), .A2(n_828), .B(n_835), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_490), .A2(n_505), .B1(n_879), .B2(n_890), .C(n_900), .Y(n_878) );
OAI31xp33_ASAP7_75t_SL g1021 ( .A1(n_490), .A2(n_1022), .A3(n_1023), .B(n_1027), .Y(n_1021) );
OAI21xp5_ASAP7_75t_L g1060 ( .A1(n_490), .A2(n_1061), .B(n_1066), .Y(n_1060) );
OAI21xp5_ASAP7_75t_L g1104 ( .A1(n_490), .A2(n_1105), .B(n_1111), .Y(n_1104) );
OAI31xp33_ASAP7_75t_L g1169 ( .A1(n_490), .A2(n_1170), .A3(n_1171), .B(n_1173), .Y(n_1169) );
OAI31xp33_ASAP7_75t_SL g1210 ( .A1(n_490), .A2(n_1211), .A3(n_1212), .B(n_1219), .Y(n_1210) );
AOI221xp5_ASAP7_75t_L g1487 ( .A1(n_490), .A2(n_1488), .B1(n_1499), .B2(n_1508), .C(n_1509), .Y(n_1487) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
AOI31xp33_ASAP7_75t_L g598 ( .A1(n_491), .A2(n_599), .A3(n_604), .B(n_608), .Y(n_598) );
AOI31xp33_ASAP7_75t_SL g680 ( .A1(n_491), .A2(n_681), .A3(n_684), .B(n_686), .Y(n_680) );
AOI31xp33_ASAP7_75t_L g740 ( .A1(n_491), .A2(n_741), .A3(n_745), .B(n_748), .Y(n_740) );
AOI31xp33_ASAP7_75t_L g768 ( .A1(n_491), .A2(n_769), .A3(n_772), .B(n_775), .Y(n_768) );
AOI31xp33_ASAP7_75t_L g1127 ( .A1(n_491), .A2(n_1128), .A3(n_1130), .B(n_1133), .Y(n_1127) );
INVxp67_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
BUFx4f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_L g560 ( .A(n_502), .Y(n_560) );
OAI31xp33_ASAP7_75t_L g550 ( .A1(n_504), .A2(n_551), .A3(n_552), .B(n_560), .Y(n_550) );
AOI211x1_ASAP7_75t_SL g691 ( .A1(n_504), .A2(n_692), .B(n_704), .C(n_740), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g756 ( .A1(n_504), .A2(n_757), .B(n_768), .C(n_777), .Y(n_756) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g626 ( .A(n_505), .Y(n_626) );
AO211x2_ASAP7_75t_L g1113 ( .A1(n_505), .A2(n_1114), .B(n_1127), .C(n_1136), .Y(n_1113) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND3xp33_ASAP7_75t_L g537 ( .A(n_507), .B(n_538), .C(n_550), .Y(n_537) );
AND4x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .C(n_522), .D(n_529), .Y(n_507) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_SL g585 ( .A(n_518), .Y(n_585) );
INVx2_ASAP7_75t_L g903 ( .A(n_518), .Y(n_903) );
INVx2_ASAP7_75t_L g1197 ( .A(n_518), .Y(n_1197) );
INVx2_ASAP7_75t_L g1201 ( .A(n_518), .Y(n_1201) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g661 ( .A(n_519), .Y(n_661) );
INVx3_ASAP7_75t_L g783 ( .A(n_519), .Y(n_783) );
BUFx3_ASAP7_75t_L g737 ( .A(n_526), .Y(n_737) );
INVx2_ASAP7_75t_L g1093 ( .A(n_526), .Y(n_1093) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g731 ( .A(n_532), .Y(n_731) );
INVx2_ASAP7_75t_L g917 ( .A(n_532), .Y(n_917) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_543), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g1011 ( .A1(n_543), .A2(n_998), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
OAI22xp33_ASAP7_75t_L g1042 ( .A1(n_543), .A2(n_1043), .B1(n_1044), .B2(n_1045), .Y(n_1042) );
OAI22xp33_ASAP7_75t_SL g1049 ( .A1(n_543), .A2(n_845), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g1025 ( .A(n_544), .Y(n_1025) );
INVx2_ASAP7_75t_L g1215 ( .A(n_544), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_547), .A2(n_548), .B1(n_1163), .B2(n_1164), .Y(n_1172) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g823 ( .A(n_555), .Y(n_823) );
INVx2_ASAP7_75t_L g867 ( .A(n_555), .Y(n_867) );
BUFx4f_ASAP7_75t_L g873 ( .A(n_555), .Y(n_873) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OR2x2_ASAP7_75t_L g815 ( .A(n_556), .B(n_557), .Y(n_815) );
NAND4xp25_ASAP7_75t_L g879 ( .A(n_558), .B(n_880), .C(n_883), .D(n_886), .Y(n_879) );
NAND4xp25_ASAP7_75t_L g926 ( .A(n_558), .B(n_927), .C(n_930), .D(n_936), .Y(n_926) );
NAND2xp5_ASAP7_75t_SL g1017 ( .A(n_558), .B(n_1018), .Y(n_1017) );
NAND4xp25_ASAP7_75t_SL g1114 ( .A(n_558), .B(n_1115), .C(n_1118), .D(n_1121), .Y(n_1114) );
NAND3xp33_ASAP7_75t_SL g1158 ( .A(n_558), .B(n_1159), .C(n_1165), .Y(n_1158) );
NAND3xp33_ASAP7_75t_SL g1221 ( .A(n_558), .B(n_1222), .C(n_1225), .Y(n_1221) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_579), .B(n_583), .C(n_587), .D(n_593), .Y(n_578) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_582), .Y(n_601) );
INVx2_ASAP7_75t_SL g711 ( .A(n_582), .Y(n_711) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_689), .B2(n_751), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_627), .C(n_680), .Y(n_613) );
AOI31xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .A3(n_623), .B(n_626), .Y(n_614) );
INVx1_ASAP7_75t_L g1508 ( .A(n_626), .Y(n_1508) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_644), .C(n_656), .D(n_669), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_635), .C(n_642), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g1102 ( .A(n_637), .Y(n_1102) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g807 ( .A(n_639), .Y(n_807) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx2_ASAP7_75t_L g950 ( .A(n_640), .Y(n_950) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g738 ( .A(n_641), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g1150 ( .A(n_642), .B(n_1151), .C(n_1152), .Y(n_1150) );
BUFx4f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx4f_ASAP7_75t_L g739 ( .A(n_643), .Y(n_739) );
INVx4_ASAP7_75t_L g870 ( .A(n_643), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .C(n_653), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g1099 ( .A(n_647), .Y(n_1099) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g978 ( .A(n_650), .Y(n_978) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI33xp33_ASAP7_75t_L g725 ( .A1(n_653), .A2(n_726), .A3(n_730), .B1(n_733), .B2(n_736), .B3(n_739), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g1149 ( .A(n_654), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g1524 ( .A(n_654), .Y(n_1524) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_662), .C(n_665), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g853 ( .A(n_659), .Y(n_853) );
INVx1_ASAP7_75t_L g1177 ( .A(n_659), .Y(n_1177) );
BUFx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g1005 ( .A(n_661), .Y(n_1005) );
INVx1_ASAP7_75t_L g1513 ( .A(n_661), .Y(n_1513) );
BUFx3_ASAP7_75t_L g709 ( .A(n_663), .Y(n_709) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g678 ( .A(n_664), .Y(n_678) );
INVx2_ASAP7_75t_SL g786 ( .A(n_664), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_665), .B(n_789), .C(n_794), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_665), .B(n_902), .C(n_904), .Y(n_901) );
NAND3xp33_ASAP7_75t_L g1086 ( .A(n_665), .B(n_1087), .C(n_1088), .Y(n_1086) );
NAND3xp33_ASAP7_75t_L g1141 ( .A(n_665), .B(n_1142), .C(n_1144), .Y(n_1141) );
NAND3xp33_ASAP7_75t_L g1181 ( .A(n_665), .B(n_1182), .C(n_1183), .Y(n_1181) );
NAND3xp33_ASAP7_75t_L g1515 ( .A(n_665), .B(n_1516), .C(n_1517), .Y(n_1515) );
INVx5_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx6_ASAP7_75t_L g724 ( .A(n_666), .Y(n_724) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_675), .C(n_679), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g910 ( .A(n_674), .Y(n_910) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx2_ASAP7_75t_L g795 ( .A(n_678), .Y(n_795) );
INVx1_ASAP7_75t_L g913 ( .A(n_678), .Y(n_913) );
BUFx2_ASAP7_75t_L g1085 ( .A(n_679), .Y(n_1085) );
INVx1_ASAP7_75t_L g751 ( .A(n_689), .Y(n_751) );
INVx1_ASAP7_75t_L g750 ( .A(n_691), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_725), .Y(n_704) );
AOI33xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .A3(n_712), .B1(n_717), .B2(n_720), .B3(n_724), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g1510 ( .A(n_706), .B(n_1511), .C(n_1514), .Y(n_1510) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g1518 ( .A(n_711), .Y(n_1518) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g831 ( .A(n_722), .Y(n_831) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_724), .A2(n_842), .B1(n_852), .B2(n_860), .C(n_861), .Y(n_841) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_724), .A2(n_860), .B1(n_1041), .B2(n_1046), .C(n_1052), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_724), .B(n_1200), .C(n_1202), .Y(n_1199) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g1103 ( .A(n_729), .Y(n_1103) );
INVx1_ASAP7_75t_L g1523 ( .A(n_729), .Y(n_1523) );
BUFx2_ASAP7_75t_L g1507 ( .A(n_732), .Y(n_1507) );
BUFx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g1097 ( .A(n_739), .B(n_1098), .C(n_1100), .Y(n_1097) );
INVx1_ASAP7_75t_L g967 ( .A(n_752), .Y(n_967) );
AO22x2_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_875), .B1(n_876), .B2(n_965), .Y(n_752) );
INVx1_ASAP7_75t_L g965 ( .A(n_753), .Y(n_965) );
XNOR2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_809), .Y(n_753) );
INVx1_ASAP7_75t_L g808 ( .A(n_756), .Y(n_808) );
NAND4xp25_ASAP7_75t_L g777 ( .A(n_778), .B(n_788), .C(n_796), .D(n_803), .Y(n_777) );
INVx2_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g1143 ( .A(n_782), .Y(n_1143) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g793 ( .A(n_783), .Y(n_793) );
INVx1_ASAP7_75t_L g855 ( .A(n_783), .Y(n_855) );
INVx2_ASAP7_75t_L g1179 ( .A(n_783), .Y(n_1179) );
BUFx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g948 ( .A(n_799), .Y(n_948) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND3x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_827), .C(n_841), .Y(n_810) );
OR2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx2_ASAP7_75t_L g865 ( .A(n_815), .Y(n_865) );
INVx1_ASAP7_75t_L g984 ( .A(n_815), .Y(n_984) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
OAI221xp5_ASAP7_75t_L g871 ( .A1(n_830), .A2(n_833), .B1(n_864), .B2(n_872), .C(n_874), .Y(n_871) );
OR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
BUFx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g1004 ( .A(n_839), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B1(n_847), .B2(n_848), .Y(n_843) );
INVx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI22xp33_ASAP7_75t_L g997 ( .A1(n_850), .A2(n_982), .B1(n_985), .B2(n_998), .Y(n_997) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g863 ( .A1(n_857), .A2(n_859), .B1(n_864), .B2(n_866), .C(n_868), .Y(n_863) );
OAI22xp5_ASAP7_75t_SL g861 ( .A1(n_862), .A2(n_863), .B1(n_870), .B2(n_871), .Y(n_861) );
OAI33xp33_ASAP7_75t_L g975 ( .A1(n_862), .A2(n_976), .A3(n_981), .B1(n_987), .B2(n_990), .B3(n_995), .Y(n_975) );
OAI22xp5_ASAP7_75t_SL g1052 ( .A1(n_862), .A2(n_870), .B1(n_1053), .B2(n_1056), .Y(n_1052) );
INVx1_ASAP7_75t_SL g1096 ( .A(n_862), .Y(n_1096) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx2_ASAP7_75t_L g1054 ( .A(n_865), .Y(n_1054) );
OAI221xp5_ASAP7_75t_L g1053 ( .A1(n_866), .A2(n_1043), .B1(n_1045), .B2(n_1054), .C(n_1055), .Y(n_1053) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_866), .A2(n_1054), .B1(n_1057), .B2(n_1058), .C(n_1059), .Y(n_1056) );
BUFx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g991 ( .A(n_869), .Y(n_991) );
INVx1_ASAP7_75t_L g1526 ( .A(n_870), .Y(n_1526) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g986 ( .A(n_873), .Y(n_986) );
INVxp67_ASAP7_75t_SL g875 ( .A(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_923), .B1(n_924), .B2(n_964), .Y(n_876) );
INVx1_ASAP7_75t_L g964 ( .A(n_877), .Y(n_964) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_891), .B(n_895), .C(n_898), .Y(n_890) );
NAND4xp25_ASAP7_75t_L g900 ( .A(n_901), .B(n_906), .C(n_915), .D(n_920), .Y(n_900) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g963 ( .A(n_925), .Y(n_963) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_945), .Y(n_939) );
INVxp67_ASAP7_75t_SL g1231 ( .A(n_968), .Y(n_1231) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_969), .A2(n_1067), .B1(n_1068), .B2(n_1230), .Y(n_968) );
INVx1_ASAP7_75t_L g1230 ( .A(n_969), .Y(n_1230) );
XNOR2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_1028), .Y(n_969) );
INVx2_ASAP7_75t_SL g970 ( .A(n_971), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
NAND3xp33_ASAP7_75t_L g973 ( .A(n_974), .B(n_1014), .C(n_1021), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_996), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g1002 ( .A1(n_977), .A2(n_979), .B1(n_1003), .B2(n_1005), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_983), .B1(n_985), .B2(n_986), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_983), .A2(n_986), .B1(n_988), .B2(n_989), .Y(n_987) );
INVx2_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .B1(n_993), .B2(n_994), .Y(n_990) );
INVx1_ASAP7_75t_L g1522 ( .A(n_991), .Y(n_1522) );
OAI33xp33_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_1000), .A3(n_1002), .B1(n_1006), .B2(n_1010), .B3(n_1011), .Y(n_996) );
INVx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1004), .Y(n_1007) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_1005), .A2(n_1007), .B1(n_1008), .B2(n_1009), .Y(n_1006) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
XNOR2xp5_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
NAND3x1_ASAP7_75t_SL g1031 ( .A(n_1032), .B(n_1040), .C(n_1060), .Y(n_1031) );
INVxp67_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
XNOR2xp5_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1153), .Y(n_1068) );
XOR2x2_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1112), .Y(n_1069) );
NAND3x1_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1079), .C(n_1104), .Y(n_1071) );
AND4x1_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1086), .C(n_1089), .D(n_1097), .Y(n_1079) );
NAND3xp33_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1084), .C(n_1085), .Y(n_1080) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
NAND3xp33_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1091), .C(n_1096), .Y(n_1089) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx2_ASAP7_75t_SL g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
NAND4xp25_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1141), .C(n_1145), .D(n_1150), .Y(n_1136) );
NAND3xp33_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1147), .C(n_1149), .Y(n_1145) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
XOR2x2_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1192), .Y(n_1154) );
NAND3x1_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1169), .C(n_1174), .Y(n_1156) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1162), .Y(n_1224) );
AND4x1_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1181), .C(n_1184), .D(n_1189), .Y(n_1174) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
XOR2xp5_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1229), .Y(n_1192) );
NAND3xp33_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1210), .C(n_1220), .Y(n_1193) );
AND4x1_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1199), .C(n_1203), .D(n_1206), .Y(n_1194) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
OAI221xp5_ASAP7_75t_L g1232 ( .A1(n_1233), .A2(n_1482), .B1(n_1485), .B2(n_1531), .C(n_1535), .Y(n_1232) );
AOI211xp5_ASAP7_75t_L g1233 ( .A1(n_1234), .A2(n_1390), .B(n_1432), .C(n_1464), .Y(n_1233) );
NAND5xp2_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1332), .C(n_1350), .D(n_1379), .E(n_1382), .Y(n_1234) );
AOI321xp33_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1279), .A3(n_1296), .B1(n_1303), .B2(n_1311), .C(n_1322), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1275), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1262), .Y(n_1238) );
CKINVDCx6p67_ASAP7_75t_R g1278 ( .A(n_1239), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1239), .B(n_1277), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1239), .B(n_1325), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1239), .B(n_1277), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1239), .B(n_1348), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1239), .B(n_1375), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1239), .B(n_1326), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1239), .B(n_1263), .Y(n_1419) );
A2O1A1Ixp33_ASAP7_75t_SL g1468 ( .A1(n_1239), .A2(n_1469), .B(n_1473), .C(n_1475), .Y(n_1468) );
OR2x6_ASAP7_75t_SL g1239 ( .A(n_1240), .B(n_1252), .Y(n_1239) );
OAI22xp5_ASAP7_75t_L g1240 ( .A1(n_1241), .A2(n_1248), .B1(n_1249), .B2(n_1251), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1245), .Y(n_1242) );
AND2x4_ASAP7_75t_L g1250 ( .A(n_1243), .B(n_1246), .Y(n_1250) );
AND2x4_ASAP7_75t_L g1291 ( .A(n_1243), .B(n_1245), .Y(n_1291) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1244), .Y(n_1257) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1247), .B(n_1257), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_1249), .A2(n_1289), .B1(n_1290), .B2(n_1292), .Y(n_1288) );
INVx1_ASAP7_75t_SL g1249 ( .A(n_1250), .Y(n_1249) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1250), .Y(n_1302) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_1253), .A2(n_1258), .B1(n_1259), .B2(n_1261), .Y(n_1252) );
OAI22xp33_ASAP7_75t_L g1283 ( .A1(n_1253), .A2(n_1284), .B1(n_1285), .B2(n_1286), .Y(n_1283) );
OAI22xp33_ASAP7_75t_L g1306 ( .A1(n_1253), .A2(n_1259), .B1(n_1307), .B2(n_1308), .Y(n_1306) );
BUFx3_ASAP7_75t_L g1365 ( .A(n_1253), .Y(n_1365) );
BUFx6f_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_1254), .A2(n_1259), .B1(n_1273), .B2(n_1274), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1256), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1255), .B(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1255), .Y(n_1267) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1256), .Y(n_1266) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1259), .Y(n_1287) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1260), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1262), .B(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1262), .Y(n_1327) );
OAI32xp33_ASAP7_75t_L g1394 ( .A1(n_1262), .A2(n_1293), .A3(n_1333), .B1(n_1395), .B2(n_1397), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1262), .B(n_1278), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1444 ( .A(n_1262), .B(n_1337), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1271), .Y(n_1262) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1263), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1263), .B(n_1271), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1263), .B(n_1349), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1270), .Y(n_1263) );
AND2x4_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1267), .Y(n_1265) );
AND2x4_ASAP7_75t_L g1268 ( .A(n_1267), .B(n_1269), .Y(n_1268) );
HB1xp67_ASAP7_75t_L g1545 ( .A(n_1269), .Y(n_1545) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1271), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1271), .B(n_1278), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1271), .B(n_1277), .Y(n_1375) );
XNOR2xp5_ASAP7_75t_L g1486 ( .A(n_1274), .B(n_1487), .Y(n_1486) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_1275), .A2(n_1310), .B1(n_1352), .B2(n_1354), .C(n_1357), .Y(n_1351) );
O2A1O1Ixp33_ASAP7_75t_L g1413 ( .A1(n_1275), .A2(n_1377), .B(n_1414), .C(n_1415), .Y(n_1413) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
A2O1A1Ixp33_ASAP7_75t_L g1428 ( .A1(n_1276), .A2(n_1297), .B(n_1386), .C(n_1429), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1278), .B(n_1298), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1278), .B(n_1375), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1278), .B(n_1348), .Y(n_1381) );
NOR2xp33_ASAP7_75t_L g1396 ( .A(n_1278), .B(n_1298), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_1278), .B(n_1349), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1278), .B(n_1320), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1278), .B(n_1349), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1279), .B(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
OAI22xp5_ASAP7_75t_SL g1437 ( .A1(n_1280), .A2(n_1346), .B1(n_1438), .B2(n_1439), .Y(n_1437) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1293), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1281), .B(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1281), .Y(n_1316) );
INVx3_ASAP7_75t_L g1378 ( .A(n_1281), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1281), .B(n_1373), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1281), .B(n_1343), .Y(n_1424) );
AOI221xp5_ASAP7_75t_L g1441 ( .A1(n_1281), .A2(n_1442), .B1(n_1443), .B2(n_1445), .C(n_1449), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1281), .B(n_1293), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1281), .B(n_1331), .Y(n_1475) );
INVx3_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_1282), .B(n_1318), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1282), .B(n_1293), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1288), .Y(n_1282) );
HB1xp67_ASAP7_75t_L g1367 ( .A(n_1286), .Y(n_1367) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1291), .Y(n_1361) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1293), .Y(n_1310) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1293), .B(n_1305), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1293), .B(n_1305), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1293), .B(n_1340), .Y(n_1339) );
OR2x2_ASAP7_75t_L g1345 ( .A(n_1293), .B(n_1343), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1293), .B(n_1343), .Y(n_1353) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1295), .Y(n_1293) );
NOR2x1_ASAP7_75t_L g1398 ( .A(n_1296), .B(n_1399), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1296), .B(n_1313), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1296), .B(n_1385), .Y(n_1404) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1296), .B(n_1345), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1296), .B(n_1403), .Y(n_1438) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1297), .B(n_1356), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1297), .B(n_1372), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1297), .B(n_1385), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1297), .B(n_1478), .Y(n_1477) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx4_ASAP7_75t_L g1321 ( .A(n_1298), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1298), .B(n_1343), .Y(n_1342) );
OR2x2_ASAP7_75t_L g1393 ( .A(n_1298), .B(n_1326), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1298), .B(n_1373), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_1298), .B(n_1372), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1298), .B(n_1347), .Y(n_1467) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1298), .B(n_1389), .Y(n_1474) );
AND2x6_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1300), .Y(n_1298) );
INVx2_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
OAI22xp5_ASAP7_75t_L g1359 ( .A1(n_1302), .A2(n_1360), .B1(n_1361), .B2(n_1362), .Y(n_1359) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1303), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1309), .Y(n_1303) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1304), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1304), .B(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1304), .Y(n_1446) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1304), .Y(n_1463) );
HB1xp67_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1343 ( .A(n_1305), .Y(n_1343) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1310), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1314), .B1(n_1316), .B2(n_1319), .Y(n_1311) );
INVxp67_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1313), .B(n_1321), .Y(n_1411) );
INVxp67_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1317), .Y(n_1315) );
AOI21xp5_ASAP7_75t_L g1427 ( .A1(n_1316), .A2(n_1335), .B(n_1357), .Y(n_1427) );
AOI22xp5_ASAP7_75t_L g1453 ( .A1(n_1316), .A2(n_1454), .B1(n_1457), .B2(n_1461), .Y(n_1453) );
OAI211xp5_ASAP7_75t_L g1390 ( .A1(n_1317), .A2(n_1391), .B(n_1402), .C(n_1416), .Y(n_1390) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVxp67_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1321), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1321), .B(n_1353), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1321), .B(n_1381), .Y(n_1380) );
AOI21xp5_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1327), .B(n_1328), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1323), .B(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
OAI31xp33_ASAP7_75t_L g1476 ( .A1(n_1324), .A2(n_1355), .A3(n_1477), .B(n_1479), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1325), .B(n_1337), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1325), .B(n_1396), .Y(n_1448) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1331), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1330), .B(n_1419), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1330), .B(n_1348), .Y(n_1429) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1331), .Y(n_1431) );
AOI211xp5_ASAP7_75t_SL g1332 ( .A1(n_1333), .A2(n_1335), .B(n_1338), .C(n_1344), .Y(n_1332) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_1333), .A2(n_1418), .B1(n_1420), .B2(n_1421), .Y(n_1417) );
AOI21xp5_ASAP7_75t_L g1433 ( .A1(n_1333), .A2(n_1434), .B(n_1437), .Y(n_1433) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1335), .B(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1336), .B(n_1463), .Y(n_1462) );
INVxp67_ASAP7_75t_SL g1338 ( .A(n_1339), .Y(n_1338) );
INVxp33_ASAP7_75t_L g1450 ( .A(n_1340), .Y(n_1450) );
NOR2xp33_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1342), .Y(n_1340) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1341), .Y(n_1478) );
INVx2_ASAP7_75t_SL g1373 ( .A(n_1343), .Y(n_1373) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1346), .Y(n_1344) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1345), .Y(n_1403) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
OAI21xp33_ASAP7_75t_SL g1410 ( .A1(n_1347), .A2(n_1411), .B(n_1412), .Y(n_1410) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1348), .Y(n_1471) );
OAI21xp5_ASAP7_75t_L g1350 ( .A1(n_1351), .A2(n_1368), .B(n_1376), .Y(n_1350) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1353), .Y(n_1420) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVxp67_ASAP7_75t_L g1421 ( .A(n_1356), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1357), .B(n_1377), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_1358), .Y(n_1357) );
OR2x6_ASAP7_75t_SL g1358 ( .A(n_1359), .B(n_1363), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1365), .B1(n_1366), .B2(n_1367), .Y(n_1363) );
BUFx2_ASAP7_75t_SL g1484 ( .A(n_1367), .Y(n_1484) );
INVxp67_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1374), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
AOI221xp5_ASAP7_75t_L g1391 ( .A1(n_1373), .A2(n_1378), .B1(n_1392), .B2(n_1394), .C(n_1400), .Y(n_1391) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_1373), .B(n_1401), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1373), .B(n_1393), .Y(n_1409) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1373), .Y(n_1481) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1375), .Y(n_1472) );
AOI211xp5_ASAP7_75t_L g1416 ( .A1(n_1377), .A2(n_1417), .B(n_1422), .C(n_1430), .Y(n_1416) );
NOR2xp33_ASAP7_75t_L g1459 ( .A(n_1377), .B(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_SL g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1381), .Y(n_1456) );
AOI21xp5_ASAP7_75t_L g1382 ( .A1(n_1383), .A2(n_1386), .B(n_1387), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
NOR2xp33_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1389), .Y(n_1387) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1388), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g1430 ( .A(n_1389), .B(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
AOI211xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1404), .B(n_1405), .C(n_1413), .Y(n_1402) );
OAI21xp33_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1408), .B(n_1410), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVxp67_ASAP7_75t_SL g1408 ( .A(n_1409), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1415), .B(n_1458), .Y(n_1457) );
OAI211xp5_ASAP7_75t_L g1422 ( .A1(n_1423), .A2(n_1425), .B(n_1427), .C(n_1428), .Y(n_1422) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
AOI21xp33_ASAP7_75t_SL g1449 ( .A1(n_1425), .A2(n_1450), .B(n_1451), .Y(n_1449) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
NAND3xp33_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1441), .C(n_1453), .Y(n_1432) );
INVxp67_ASAP7_75t_SL g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1447), .Y(n_1445) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVxp67_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
INVxp67_ASAP7_75t_SL g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
OAI211xp5_ASAP7_75t_L g1464 ( .A1(n_1465), .A2(n_1467), .B(n_1468), .C(n_1476), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1466), .B(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1472), .Y(n_1470) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
CKINVDCx5p33_ASAP7_75t_R g1482 ( .A(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_SL g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
HB1xp67_ASAP7_75t_L g1542 ( .A(n_1487), .Y(n_1542) );
NAND4xp25_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1515), .C(n_1519), .D(n_1525), .Y(n_1509) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
NAND3xp33_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1521), .C(n_1524), .Y(n_1519) );
NAND3xp33_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1527), .C(n_1530), .Y(n_1525) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx2_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx2_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
CKINVDCx5p33_ASAP7_75t_R g1537 ( .A(n_1538), .Y(n_1537) );
OAI21xp5_ASAP7_75t_L g1544 ( .A1(n_1539), .A2(n_1545), .B(n_1546), .Y(n_1544) );
INVxp33_ASAP7_75t_SL g1540 ( .A(n_1541), .Y(n_1540) );
BUFx2_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
endmodule