module real_jpeg_29940_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_1),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_1),
.A2(n_25),
.B1(n_58),
.B2(n_62),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_1),
.A2(n_25),
.B1(n_49),
.B2(n_50),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_52),
.B1(n_58),
.B2(n_62),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_6),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_6),
.A2(n_30),
.B(n_34),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_6),
.A2(n_26),
.B1(n_28),
.B2(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_6),
.B(n_32),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_6),
.A2(n_49),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_6),
.B(n_49),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_6),
.B(n_53),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_6),
.A2(n_56),
.B1(n_223),
.B2(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_6),
.A2(n_33),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_26),
.B1(n_28),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_7),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_96),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_7),
.A2(n_58),
.B1(n_62),
.B2(n_96),
.Y(n_217)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_9),
.A2(n_58),
.B1(n_62),
.B2(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_10),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_10),
.A2(n_37),
.B1(n_58),
.B2(n_62),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_26),
.B1(n_28),
.B2(n_40),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_11),
.A2(n_40),
.B1(n_58),
.B2(n_62),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_12),
.A2(n_58),
.B1(n_62),
.B2(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_72),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_12),
.A2(n_49),
.A3(n_62),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_13),
.A2(n_58),
.B1(n_62),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_67),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_16),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_17),
.A2(n_26),
.B1(n_28),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_17),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_133),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_17),
.A2(n_49),
.B1(n_50),
.B2(n_133),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_17),
.A2(n_58),
.B1(n_62),
.B2(n_133),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_99),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_21),
.B(n_99),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_76),
.C(n_86),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_22),
.B(n_76),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_22),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_38),
.CI(n_54),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_38),
.C(n_54),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_26),
.A2(n_35),
.B(n_137),
.C(n_138),
.Y(n_136)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_29),
.A2(n_32),
.B1(n_132),
.B2(n_162),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_32),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_43),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_33),
.A2(n_47),
.A3(n_50),
.B1(n_240),
.B2(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_34),
.B(n_137),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_36),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_51),
.B2(n_53),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_39),
.A2(n_41),
.B1(n_53),
.B2(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_41),
.A2(n_53),
.B1(n_160),
.B2(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_46),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_42),
.A2(n_46),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_42),
.A2(n_46),
.B1(n_143),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_42),
.A2(n_46),
.B1(n_180),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_47),
.Y(n_249)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_49),
.B(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_68),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_55),
.B(n_68),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_63),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_60),
.B1(n_65),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_56),
.A2(n_65),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_56),
.A2(n_65),
.B1(n_217),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_56),
.A2(n_212),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_57),
.A2(n_90),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_57),
.A2(n_64),
.B1(n_140),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_57),
.A2(n_64),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_58),
.B(n_72),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_58),
.B(n_229),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g251 ( 
.A(n_64),
.Y(n_251)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_65),
.B(n_137),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_71),
.B1(n_82),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_70),
.A2(n_71),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_70),
.A2(n_71),
.B1(n_198),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_70),
.A2(n_71),
.B1(n_165),
.B2(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_71),
.B(n_137),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_85),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_80),
.A2(n_83),
.B1(n_93),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_80),
.A2(n_83),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_85),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.C(n_97),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_91),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_97),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_98),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_120),
.B2(n_121),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B(n_108),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_106),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_116),
.B1(n_131),
.B2(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_120),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_148),
.B(n_276),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_146),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_126),
.B(n_146),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.C(n_145),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_145),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.C(n_142),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_142),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_139),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_185),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_168),
.B(n_184),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_166),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_166),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_156),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_156),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.C(n_163),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_172),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_175),
.Y(n_274)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_178),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_181),
.B(n_183),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_182),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.C(n_188),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_270),
.B(n_275),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_256),
.B(n_269),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_233),
.B(n_255),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_213),
.B(n_232),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_203),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_193),
.B(n_203),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_208),
.C(n_210),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_220),
.B(n_231),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_219),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_225),
.B(n_230),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_235),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_246),
.B1(n_253),
.B2(n_254),
.Y(n_235)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_241),
.B1(n_244),
.B2(n_245),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_245),
.C(n_254),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_246),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_258),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_265),
.C(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);


endmodule