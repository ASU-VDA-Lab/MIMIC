module fake_jpeg_18608_n_143 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_29),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_11),
.B(n_20),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_21),
.B1(n_17),
.B2(n_11),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_47),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_48),
.B1(n_50),
.B2(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_38),
.Y(n_47)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_12),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_48),
.B(n_45),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_50),
.B(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_50),
.B1(n_58),
.B2(n_48),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_83),
.B1(n_72),
.B2(n_67),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_58),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_81),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_56),
.B(n_63),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_20),
.B(n_18),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_84),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_56),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_71),
.B(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_71),
.Y(n_88)
);

OA21x2_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_16),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_23),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_7),
.B(n_1),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_66),
.B(n_51),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_32),
.B(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_43),
.B1(n_65),
.B2(n_35),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_97),
.B1(n_37),
.B2(n_23),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_32),
.C(n_35),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_49),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_32),
.B1(n_35),
.B2(n_64),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_37),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_103),
.B(n_22),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_105),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_17),
.B(n_16),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_94),
.Y(n_112)
);

AOI31xp67_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_110),
.A3(n_7),
.B(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_113),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_114),
.B(n_116),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_119),
.B(n_0),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_87),
.B1(n_2),
.B2(n_3),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_87),
.C(n_22),
.Y(n_119)
);

AOI211xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_103),
.B(n_100),
.C(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_119),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_4),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_2),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_2),
.B(n_4),
.C(n_6),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_6),
.B(n_8),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_113),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_4),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_6),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.C(n_15),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_120),
.C(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.C(n_8),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_120),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_128),
.B(n_8),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_9),
.B(n_139),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_137),
.C(n_134),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);


endmodule