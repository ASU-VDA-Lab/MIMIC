module fake_ariane_2804_n_2931 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2931);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2931;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_2238;
wire n_1503;
wire n_764;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2391;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_661;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_1253;
wire n_1468;
wire n_762;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_1623;
wire n_990;
wire n_1903;
wire n_2147;
wire n_867;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_1832;
wire n_767;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_1914;
wire n_965;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_1689;
wire n_970;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_590;
wire n_2075;
wire n_699;
wire n_727;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2774;
wire n_2707;
wire n_2754;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_710;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_1700;
wire n_862;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_642;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_1118;
wire n_943;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_756;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_807;
wire n_891;
wire n_1659;
wire n_885;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_820;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_1809;
wire n_765;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2556;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_2351;
wire n_1619;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_2206;
wire n_635;
wire n_997;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2917;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1477;
wire n_1777;
wire n_1019;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1983;
wire n_1273;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2869;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_803;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g584 ( 
.A(n_159),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_283),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_427),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_281),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_581),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_545),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_188),
.Y(n_590)
);

BUFx5_ASAP7_75t_L g591 ( 
.A(n_320),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_35),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_103),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_521),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_292),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_405),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_486),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_136),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_230),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_404),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_170),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_515),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_1),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_343),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_149),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_497),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_502),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_536),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_305),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_86),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_458),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_437),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_144),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_260),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_299),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_538),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_244),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_453),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_416),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_284),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_154),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_111),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_354),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_34),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_232),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_102),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_512),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_438),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_567),
.Y(n_630)
);

CKINVDCx16_ASAP7_75t_R g631 ( 
.A(n_97),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_516),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_251),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_421),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_559),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_298),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_231),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_484),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_143),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_271),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_503),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_296),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_273),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_109),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_65),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_191),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_234),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_388),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_1),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_11),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_182),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_443),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_436),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_336),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_555),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_25),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_365),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_246),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_363),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_480),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_57),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_426),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_277),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_552),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_299),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_349),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_386),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_19),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_16),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_396),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_52),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_85),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_249),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_460),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_429),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_259),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_467),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_482),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_523),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_532),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_471),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_366),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_504),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_501),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_553),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_120),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_556),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_39),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_289),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_148),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_471),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_57),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_540),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_528),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_514),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_159),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_216),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_125),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_184),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_157),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_305),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_439),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_466),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_297),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_399),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_274),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_566),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_52),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_268),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_180),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_550),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_335),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_439),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_465),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_5),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_539),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_312),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_527),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_335),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_108),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_227),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_255),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_525),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_338),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_3),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_524),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_482),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_580),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_522),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_360),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_81),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_73),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_513),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_385),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_308),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_564),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_579),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_163),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_517),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_87),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_201),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_96),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_219),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_133),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_36),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_68),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_201),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_498),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_88),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_547),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_93),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_535),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_370),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_199),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_563),
.Y(n_756)
);

BUFx10_ASAP7_75t_L g757 ( 
.A(n_369),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_245),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_62),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_39),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_565),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_156),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_40),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_533),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_300),
.Y(n_765)
);

BUFx2_ASAP7_75t_SL g766 ( 
.A(n_24),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_98),
.Y(n_767)
);

BUFx5_ASAP7_75t_L g768 ( 
.A(n_223),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_390),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_190),
.Y(n_770)
);

CKINVDCx16_ASAP7_75t_R g771 ( 
.A(n_334),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_106),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_281),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_583),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_120),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_290),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_344),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_195),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_106),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_317),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_17),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_521),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_494),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_372),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_570),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_354),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_19),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_379),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_172),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_389),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_294),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_226),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_473),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_326),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_275),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_560),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_375),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_124),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_414),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_59),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_209),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_390),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_531),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_549),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_575),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_228),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_546),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_132),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_383),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_358),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_129),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_127),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_537),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_530),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_513),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_499),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_508),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_139),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_407),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_140),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_423),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_526),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_72),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_561),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_353),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_222),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_573),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_415),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_392),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_548),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_495),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_520),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_243),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_503),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_519),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_98),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_541),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_89),
.Y(n_838)
);

INVxp33_ASAP7_75t_R g839 ( 
.A(n_475),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_453),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_222),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_442),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_465),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_343),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_569),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_26),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_293),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_100),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_383),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_496),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_278),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_554),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_130),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_388),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_60),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_568),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_71),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_71),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_249),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_313),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_582),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_458),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_493),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_282),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_23),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_22),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_358),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_315),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_235),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_507),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_511),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_576),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_101),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_199),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_22),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_352),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_186),
.Y(n_877)
);

BUFx10_ASAP7_75t_L g878 ( 
.A(n_141),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_534),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_316),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_356),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_208),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_14),
.Y(n_883)
);

CKINVDCx14_ASAP7_75t_R g884 ( 
.A(n_82),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_455),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_61),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_90),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_14),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_165),
.Y(n_889)
);

BUFx10_ASAP7_75t_L g890 ( 
.A(n_543),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_328),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_152),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_261),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_264),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_510),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_256),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_209),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_455),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_303),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_280),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_258),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_276),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_94),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_142),
.Y(n_904)
);

BUFx8_ASAP7_75t_SL g905 ( 
.A(n_180),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_416),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_551),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_104),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_190),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_84),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_526),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_54),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_341),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_200),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_284),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_577),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_370),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_542),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_463),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_514),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_248),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_224),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_55),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_440),
.Y(n_924)
);

BUFx10_ASAP7_75t_L g925 ( 
.A(n_463),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_123),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_518),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_280),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_49),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_423),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_145),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_20),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_449),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_194),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_378),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_373),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_485),
.Y(n_937)
);

BUFx10_ASAP7_75t_L g938 ( 
.A(n_499),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_529),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_419),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_345),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_519),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_457),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_183),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_192),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_574),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_359),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_386),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_376),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_558),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_456),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_33),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_242),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_294),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_172),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_137),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_324),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_510),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_45),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_35),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_422),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_572),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_181),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_230),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_56),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_257),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_55),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_366),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_505),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_509),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_404),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_481),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_103),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_91),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_112),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_36),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_101),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_210),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_121),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_506),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_377),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_169),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_202),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_418),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_467),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_361),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_204),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_102),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_34),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_375),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_117),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_523),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_578),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_289),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_412),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_496),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_162),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_219),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_328),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_188),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_270),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_544),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_557),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_352),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_223),
.Y(n_1005)
);

BUFx8_ASAP7_75t_SL g1006 ( 
.A(n_500),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_278),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_38),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_95),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_112),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_100),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_137),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_9),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_77),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_408),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_31),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_82),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_571),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_480),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_117),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_293),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_473),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_591),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_591),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_591),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_784),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_784),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_659),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_905),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_591),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_591),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_591),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_591),
.Y(n_1033)
);

INVxp33_ASAP7_75t_L g1034 ( 
.A(n_598),
.Y(n_1034)
);

INVxp67_ASAP7_75t_SL g1035 ( 
.A(n_1001),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_591),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_768),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_768),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_768),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_884),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_768),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_768),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_768),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_1006),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_1001),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_659),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_768),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_768),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_665),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_665),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_688),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_631),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_671),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_688),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_708),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_771),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_951),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_632),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_708),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_632),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_737),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_737),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_879),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_671),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_786),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_589),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_761),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_879),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_761),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_630),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_814),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_786),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_814),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_822),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_824),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_824),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_827),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_822),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_632),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_827),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_830),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_830),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_852),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_632),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_632),
.Y(n_1085)
);

CKINVDCx16_ASAP7_75t_R g1086 ( 
.A(n_785),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_852),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_700),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_872),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_918),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_637),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_950),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_602),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_872),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_907),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_907),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_980),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_1052),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1023),
.Y(n_1099)
);

OAI22x1_ASAP7_75t_L g1100 ( 
.A1(n_1078),
.A2(n_980),
.B1(n_683),
.B2(n_895),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_1048),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1048),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1023),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1058),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1053),
.A2(n_640),
.B1(n_668),
.B2(n_628),
.Y(n_1105)
);

CKINVDCx11_ASAP7_75t_R g1106 ( 
.A(n_1093),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1024),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1058),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1060),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1060),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1064),
.A2(n_696),
.B1(n_719),
.B2(n_679),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1024),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1079),
.B(n_916),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1025),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_1085),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1028),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1085),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_1025),
.A2(n_1018),
.B(n_993),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1088),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1088),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1030),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_SL g1122 ( 
.A1(n_1029),
.A2(n_742),
.B1(n_773),
.B2(n_731),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1084),
.B(n_916),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1030),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1031),
.Y(n_1125)
);

OAI22x1_ASAP7_75t_R g1126 ( 
.A1(n_1044),
.A2(n_835),
.B1(n_848),
.B2(n_791),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_1049),
.B(n_672),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1031),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1032),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1032),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1049),
.B(n_650),
.Y(n_1131)
);

OAI22x1_ASAP7_75t_R g1132 ( 
.A1(n_1066),
.A2(n_849),
.B1(n_896),
.B2(n_889),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1070),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1033),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1033),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1036),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1036),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1050),
.B(n_650),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1065),
.A2(n_899),
.B1(n_906),
.B2(n_897),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1037),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1037),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1038),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1050),
.B(n_720),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1038),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1039),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_1063),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1026),
.B(n_1027),
.Y(n_1147)
);

OAI22x1_ASAP7_75t_SL g1148 ( 
.A1(n_1056),
.A2(n_915),
.B1(n_947),
.B2(n_920),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1078),
.A2(n_998),
.B1(n_958),
.B2(n_1020),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1090),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1039),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1057),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1041),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_1041),
.A2(n_1018),
.B(n_993),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1042),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1042),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1043),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1043),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1047),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1125),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_1106),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1133),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1133),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1150),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1102),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1150),
.Y(n_1166)
);

AND3x2_ASAP7_75t_L g1167 ( 
.A(n_1098),
.B(n_1097),
.C(n_739),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1106),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1098),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1098),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1102),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_1146),
.B(n_1051),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1152),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_R g1174 ( 
.A(n_1152),
.B(n_1092),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1152),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1148),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1148),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1146),
.B(n_1035),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1122),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1122),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_1101),
.B(n_1086),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1125),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1147),
.B(n_1091),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1125),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1102),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1105),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1121),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_R g1188 ( 
.A(n_1101),
.B(n_1040),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1105),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1128),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1128),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_R g1192 ( 
.A(n_1101),
.B(n_1072),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1132),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1128),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1130),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1130),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1130),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_R g1198 ( 
.A(n_1147),
.B(n_1097),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_1132),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_SL g1200 ( 
.A(n_1127),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1134),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1111),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1149),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1134),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1116),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_R g1206 ( 
.A(n_1101),
.B(n_1129),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1134),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1111),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1116),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1136),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1139),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1139),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1136),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1149),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1121),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1146),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1146),
.Y(n_1217)
);

AND2x6_ASAP7_75t_L g1218 ( 
.A(n_1178),
.B(n_1190),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1165),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1165),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1171),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1191),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1195),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1171),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1183),
.B(n_1131),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1185),
.Y(n_1226)
);

NOR3xp33_ASAP7_75t_L g1227 ( 
.A(n_1163),
.B(n_732),
.C(n_645),
.Y(n_1227)
);

INVxp33_ASAP7_75t_SL g1228 ( 
.A(n_1163),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1178),
.B(n_1127),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1178),
.B(n_1127),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1190),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1187),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1196),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1209),
.B(n_1131),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1185),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1201),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1170),
.A2(n_1068),
.B1(n_1063),
.B2(n_1100),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1187),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1213),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1187),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1194),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1194),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1200),
.A2(n_1100),
.B1(n_1068),
.B2(n_1127),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1205),
.B(n_1146),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1197),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1173),
.B(n_1146),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1197),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1204),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1204),
.Y(n_1249)
);

NOR3xp33_ASAP7_75t_L g1250 ( 
.A(n_1164),
.B(n_840),
.C(n_794),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1160),
.B(n_1146),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1200),
.A2(n_1100),
.B1(n_1127),
.B2(n_1034),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1207),
.Y(n_1253)
);

NOR2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1170),
.B(n_1045),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1182),
.A2(n_1142),
.B(n_1136),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1175),
.A2(n_585),
.B1(n_596),
.B2(n_593),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1207),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1210),
.B(n_1099),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1210),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1192),
.B(n_1131),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1174),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1184),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1187),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1162),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_L g1265 ( 
.A(n_1187),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1215),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1215),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1215),
.B(n_1099),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1215),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1215),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1169),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1206),
.Y(n_1272)
);

AND2x6_ASAP7_75t_L g1273 ( 
.A(n_1200),
.B(n_1138),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1216),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1181),
.B(n_1146),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1172),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1216),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1164),
.B(n_1113),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1217),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1167),
.B(n_1138),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1217),
.B(n_1103),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1166),
.B(n_1046),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1188),
.B(n_1103),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1166),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1214),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1186),
.B(n_1138),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1189),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1212),
.Y(n_1288)
);

AND2x2_ASAP7_75t_SL g1289 ( 
.A(n_1198),
.B(n_1154),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1189),
.B(n_1113),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1212),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1161),
.Y(n_1292)
);

AND2x2_ASAP7_75t_SL g1293 ( 
.A(n_1202),
.B(n_1118),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1202),
.B(n_1123),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1208),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1294),
.B(n_1290),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1225),
.B(n_1123),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1285),
.B(n_1208),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1231),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1225),
.B(n_1260),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1260),
.B(n_1143),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1265),
.B(n_1129),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1218),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1254),
.A2(n_1211),
.B1(n_1203),
.B2(n_1143),
.Y(n_1304)
);

NAND2xp33_ASAP7_75t_L g1305 ( 
.A(n_1232),
.B(n_1129),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1271),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1268),
.A2(n_1112),
.B(n_1107),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1284),
.A2(n_1211),
.B1(n_595),
.B2(n_687),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1271),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_L g1310 ( 
.A(n_1282),
.B(n_1168),
.C(n_973),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1228),
.A2(n_1193),
.B1(n_1199),
.B2(n_1168),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1222),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1231),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1231),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1222),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1286),
.B(n_1143),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1223),
.Y(n_1317)
);

AND2x2_ASAP7_75t_SL g1318 ( 
.A(n_1289),
.B(n_1118),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1231),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1286),
.B(n_1129),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1219),
.Y(n_1321)
);

NOR2x2_ASAP7_75t_L g1322 ( 
.A(n_1285),
.B(n_1126),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1223),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1289),
.A2(n_1054),
.B1(n_1055),
.B2(n_1051),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1284),
.A2(n_707),
.B1(n_713),
.B2(n_584),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1265),
.B(n_1129),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1229),
.B(n_1137),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1289),
.A2(n_1055),
.B1(n_1059),
.B2(n_1054),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1233),
.A2(n_1061),
.B(n_1062),
.C(n_1059),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1229),
.B(n_1137),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1229),
.B(n_1137),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1249),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1229),
.B(n_1137),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1285),
.B(n_839),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1233),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1278),
.B(n_1137),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1230),
.B(n_1107),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1288),
.B(n_1061),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1230),
.B(n_1112),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1284),
.B(n_1114),
.Y(n_1340)
);

INVx8_ASAP7_75t_L g1341 ( 
.A(n_1273),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_L g1342 ( 
.A(n_1232),
.B(n_1114),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1265),
.B(n_1144),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1284),
.B(n_1124),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1265),
.B(n_1144),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1249),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1288),
.B(n_1124),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1232),
.B(n_1155),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1288),
.B(n_1074),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1288),
.B(n_1135),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1230),
.B(n_1135),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1236),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1232),
.B(n_1155),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1291),
.B(n_1287),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1230),
.B(n_1140),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1232),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1236),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1239),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1239),
.Y(n_1359)
);

NOR2xp67_ASAP7_75t_L g1360 ( 
.A(n_1264),
.B(n_1176),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1291),
.B(n_1140),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1232),
.B(n_1157),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1291),
.B(n_1177),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1249),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1262),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_SL g1366 ( 
.A(n_1280),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1249),
.Y(n_1367)
);

AO221x1_ASAP7_75t_L g1368 ( 
.A1(n_1237),
.A2(n_1256),
.B1(n_1291),
.B2(n_1261),
.C(n_1272),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1272),
.B(n_1157),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1263),
.B(n_1159),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1261),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1262),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1219),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1283),
.B(n_1159),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1263),
.B(n_1142),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1283),
.B(n_1142),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1219),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1234),
.B(n_637),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1262),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1220),
.Y(n_1380)
);

O2A1O1Ixp5_ASAP7_75t_L g1381 ( 
.A1(n_1281),
.A2(n_1151),
.B(n_1158),
.C(n_1145),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1234),
.B(n_1145),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1220),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1287),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1220),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1295),
.B(n_1145),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1241),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1241),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1293),
.A2(n_1067),
.B1(n_1069),
.B2(n_1062),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1295),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1247),
.Y(n_1391)
);

AND2x2_ASAP7_75t_SL g1392 ( 
.A(n_1293),
.B(n_1118),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1293),
.A2(n_1069),
.B1(n_1071),
.B2(n_1067),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1221),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1273),
.B(n_1151),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1254),
.A2(n_722),
.B1(n_745),
.B2(n_735),
.Y(n_1396)
);

OAI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1256),
.A2(n_819),
.B1(n_1005),
.B2(n_994),
.C(n_919),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1273),
.B(n_1151),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1312),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1340),
.A2(n_1281),
.B(n_1268),
.Y(n_1400)
);

BUFx4f_ASAP7_75t_L g1401 ( 
.A(n_1371),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1381),
.A2(n_1258),
.B(n_1247),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1325),
.A2(n_1250),
.B(n_1227),
.C(n_683),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1340),
.A2(n_1258),
.B(n_1263),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1300),
.B(n_1243),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1296),
.B(n_1252),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1347),
.B(n_1273),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1347),
.B(n_1273),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1338),
.B(n_1273),
.Y(n_1409)
);

AND2x2_ASAP7_75t_SL g1410 ( 
.A(n_1389),
.B(n_1393),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1315),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1350),
.B(n_1273),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1324),
.A2(n_1274),
.B1(n_1279),
.B2(n_1277),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1344),
.A2(n_1270),
.B(n_1263),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1356),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1303),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_SL g1417 ( 
.A(n_1311),
.B(n_1292),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1324),
.A2(n_1274),
.B1(n_1279),
.B2(n_1277),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1303),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1350),
.A2(n_1244),
.B(n_1279),
.C(n_1277),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_R g1421 ( 
.A(n_1349),
.B(n_1292),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1328),
.A2(n_1274),
.B1(n_1240),
.B2(n_1266),
.Y(n_1422)
);

O2A1O1Ixp5_ASAP7_75t_L g1423 ( 
.A1(n_1344),
.A2(n_1246),
.B(n_1240),
.C(n_1238),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1306),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1296),
.B(n_1280),
.Y(n_1425)
);

OAI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1361),
.A2(n_587),
.B(n_586),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1310),
.B(n_1276),
.C(n_1073),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1297),
.B(n_1273),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1361),
.A2(n_1245),
.B(n_1242),
.Y(n_1429)
);

AO21x1_ASAP7_75t_L g1430 ( 
.A1(n_1386),
.A2(n_1269),
.B(n_1267),
.Y(n_1430)
);

BUFx4f_ASAP7_75t_L g1431 ( 
.A(n_1354),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1338),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1305),
.A2(n_1270),
.B(n_1263),
.Y(n_1433)
);

BUFx4f_ASAP7_75t_L g1434 ( 
.A(n_1363),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1308),
.A2(n_1280),
.B1(n_1218),
.B2(n_1274),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1321),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1321),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1298),
.B(n_1280),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1385),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1385),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1298),
.B(n_1301),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1309),
.B(n_1267),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1341),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1342),
.A2(n_1270),
.B(n_1263),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1317),
.Y(n_1445)
);

OAI21xp33_ASAP7_75t_L g1446 ( 
.A1(n_1320),
.A2(n_592),
.B(n_590),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1389),
.B(n_1218),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1341),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1323),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1307),
.A2(n_1245),
.B(n_1242),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1365),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1372),
.Y(n_1452)
);

AO21x1_ASAP7_75t_L g1453 ( 
.A1(n_1386),
.A2(n_1375),
.B(n_1353),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1375),
.A2(n_1270),
.B(n_1269),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1343),
.A2(n_1270),
.B(n_1251),
.Y(n_1455)
);

OAI321xp33_ASAP7_75t_L g1456 ( 
.A1(n_1397),
.A2(n_932),
.A3(n_873),
.B1(n_967),
.B2(n_895),
.C(n_672),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1322),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1393),
.B(n_1335),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1379),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1334),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1384),
.B(n_1218),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1390),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1316),
.B(n_1242),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1352),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1357),
.B(n_1218),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1373),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1343),
.A2(n_1270),
.B(n_1240),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1328),
.A2(n_1240),
.B1(n_1266),
.B2(n_1238),
.Y(n_1468)
);

OAI21xp33_ASAP7_75t_L g1469 ( 
.A1(n_1336),
.A2(n_600),
.B(n_594),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1470)
);

AO21x1_ASAP7_75t_L g1471 ( 
.A1(n_1348),
.A2(n_1266),
.B(n_1238),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1345),
.A2(n_1266),
.B(n_1238),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1377),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1337),
.A2(n_593),
.B1(n_596),
.B2(n_585),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1345),
.A2(n_1255),
.B(n_1248),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1380),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1378),
.B(n_1218),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1304),
.B(n_637),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1382),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1387),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1302),
.A2(n_1255),
.B(n_1248),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1302),
.A2(n_1255),
.B(n_1248),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1388),
.Y(n_1483)
);

CKINVDCx10_ASAP7_75t_R g1484 ( 
.A(n_1366),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1374),
.B(n_1218),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1326),
.A2(n_1255),
.B(n_1253),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1326),
.A2(n_1253),
.B(n_1245),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1369),
.A2(n_1257),
.B(n_1253),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1383),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1348),
.A2(n_1259),
.B(n_1257),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1353),
.A2(n_1259),
.B(n_1257),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1360),
.B(n_1276),
.Y(n_1492)
);

BUFx4f_ASAP7_75t_L g1493 ( 
.A(n_1341),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1368),
.B(n_1334),
.Y(n_1494)
);

AOI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1392),
.A2(n_1259),
.B(n_1073),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1336),
.A2(n_1075),
.B(n_1076),
.C(n_1071),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1410),
.A2(n_1396),
.B1(n_1392),
.B2(n_1366),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1400),
.A2(n_1356),
.B(n_1318),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1481),
.A2(n_1398),
.B(n_1395),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1424),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1441),
.A2(n_1425),
.B(n_1494),
.C(n_1403),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1404),
.A2(n_1356),
.B(n_1318),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1420),
.A2(n_1351),
.B(n_1339),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_L g1504 ( 
.A(n_1438),
.Y(n_1504)
);

O2A1O1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1462),
.A2(n_1329),
.B(n_932),
.C(n_967),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1406),
.B(n_1391),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1460),
.B(n_1179),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1414),
.A2(n_1356),
.B(n_1362),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1405),
.A2(n_1355),
.B1(n_1218),
.B2(n_1327),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1451),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1417),
.A2(n_1330),
.B1(n_1333),
.B2(n_1331),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1401),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1431),
.B(n_1376),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1431),
.B(n_1421),
.Y(n_1514)
);

NOR3xp33_ASAP7_75t_L g1515 ( 
.A(n_1427),
.B(n_873),
.C(n_599),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1407),
.A2(n_1370),
.B(n_1362),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1479),
.B(n_1329),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1401),
.B(n_1180),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1426),
.A2(n_1076),
.B(n_1077),
.C(n_1075),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1457),
.B(n_1299),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1399),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1432),
.B(n_1394),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1411),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1407),
.A2(n_1370),
.B(n_1314),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1434),
.B(n_1313),
.Y(n_1525)
);

OAI22x1_ASAP7_75t_L g1526 ( 
.A1(n_1478),
.A2(n_1126),
.B1(n_599),
.B2(n_604),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1463),
.A2(n_1080),
.B(n_1081),
.C(n_1077),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1435),
.A2(n_604),
.B1(n_607),
.B2(n_597),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1445),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1408),
.A2(n_1412),
.B(n_1433),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1447),
.A2(n_624),
.B1(n_647),
.B2(n_616),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1449),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1415),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1469),
.A2(n_1081),
.B(n_1082),
.C(n_1080),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1434),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1415),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1470),
.B(n_1364),
.Y(n_1537)
);

CKINVDCx14_ASAP7_75t_R g1538 ( 
.A(n_1484),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1464),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1493),
.B(n_1319),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1415),
.Y(n_1541)
);

AOI21x1_ASAP7_75t_SL g1542 ( 
.A1(n_1470),
.A2(n_766),
.B(n_603),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1408),
.A2(n_1346),
.B(n_1332),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1412),
.A2(n_1367),
.B1(n_766),
.B2(n_605),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1442),
.A2(n_606),
.B1(n_611),
.B2(n_601),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1422),
.A2(n_1224),
.B(n_1221),
.Y(n_1546)
);

AOI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1430),
.A2(n_1275),
.B(n_1083),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1480),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1422),
.A2(n_1224),
.B(n_1221),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_1492),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1461),
.Y(n_1551)
);

NOR2xp67_ASAP7_75t_L g1552 ( 
.A(n_1483),
.B(n_1224),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1493),
.B(n_1226),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1474),
.B(n_1082),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1474),
.B(n_1083),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1461),
.B(n_1087),
.Y(n_1556)
);

OAI22x1_ASAP7_75t_L g1557 ( 
.A1(n_1456),
.A2(n_607),
.B1(n_609),
.B2(n_597),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1444),
.A2(n_1235),
.B(n_1226),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1477),
.A2(n_1089),
.B(n_1094),
.C(n_1087),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1409),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1452),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1459),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1466),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_R g1564 ( 
.A(n_1443),
.B(n_641),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1473),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1409),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1476),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1413),
.A2(n_610),
.B1(n_613),
.B2(n_612),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1496),
.B(n_641),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1489),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1458),
.B(n_1446),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1436),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1485),
.B(n_1226),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1437),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1443),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1439),
.Y(n_1576)
);

NAND2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1448),
.B(n_1235),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1456),
.A2(n_1089),
.B(n_1095),
.C(n_1094),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1465),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1416),
.B(n_1095),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1458),
.B(n_1235),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1440),
.B(n_1096),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1429),
.A2(n_1154),
.B(n_1118),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1429),
.A2(n_1154),
.B(n_1118),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1465),
.Y(n_1585)
);

BUFx4f_ASAP7_75t_L g1586 ( 
.A(n_1448),
.Y(n_1586)
);

A2O1A1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1428),
.A2(n_1096),
.B(n_617),
.C(n_939),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1468),
.A2(n_1154),
.B(n_1158),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1447),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1468),
.A2(n_1154),
.B(n_1158),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1416),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1453),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1488),
.Y(n_1593)
);

NAND2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1413),
.B(n_614),
.Y(n_1594)
);

INVx3_ASAP7_75t_SL g1595 ( 
.A(n_1419),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1495),
.A2(n_749),
.B1(n_757),
.B2(n_641),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1450),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1419),
.B(n_619),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1561),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1500),
.B(n_620),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_SL g1601 ( 
.A1(n_1501),
.A2(n_1418),
.B(n_1495),
.C(n_618),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1506),
.B(n_1475),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1530),
.A2(n_1486),
.B(n_1482),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1594),
.A2(n_1418),
.B(n_1467),
.Y(n_1604)
);

INVx3_ASAP7_75t_SL g1605 ( 
.A(n_1512),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1521),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1510),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1547),
.A2(n_1454),
.B(n_1455),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1562),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1589),
.B(n_1402),
.Y(n_1610)
);

AO31x2_ASAP7_75t_L g1611 ( 
.A1(n_1592),
.A2(n_1471),
.A3(n_1487),
.B(n_1490),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1498),
.A2(n_1402),
.B(n_1450),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1499),
.A2(n_1491),
.B(n_1472),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1523),
.B(n_1529),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1535),
.B(n_749),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_SL g1616 ( 
.A(n_1528),
.B(n_890),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1546),
.A2(n_1423),
.B(n_1101),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1502),
.A2(n_617),
.B(n_717),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1579),
.B(n_609),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1532),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1520),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1588),
.A2(n_717),
.B(n_729),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1538),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1590),
.A2(n_807),
.B(n_796),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1549),
.A2(n_1108),
.B(n_1104),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1560),
.Y(n_1626)
);

O2A1O1Ixp5_ASAP7_75t_L g1627 ( 
.A1(n_1568),
.A2(n_623),
.B(n_625),
.C(n_618),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1514),
.Y(n_1628)
);

NOR4xp25_ASAP7_75t_L g1629 ( 
.A(n_1505),
.B(n_1554),
.C(n_1555),
.D(n_1571),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1503),
.A2(n_625),
.B(n_623),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1508),
.A2(n_813),
.B(n_741),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1558),
.A2(n_1108),
.B(n_1104),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_R g1633 ( 
.A(n_1550),
.B(n_749),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1533),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_R g1635 ( 
.A(n_1585),
.B(n_757),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1593),
.A2(n_1108),
.B(n_1104),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1533),
.Y(n_1637)
);

AOI221x1_ASAP7_75t_L g1638 ( 
.A1(n_1557),
.A2(n_629),
.B1(n_638),
.B2(n_635),
.C(n_627),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1597),
.A2(n_741),
.B(n_720),
.Y(n_1639)
);

A2O1A1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1569),
.A2(n_627),
.B(n_635),
.C(n_629),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1524),
.A2(n_1110),
.B(n_1109),
.Y(n_1641)
);

AO21x1_ASAP7_75t_L g1642 ( 
.A1(n_1517),
.A2(n_644),
.B(n_638),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1595),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1537),
.B(n_644),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1533),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1539),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1543),
.A2(n_1573),
.B(n_1581),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1560),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1563),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1583),
.A2(n_789),
.B(n_762),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1504),
.B(n_757),
.Y(n_1651)
);

AO31x2_ASAP7_75t_L g1652 ( 
.A1(n_1584),
.A2(n_1110),
.A3(n_1117),
.B(n_1109),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_R g1653 ( 
.A(n_1560),
.B(n_621),
.Y(n_1653)
);

AO31x2_ASAP7_75t_L g1654 ( 
.A1(n_1544),
.A2(n_1110),
.A3(n_1117),
.B(n_1109),
.Y(n_1654)
);

BUFx8_ASAP7_75t_L g1655 ( 
.A(n_1536),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1509),
.A2(n_649),
.B(n_648),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1518),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1507),
.Y(n_1658)
);

AOI21x1_ASAP7_75t_SL g1659 ( 
.A1(n_1598),
.A2(n_0),
.B(n_2),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1504),
.B(n_878),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1548),
.B(n_648),
.Y(n_1661)
);

INVxp67_ASAP7_75t_SL g1662 ( 
.A(n_1522),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1536),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1509),
.A2(n_789),
.B(n_762),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1525),
.B(n_649),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1526),
.B(n_1497),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1528),
.A2(n_893),
.B(n_854),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1536),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1565),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_SL g1670 ( 
.A(n_1564),
.B(n_626),
.C(n_622),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1566),
.B(n_1117),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1541),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1553),
.B(n_890),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1567),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1551),
.B(n_1119),
.Y(n_1675)
);

NOR2xp67_ASAP7_75t_L g1676 ( 
.A(n_1591),
.B(n_1541),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1527),
.A2(n_653),
.B(n_651),
.Y(n_1677)
);

AO221x2_ASAP7_75t_L g1678 ( 
.A1(n_1545),
.A2(n_655),
.B1(n_663),
.B2(n_653),
.C(n_651),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1576),
.B(n_655),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1513),
.A2(n_893),
.B(n_854),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1541),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1603),
.A2(n_1516),
.B(n_1542),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1630),
.A2(n_1578),
.B(n_1531),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1606),
.B(n_1531),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1620),
.B(n_1552),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1611),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1608),
.A2(n_1613),
.B(n_1617),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1604),
.A2(n_1577),
.B(n_1553),
.Y(n_1688)
);

BUFx8_ASAP7_75t_SL g1689 ( 
.A(n_1623),
.Y(n_1689)
);

NOR2x1_ASAP7_75t_R g1690 ( 
.A(n_1658),
.B(n_633),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1614),
.B(n_1570),
.Y(n_1691)
);

NAND2x1p5_ASAP7_75t_L g1692 ( 
.A(n_1647),
.B(n_1645),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1612),
.A2(n_1577),
.B(n_1559),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1629),
.A2(n_1596),
.B1(n_723),
.B2(n_724),
.C(n_716),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

AOI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1616),
.A2(n_1556),
.B(n_1582),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1611),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1618),
.A2(n_1625),
.B(n_1622),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1643),
.B(n_634),
.Y(n_1699)
);

BUFx4_ASAP7_75t_SL g1700 ( 
.A(n_1657),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1630),
.A2(n_1515),
.B(n_1587),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1636),
.A2(n_1580),
.B(n_1574),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1662),
.B(n_1572),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1602),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1602),
.B(n_663),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1616),
.A2(n_1534),
.B(n_1511),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1652),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1599),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1681),
.B(n_1575),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1624),
.A2(n_1511),
.B(n_1519),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1645),
.B(n_1586),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1632),
.A2(n_1120),
.B(n_1119),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1656),
.A2(n_1586),
.B(n_675),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1655),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1656),
.B(n_664),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1655),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1650),
.A2(n_1540),
.B(n_1120),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1621),
.B(n_664),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1669),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1674),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1610),
.B(n_1634),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1607),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1640),
.A2(n_1575),
.B1(n_677),
.B2(n_684),
.Y(n_1723)
);

CKINVDCx20_ASAP7_75t_R g1724 ( 
.A(n_1635),
.Y(n_1724)
);

INVx4_ASAP7_75t_SL g1725 ( 
.A(n_1611),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1609),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1681),
.B(n_1575),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1628),
.B(n_1119),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1672),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1641),
.A2(n_1120),
.B(n_1047),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1663),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1664),
.B(n_748),
.C(n_697),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1610),
.B(n_675),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1631),
.A2(n_684),
.B(n_677),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1642),
.B(n_615),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1652),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1643),
.A2(n_690),
.B1(n_692),
.B2(n_689),
.Y(n_1737)
);

A2O1A1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1667),
.A2(n_689),
.B(n_692),
.C(n_690),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1652),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1663),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1601),
.A2(n_1629),
.B(n_1673),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_1705),
.B(n_1619),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1721),
.B(n_1666),
.Y(n_1743)
);

OAI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1694),
.A2(n_1677),
.B(n_698),
.C(n_701),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1741),
.A2(n_1673),
.B(n_1678),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1687),
.A2(n_1659),
.B(n_1639),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1722),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1704),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1729),
.Y(n_1749)
);

AOI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1686),
.A2(n_1661),
.B(n_1644),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1706),
.A2(n_1678),
.B(n_1644),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1705),
.B(n_1661),
.Y(n_1752)
);

AOI22x1_ASAP7_75t_L g1753 ( 
.A1(n_1683),
.A2(n_1714),
.B1(n_1701),
.B2(n_1711),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1715),
.A2(n_1627),
.B(n_1677),
.C(n_1660),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1721),
.B(n_1665),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1695),
.Y(n_1756)
);

BUFx3_ASAP7_75t_L g1757 ( 
.A(n_1729),
.Y(n_1757)
);

NAND2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1688),
.B(n_1637),
.Y(n_1758)
);

AO21x2_ASAP7_75t_L g1759 ( 
.A1(n_1739),
.A2(n_1679),
.B(n_1619),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1685),
.B(n_1663),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1715),
.A2(n_1651),
.B(n_1600),
.C(n_1670),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1726),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1686),
.B(n_1654),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1685),
.B(n_1708),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1687),
.A2(n_1638),
.B(n_1679),
.Y(n_1765)
);

AOI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1697),
.A2(n_1676),
.B(n_1680),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1719),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1720),
.B(n_1654),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1710),
.A2(n_1637),
.B(n_1668),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1692),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1697),
.B(n_1654),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1692),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1707),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1692),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1682),
.A2(n_1626),
.B(n_1649),
.Y(n_1775)
);

AO21x2_ASAP7_75t_L g1776 ( 
.A1(n_1739),
.A2(n_1671),
.B(n_1675),
.Y(n_1776)
);

AOI21xp33_ASAP7_75t_L g1777 ( 
.A1(n_1735),
.A2(n_1733),
.B(n_1718),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1684),
.B(n_1668),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1738),
.A2(n_1713),
.B(n_1710),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1711),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1707),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1688),
.B(n_1668),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1691),
.Y(n_1783)
);

OA21x2_ASAP7_75t_L g1784 ( 
.A1(n_1682),
.A2(n_1736),
.B(n_1693),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1725),
.B(n_1626),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1690),
.B(n_1605),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1724),
.B(n_1653),
.Y(n_1787)
);

OA21x2_ASAP7_75t_L g1788 ( 
.A1(n_1736),
.A2(n_698),
.B(n_697),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1693),
.A2(n_1648),
.B(n_1671),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1685),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1767),
.Y(n_1791)
);

BUFx8_ASAP7_75t_L g1792 ( 
.A(n_1749),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1773),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1757),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1773),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1767),
.Y(n_1796)
);

AO21x2_ASAP7_75t_L g1797 ( 
.A1(n_1750),
.A2(n_1771),
.B(n_1763),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1781),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1768),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1743),
.B(n_1725),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1784),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1768),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1748),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1748),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1763),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1781),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1771),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1775),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1784),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1784),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1770),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1775),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1770),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1751),
.A2(n_1735),
.B1(n_1684),
.B2(n_1696),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1743),
.B(n_1725),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1745),
.A2(n_1732),
.B(n_1735),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1756),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_1757),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1783),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1774),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1784),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1774),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1788),
.Y(n_1823)
);

NAND2x1p5_ASAP7_75t_L g1824 ( 
.A(n_1788),
.B(n_1698),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1747),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1788),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1747),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1788),
.Y(n_1828)
);

AO21x2_ASAP7_75t_L g1829 ( 
.A1(n_1750),
.A2(n_1703),
.B(n_1717),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1762),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1764),
.B(n_1725),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1755),
.B(n_1733),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1762),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1772),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1758),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1764),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1772),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1782),
.Y(n_1838)
);

AO21x2_ASAP7_75t_L g1839 ( 
.A1(n_1779),
.A2(n_1717),
.B(n_1702),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1758),
.Y(n_1840)
);

OA21x2_ASAP7_75t_L g1841 ( 
.A1(n_1746),
.A2(n_1702),
.B(n_1698),
.Y(n_1841)
);

OA21x2_ASAP7_75t_L g1842 ( 
.A1(n_1746),
.A2(n_1730),
.B(n_1712),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1764),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1749),
.Y(n_1844)
);

OA21x2_ASAP7_75t_L g1845 ( 
.A1(n_1821),
.A2(n_1769),
.B(n_1789),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1814),
.A2(n_1753),
.B1(n_1742),
.B2(n_1735),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1818),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1799),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1814),
.A2(n_1753),
.B1(n_1742),
.B2(n_1759),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1818),
.A2(n_1754),
.B1(n_1752),
.B2(n_1777),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1797),
.A2(n_1816),
.B1(n_1809),
.B2(n_1810),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1801),
.A2(n_1766),
.B(n_1758),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1816),
.A2(n_1759),
.B1(n_1776),
.B2(n_1790),
.Y(n_1853)
);

OAI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1817),
.A2(n_706),
.B(n_701),
.Y(n_1854)
);

OAI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1832),
.A2(n_1790),
.B1(n_1780),
.B2(n_1778),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1797),
.A2(n_1759),
.B1(n_1776),
.B2(n_1765),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1794),
.B(n_1689),
.Y(n_1857)
);

A2O1A1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1805),
.A2(n_1761),
.B(n_1787),
.C(n_1744),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1821),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1821),
.Y(n_1860)
);

OAI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1832),
.A2(n_1780),
.B1(n_1711),
.B2(n_1783),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1821),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1832),
.A2(n_1737),
.B1(n_730),
.B2(n_736),
.C(n_709),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1824),
.Y(n_1864)
);

OA21x2_ASAP7_75t_L g1865 ( 
.A1(n_1808),
.A2(n_1766),
.B(n_1785),
.Y(n_1865)
);

OAI211xp5_ASAP7_75t_L g1866 ( 
.A1(n_1817),
.A2(n_1699),
.B(n_709),
.C(n_730),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1824),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1792),
.Y(n_1868)
);

AOI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1801),
.A2(n_706),
.B(n_744),
.C(n_736),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1792),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1799),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1797),
.A2(n_1776),
.B1(n_1765),
.B2(n_1717),
.Y(n_1872)
);

AOI33xp33_ASAP7_75t_L g1873 ( 
.A1(n_1805),
.A2(n_748),
.A3(n_755),
.B1(n_776),
.B2(n_758),
.B3(n_744),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1797),
.A2(n_1765),
.B1(n_1633),
.B2(n_1760),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1836),
.B(n_1749),
.Y(n_1875)
);

OAI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1805),
.A2(n_1780),
.B1(n_1728),
.B2(n_1749),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1859),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1859),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1864),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1848),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1848),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1871),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1859),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1864),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1871),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1860),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1860),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1860),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1852),
.B(n_1801),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1847),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1864),
.Y(n_1891)
);

NOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1847),
.B(n_1803),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1862),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1862),
.Y(n_1894)
);

OAI222xp33_ASAP7_75t_L g1895 ( 
.A1(n_1850),
.A2(n_1807),
.B1(n_1815),
.B2(n_1800),
.C1(n_1826),
.C2(n_1823),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1862),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1875),
.B(n_1836),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1875),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1851),
.B(n_1843),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1865),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1851),
.B(n_1843),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1865),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1850),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1845),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1845),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1847),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1845),
.Y(n_1907)
);

OAI31xp33_ASAP7_75t_L g1908 ( 
.A1(n_1895),
.A2(n_1858),
.A3(n_1874),
.B(n_1849),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1890),
.B(n_1868),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1900),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1903),
.B(n_1819),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1900),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1890),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1880),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1897),
.B(n_1843),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1880),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1897),
.B(n_1868),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1906),
.B(n_1689),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1903),
.B(n_1803),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1900),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1881),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1897),
.B(n_1868),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1881),
.B(n_1803),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1882),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1898),
.B(n_1870),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1882),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1898),
.B(n_1870),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1892),
.B(n_1870),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1906),
.B(n_1819),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1885),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1885),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1899),
.B(n_1804),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1899),
.B(n_1804),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1895),
.B(n_1857),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1894),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1899),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1894),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1902),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1892),
.B(n_1724),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1886),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1928),
.B(n_1901),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1928),
.B(n_1901),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1909),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1917),
.B(n_1901),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1936),
.A2(n_1908),
.B1(n_1934),
.B2(n_1863),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1928),
.B(n_1902),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1918),
.B(n_1786),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1919),
.B(n_1911),
.Y(n_1948)
);

OAI31xp33_ASAP7_75t_L g1949 ( 
.A1(n_1939),
.A2(n_1866),
.A3(n_1863),
.B(n_1854),
.Y(n_1949)
);

BUFx2_ASAP7_75t_L g1950 ( 
.A(n_1909),
.Y(n_1950)
);

OAI31xp33_ASAP7_75t_L g1951 ( 
.A1(n_1932),
.A2(n_1866),
.A3(n_1854),
.B(n_1904),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1936),
.A2(n_1853),
.B1(n_1846),
.B2(n_1856),
.Y(n_1952)
);

NOR2x1_ASAP7_75t_L g1953 ( 
.A(n_1913),
.B(n_1716),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1932),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1919),
.B(n_1886),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1910),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1917),
.B(n_1922),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1926),
.B(n_1888),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1922),
.B(n_1889),
.Y(n_1959)
);

NAND4xp25_ASAP7_75t_SL g1960 ( 
.A(n_1933),
.B(n_1873),
.C(n_1869),
.D(n_1904),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1909),
.B(n_1855),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1910),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1925),
.B(n_1889),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1914),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_L g1965 ( 
.A(n_1937),
.B(n_1716),
.Y(n_1965)
);

AO21x2_ASAP7_75t_L g1966 ( 
.A1(n_1912),
.A2(n_1907),
.B(n_1905),
.Y(n_1966)
);

AO21x2_ASAP7_75t_L g1967 ( 
.A1(n_1912),
.A2(n_1907),
.B(n_1905),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1925),
.B(n_1889),
.Y(n_1968)
);

AOI221xp5_ASAP7_75t_L g1969 ( 
.A1(n_1933),
.A2(n_1902),
.B1(n_755),
.B2(n_778),
.C(n_776),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1927),
.B(n_1889),
.Y(n_1970)
);

OAI31xp33_ASAP7_75t_L g1971 ( 
.A1(n_1937),
.A2(n_1872),
.A3(n_1861),
.B(n_1889),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1964),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1957),
.B(n_1927),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1966),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1951),
.B(n_1929),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1948),
.B(n_1935),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1966),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1964),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1954),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1954),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1954),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1951),
.B(n_1915),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1966),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1953),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1943),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1954),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1945),
.B(n_1915),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1956),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1945),
.B(n_1930),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1941),
.Y(n_1990)
);

OAI221xp5_ASAP7_75t_L g1991 ( 
.A1(n_1971),
.A2(n_1938),
.B1(n_1920),
.B2(n_1869),
.C(n_1940),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1969),
.B(n_1931),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1953),
.B(n_1714),
.Y(n_1993)
);

AOI21xp33_ASAP7_75t_L g1994 ( 
.A1(n_1965),
.A2(n_1938),
.B(n_1920),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1960),
.A2(n_1916),
.B(n_1914),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1957),
.B(n_1916),
.Y(n_1996)
);

NAND4xp25_ASAP7_75t_L g1997 ( 
.A(n_1943),
.B(n_1924),
.C(n_1921),
.D(n_1923),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1956),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1941),
.A2(n_1879),
.B1(n_1891),
.B2(n_1884),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1966),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1956),
.Y(n_2001)
);

AND2x4_ASAP7_75t_SL g2002 ( 
.A(n_1941),
.B(n_1942),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1944),
.B(n_1921),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1969),
.B(n_1924),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1962),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1950),
.B(n_1944),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1967),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1950),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1941),
.B(n_1923),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1949),
.B(n_1940),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1967),
.Y(n_2011)
);

INVx4_ASAP7_75t_L g2012 ( 
.A(n_1942),
.Y(n_2012)
);

AND2x2_ASAP7_75t_SL g2013 ( 
.A(n_1942),
.B(n_1700),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1948),
.B(n_1888),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1962),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_2006),
.B(n_1942),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_1949),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1987),
.B(n_1960),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1985),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1990),
.Y(n_2020)
);

NOR2xp67_ASAP7_75t_SL g2021 ( 
.A(n_1990),
.B(n_1961),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2008),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2013),
.B(n_1968),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1990),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2013),
.B(n_1968),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_2012),
.B(n_1947),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2003),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1997),
.B(n_1982),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1974),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1973),
.B(n_1970),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2004),
.B(n_1955),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_2003),
.B(n_1955),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1973),
.B(n_1970),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1972),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1996),
.B(n_1958),
.Y(n_2035)
);

OAI22xp33_ASAP7_75t_SL g2036 ( 
.A1(n_1991),
.A2(n_1975),
.B1(n_1984),
.B2(n_1989),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1984),
.B(n_1965),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_2002),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_2002),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2012),
.B(n_1959),
.Y(n_2040)
);

NOR2x1_ASAP7_75t_L g2041 ( 
.A(n_2012),
.B(n_1946),
.Y(n_2041)
);

NAND2x1p5_ASAP7_75t_L g2042 ( 
.A(n_1993),
.B(n_1946),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1996),
.B(n_1958),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2009),
.B(n_1959),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1972),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2009),
.B(n_1946),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1992),
.B(n_1962),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1995),
.B(n_1946),
.Y(n_2048)
);

INVxp67_ASAP7_75t_L g2049 ( 
.A(n_1988),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1978),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1979),
.B(n_1963),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1976),
.B(n_1986),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1978),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1976),
.B(n_2014),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1980),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1980),
.B(n_1952),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_2014),
.B(n_1967),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1981),
.B(n_1998),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1981),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2001),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1999),
.B(n_1967),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2001),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_1974),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1994),
.B(n_1879),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1977),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2005),
.B(n_1879),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1977),
.B(n_1971),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2015),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1983),
.B(n_1893),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1983),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2000),
.Y(n_2071)
);

NOR2xp67_ASAP7_75t_SL g2072 ( 
.A(n_2000),
.B(n_1615),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2007),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2007),
.B(n_1893),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2011),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2011),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1985),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1985),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_2002),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_2028),
.A2(n_1884),
.B1(n_1891),
.B2(n_1879),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2055),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2017),
.A2(n_1878),
.B1(n_1883),
.B2(n_1877),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2017),
.A2(n_1878),
.B1(n_1883),
.B2(n_1877),
.Y(n_2083)
);

AOI322xp5_ASAP7_75t_L g2084 ( 
.A1(n_2067),
.A2(n_1877),
.A3(n_1883),
.B1(n_1887),
.B2(n_1878),
.C1(n_1896),
.C2(n_1807),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_2016),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2055),
.Y(n_2086)
);

OAI21xp5_ASAP7_75t_SL g2087 ( 
.A1(n_2048),
.A2(n_2025),
.B(n_2023),
.Y(n_2087)
);

OR2x2_ASAP7_75t_L g2088 ( 
.A(n_2054),
.B(n_1884),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2067),
.A2(n_1887),
.B1(n_1896),
.B2(n_1891),
.Y(n_2089)
);

NAND3xp33_ASAP7_75t_L g2090 ( 
.A(n_2018),
.B(n_780),
.C(n_778),
.Y(n_2090)
);

OAI221xp5_ASAP7_75t_L g2091 ( 
.A1(n_2021),
.A2(n_1891),
.B1(n_1884),
.B2(n_1887),
.C(n_1810),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_2032),
.B(n_2027),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2063),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_2026),
.B(n_1864),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2046),
.B(n_1804),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2063),
.Y(n_2096)
);

AOI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_2036),
.A2(n_1845),
.B(n_1865),
.Y(n_2097)
);

AOI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_2037),
.A2(n_780),
.B(n_758),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2019),
.Y(n_2099)
);

OAI21xp33_ASAP7_75t_L g2100 ( 
.A1(n_2079),
.A2(n_1834),
.B(n_1844),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2030),
.B(n_783),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2033),
.B(n_783),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2022),
.Y(n_2103)
);

INVxp67_ASAP7_75t_SL g2104 ( 
.A(n_2026),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2077),
.Y(n_2105)
);

CKINVDCx14_ASAP7_75t_R g2106 ( 
.A(n_2039),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2078),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2020),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2020),
.Y(n_2109)
);

O2A1O1Ixp33_ASAP7_75t_L g2110 ( 
.A1(n_2047),
.A2(n_790),
.B(n_793),
.C(n_792),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2024),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_2039),
.B(n_1864),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2024),
.Y(n_2113)
);

INVxp67_ASAP7_75t_SL g2114 ( 
.A(n_2037),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2032),
.B(n_1791),
.Y(n_2115)
);

OAI33xp33_ASAP7_75t_L g2116 ( 
.A1(n_2031),
.A2(n_790),
.A3(n_792),
.B1(n_816),
.B2(n_793),
.B3(n_788),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_2038),
.Y(n_2117)
);

AOI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2056),
.A2(n_1797),
.B1(n_1867),
.B2(n_1864),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_2038),
.Y(n_2119)
);

AOI31xp33_ASAP7_75t_L g2120 ( 
.A1(n_2052),
.A2(n_816),
.A3(n_817),
.B(n_788),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_2047),
.A2(n_1867),
.B1(n_1809),
.B2(n_1810),
.Y(n_2121)
);

OAI221xp5_ASAP7_75t_L g2122 ( 
.A1(n_2031),
.A2(n_2057),
.B1(n_2042),
.B2(n_2049),
.C(n_2041),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2059),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2035),
.B(n_817),
.Y(n_2124)
);

INVx2_ASAP7_75t_SL g2125 ( 
.A(n_2040),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2044),
.B(n_1791),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2034),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2042),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_L g2129 ( 
.A(n_2043),
.B(n_1867),
.Y(n_2129)
);

OAI21xp5_ASAP7_75t_L g2130 ( 
.A1(n_2049),
.A2(n_1852),
.B(n_829),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_2051),
.Y(n_2131)
);

INVx1_ASAP7_75t_SL g2132 ( 
.A(n_2064),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2045),
.Y(n_2133)
);

A2O1A1Ixp33_ASAP7_75t_SL g2134 ( 
.A1(n_2050),
.A2(n_829),
.B(n_834),
.C(n_825),
.Y(n_2134)
);

NOR2xp67_ASAP7_75t_SL g2135 ( 
.A(n_2029),
.B(n_825),
.Y(n_2135)
);

OAI211xp5_ASAP7_75t_SL g2136 ( 
.A1(n_2058),
.A2(n_838),
.B(n_842),
.C(n_834),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2053),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2068),
.B(n_838),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_2058),
.Y(n_2139)
);

OAI21xp33_ASAP7_75t_L g2140 ( 
.A1(n_2066),
.A2(n_1834),
.B(n_1844),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_2072),
.A2(n_1867),
.B1(n_1810),
.B2(n_1809),
.Y(n_2141)
);

OAI21xp33_ASAP7_75t_L g2142 ( 
.A1(n_2061),
.A2(n_1834),
.B(n_1844),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2060),
.B(n_842),
.Y(n_2143)
);

AOI21xp33_ASAP7_75t_SL g2144 ( 
.A1(n_2062),
.A2(n_846),
.B(n_843),
.Y(n_2144)
);

NAND4xp25_ASAP7_75t_L g2145 ( 
.A(n_2070),
.B(n_846),
.C(n_847),
.D(n_843),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2029),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2071),
.Y(n_2147)
);

OAI31xp33_ASAP7_75t_L g2148 ( 
.A1(n_2073),
.A2(n_850),
.A3(n_857),
.B(n_847),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2069),
.A2(n_2074),
.B1(n_2065),
.B2(n_2075),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2076),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2065),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2069),
.B(n_2074),
.Y(n_2152)
);

OAI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_2018),
.A2(n_1867),
.B1(n_1801),
.B2(n_1810),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2046),
.B(n_850),
.Y(n_2154)
);

OAI21xp33_ASAP7_75t_L g2155 ( 
.A1(n_2028),
.A2(n_859),
.B(n_857),
.Y(n_2155)
);

AOI21xp33_ASAP7_75t_SL g2156 ( 
.A1(n_2026),
.A2(n_863),
.B(n_859),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2030),
.B(n_1791),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2046),
.B(n_863),
.Y(n_2158)
);

OAI322xp33_ASAP7_75t_L g2159 ( 
.A1(n_2028),
.A2(n_871),
.A3(n_868),
.B1(n_877),
.B2(n_882),
.C1(n_869),
.C2(n_866),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_2046),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2055),
.Y(n_2161)
);

OAI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2017),
.A2(n_1810),
.B1(n_1809),
.B2(n_1801),
.C(n_1867),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2055),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2046),
.B(n_866),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2055),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2030),
.B(n_1796),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2131),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2106),
.B(n_1796),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2117),
.Y(n_2169)
);

NOR2x1_ASAP7_75t_L g2170 ( 
.A(n_2081),
.B(n_868),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_2089),
.A2(n_1801),
.B1(n_1809),
.B2(n_1835),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2120),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2086),
.Y(n_2173)
);

OAI21xp33_ASAP7_75t_SL g2174 ( 
.A1(n_2114),
.A2(n_1796),
.B(n_1852),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2104),
.B(n_869),
.Y(n_2175)
);

OAI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2087),
.A2(n_926),
.B(n_913),
.Y(n_2176)
);

OAI22xp33_ASAP7_75t_L g2177 ( 
.A1(n_2097),
.A2(n_1809),
.B1(n_1840),
.B2(n_1835),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2159),
.A2(n_877),
.B(n_871),
.Y(n_2178)
);

A2O1A1Ixp33_ASAP7_75t_L g2179 ( 
.A1(n_2084),
.A2(n_886),
.B(n_892),
.C(n_882),
.Y(n_2179)
);

INVxp67_ASAP7_75t_L g2180 ( 
.A(n_2135),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_2085),
.B(n_1749),
.Y(n_2181)
);

OAI221xp5_ASAP7_75t_L g2182 ( 
.A1(n_2122),
.A2(n_894),
.B1(n_903),
.B2(n_892),
.C(n_886),
.Y(n_2182)
);

NAND3x2_ASAP7_75t_L g2183 ( 
.A(n_2092),
.B(n_903),
.C(n_894),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2161),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2139),
.B(n_908),
.Y(n_2185)
);

OAI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_2132),
.A2(n_1835),
.B1(n_1840),
.B2(n_1807),
.Y(n_2186)
);

OAI221xp5_ASAP7_75t_SL g2187 ( 
.A1(n_2091),
.A2(n_913),
.B1(n_917),
.B2(n_911),
.C(n_908),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2163),
.Y(n_2188)
);

INVxp67_ASAP7_75t_L g2189 ( 
.A(n_2160),
.Y(n_2189)
);

AO21x1_ASAP7_75t_L g2190 ( 
.A1(n_2165),
.A2(n_917),
.B(n_911),
.Y(n_2190)
);

INVxp33_ASAP7_75t_L g2191 ( 
.A(n_2101),
.Y(n_2191)
);

NAND3x2_ASAP7_75t_L g2192 ( 
.A(n_2099),
.B(n_926),
.C(n_924),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2125),
.Y(n_2193)
);

AOI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_2159),
.A2(n_930),
.B(n_924),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2108),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2119),
.B(n_930),
.Y(n_2196)
);

OAI322xp33_ASAP7_75t_L g2197 ( 
.A1(n_2093),
.A2(n_940),
.A3(n_936),
.B1(n_945),
.B2(n_952),
.C1(n_937),
.C2(n_931),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_R g2198 ( 
.A(n_2103),
.B(n_0),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_2136),
.B(n_931),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2109),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2156),
.B(n_936),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2111),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2113),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2102),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2134),
.B(n_937),
.Y(n_2205)
);

AOI321xp33_ASAP7_75t_L g2206 ( 
.A1(n_2149),
.A2(n_955),
.A3(n_945),
.B1(n_960),
.B2(n_952),
.C(n_940),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2154),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2146),
.A2(n_1839),
.B1(n_1865),
.B2(n_1829),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2158),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2128),
.B(n_955),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2126),
.B(n_960),
.Y(n_2211)
);

INVxp67_ASAP7_75t_L g2212 ( 
.A(n_2116),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2157),
.B(n_963),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_2164),
.Y(n_2214)
);

INVxp67_ASAP7_75t_SL g2215 ( 
.A(n_2124),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2166),
.B(n_2105),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2144),
.B(n_2155),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2096),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2143),
.Y(n_2219)
);

INVx1_ASAP7_75t_SL g2220 ( 
.A(n_2088),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2151),
.Y(n_2221)
);

O2A1O1Ixp33_ASAP7_75t_SL g2222 ( 
.A1(n_2107),
.A2(n_968),
.B(n_970),
.C(n_963),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2138),
.Y(n_2223)
);

OAI21xp33_ASAP7_75t_L g2224 ( 
.A1(n_2100),
.A2(n_970),
.B(n_968),
.Y(n_2224)
);

OAI322xp33_ASAP7_75t_L g2225 ( 
.A1(n_2147),
.A2(n_983),
.A3(n_979),
.B1(n_984),
.B2(n_985),
.C1(n_981),
.C2(n_971),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2090),
.Y(n_2226)
);

INVxp67_ASAP7_75t_L g2227 ( 
.A(n_2090),
.Y(n_2227)
);

AOI21xp33_ASAP7_75t_SL g2228 ( 
.A1(n_2080),
.A2(n_979),
.B(n_971),
.Y(n_2228)
);

AOI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2152),
.A2(n_1839),
.B1(n_1829),
.B2(n_1826),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2110),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2123),
.Y(n_2231)
);

AOI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_2082),
.A2(n_2083),
.B1(n_2118),
.B2(n_2112),
.Y(n_2232)
);

OAI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2130),
.A2(n_2094),
.B(n_2098),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_2145),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_2127),
.Y(n_2235)
);

OAI21xp33_ASAP7_75t_SL g2236 ( 
.A1(n_2133),
.A2(n_983),
.B(n_981),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2150),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2137),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2095),
.B(n_984),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2145),
.A2(n_987),
.B(n_985),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2129),
.B(n_2115),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2142),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2140),
.Y(n_2243)
);

OAI322xp33_ASAP7_75t_L g2244 ( 
.A1(n_2153),
.A2(n_2162),
.A3(n_2141),
.B1(n_996),
.B2(n_999),
.C1(n_990),
.C2(n_1012),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2121),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2148),
.A2(n_1840),
.B1(n_1835),
.B2(n_1837),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2148),
.B(n_987),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2120),
.B(n_990),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2117),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2120),
.B(n_991),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2131),
.Y(n_2251)
);

OAI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2114),
.A2(n_996),
.B(n_991),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2120),
.B(n_999),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_2085),
.B(n_878),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2106),
.B(n_1012),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2117),
.Y(n_2256)
);

OAI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2106),
.A2(n_1840),
.B1(n_1835),
.B2(n_1837),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2117),
.Y(n_2258)
);

AOI21xp33_ASAP7_75t_L g2259 ( 
.A1(n_2139),
.A2(n_974),
.B(n_928),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2160),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2117),
.Y(n_2261)
);

OAI21xp5_ASAP7_75t_L g2262 ( 
.A1(n_2114),
.A2(n_1022),
.B(n_1019),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2085),
.B(n_878),
.Y(n_2263)
);

AOI221xp5_ASAP7_75t_L g2264 ( 
.A1(n_2097),
.A2(n_1022),
.B1(n_1019),
.B2(n_797),
.C(n_798),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2117),
.Y(n_2265)
);

OAI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2114),
.A2(n_974),
.B(n_928),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2120),
.B(n_710),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2085),
.B(n_728),
.Y(n_2268)
);

OAI222xp33_ASAP7_75t_L g2269 ( 
.A1(n_2122),
.A2(n_1802),
.B1(n_1799),
.B2(n_1815),
.C1(n_1800),
.C2(n_1824),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_2120),
.B(n_799),
.Y(n_2270)
);

OAI221xp5_ASAP7_75t_L g2271 ( 
.A1(n_2097),
.A2(n_1011),
.B1(n_802),
.B2(n_806),
.C(n_801),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2120),
.B(n_800),
.Y(n_2272)
);

NAND3xp33_ASAP7_75t_L g2273 ( 
.A(n_2114),
.B(n_1011),
.C(n_811),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2160),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2120),
.B(n_809),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2117),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2117),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2106),
.B(n_1831),
.Y(n_2278)
);

A2O1A1Ixp33_ASAP7_75t_L g2279 ( 
.A1(n_2097),
.A2(n_639),
.B(n_643),
.C(n_642),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_2085),
.B(n_2),
.Y(n_2280)
);

OAI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2114),
.A2(n_652),
.B(n_646),
.Y(n_2281)
);

OAI221xp5_ASAP7_75t_L g2282 ( 
.A1(n_2097),
.A2(n_658),
.B1(n_660),
.B2(n_657),
.C(n_654),
.Y(n_2282)
);

AOI221xp5_ASAP7_75t_L g2283 ( 
.A1(n_2097),
.A2(n_666),
.B1(n_667),
.B2(n_662),
.C(n_661),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2117),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2117),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2106),
.B(n_1831),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2117),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2120),
.B(n_669),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2117),
.Y(n_2289)
);

INVx1_ASAP7_75t_SL g2290 ( 
.A(n_2131),
.Y(n_2290)
);

AO22x1_ASAP7_75t_L g2291 ( 
.A1(n_2114),
.A2(n_673),
.B1(n_674),
.B2(n_670),
.Y(n_2291)
);

NOR2x1_ASAP7_75t_L g2292 ( 
.A(n_2081),
.B(n_700),
.Y(n_2292)
);

NAND2xp33_ASAP7_75t_R g2293 ( 
.A(n_2092),
.B(n_3),
.Y(n_2293)
);

AOI222xp33_ASAP7_75t_L g2294 ( 
.A1(n_2149),
.A2(n_938),
.B1(n_925),
.B2(n_1826),
.C1(n_1828),
.C2(n_1823),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2120),
.B(n_676),
.Y(n_2295)
);

AOI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2114),
.A2(n_680),
.B(n_678),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2106),
.B(n_1831),
.Y(n_2297)
);

OAI21xp33_ASAP7_75t_L g2298 ( 
.A1(n_2087),
.A2(n_1813),
.B(n_1811),
.Y(n_2298)
);

NAND2x1_ASAP7_75t_L g2299 ( 
.A(n_2160),
.B(n_1835),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2114),
.A2(n_685),
.B(n_682),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2106),
.B(n_691),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2117),
.Y(n_2302)
);

O2A1O1Ixp5_ASAP7_75t_L g2303 ( 
.A1(n_2114),
.A2(n_1840),
.B(n_1811),
.C(n_1820),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2117),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2106),
.A2(n_1840),
.B1(n_1837),
.B2(n_1802),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2117),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2117),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2106),
.B(n_693),
.Y(n_2308)
);

INVx1_ASAP7_75t_SL g2309 ( 
.A(n_2085),
.Y(n_2309)
);

NAND2x1_ASAP7_75t_L g2310 ( 
.A(n_2160),
.B(n_700),
.Y(n_2310)
);

INVx2_ASAP7_75t_SL g2311 ( 
.A(n_2117),
.Y(n_2311)
);

AOI221xp5_ASAP7_75t_L g2312 ( 
.A1(n_2097),
.A2(n_702),
.B1(n_703),
.B2(n_699),
.C(n_695),
.Y(n_2312)
);

AOI21xp33_ASAP7_75t_L g2313 ( 
.A1(n_2139),
.A2(n_705),
.B(n_704),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2120),
.B(n_711),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2117),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2160),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2309),
.B(n_925),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2309),
.B(n_715),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_2311),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2167),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2290),
.B(n_925),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2197),
.B(n_938),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2251),
.Y(n_2323)
);

INVx1_ASAP7_75t_SL g2324 ( 
.A(n_2301),
.Y(n_2324)
);

AOI222xp33_ASAP7_75t_L g2325 ( 
.A1(n_2283),
.A2(n_938),
.B1(n_718),
.B2(n_714),
.C1(n_726),
.C2(n_725),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2291),
.B(n_727),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2255),
.Y(n_2327)
);

INVxp67_ASAP7_75t_L g2328 ( 
.A(n_2293),
.Y(n_2328)
);

AOI221xp5_ASAP7_75t_SL g2329 ( 
.A1(n_2302),
.A2(n_862),
.B1(n_898),
.B2(n_808),
.C(n_700),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2308),
.B(n_733),
.Y(n_2330)
);

AOI22xp33_ASAP7_75t_L g2331 ( 
.A1(n_2212),
.A2(n_1839),
.B1(n_1829),
.B2(n_1812),
.Y(n_2331)
);

OAI21xp33_ASAP7_75t_L g2332 ( 
.A1(n_2189),
.A2(n_1813),
.B(n_1811),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2172),
.B(n_734),
.Y(n_2333)
);

O2A1O1Ixp5_ASAP7_75t_L g2334 ( 
.A1(n_2181),
.A2(n_1813),
.B(n_1822),
.C(n_1820),
.Y(n_2334)
);

NAND2xp33_ASAP7_75t_R g2335 ( 
.A(n_2198),
.B(n_5),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2220),
.A2(n_1837),
.B1(n_1820),
.B2(n_1822),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2169),
.B(n_2249),
.Y(n_2337)
);

OAI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2256),
.A2(n_1822),
.B1(n_1802),
.B2(n_1876),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2216),
.B(n_721),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2190),
.Y(n_2340)
);

AOI221xp5_ASAP7_75t_L g2341 ( 
.A1(n_2282),
.A2(n_743),
.B1(n_747),
.B2(n_746),
.C(n_740),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2248),
.Y(n_2342)
);

AOI32xp33_ASAP7_75t_L g2343 ( 
.A1(n_2245),
.A2(n_2312),
.A3(n_2174),
.B1(n_2195),
.B2(n_2202),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_SL g2344 ( 
.A1(n_2258),
.A2(n_750),
.B1(n_775),
.B2(n_763),
.Y(n_2344)
);

NAND3xp33_ASAP7_75t_L g2345 ( 
.A(n_2206),
.B(n_754),
.C(n_752),
.Y(n_2345)
);

AOI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2232),
.A2(n_1839),
.B1(n_1760),
.B2(n_1815),
.Y(n_2346)
);

AOI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2264),
.A2(n_1839),
.B1(n_1760),
.B2(n_1800),
.Y(n_2347)
);

XOR2x2_ASAP7_75t_L g2348 ( 
.A(n_2183),
.B(n_1723),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2261),
.B(n_2265),
.Y(n_2349)
);

OAI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2276),
.A2(n_760),
.B(n_759),
.Y(n_2350)
);

AND3x1_ASAP7_75t_L g2351 ( 
.A(n_2260),
.B(n_1731),
.C(n_4),
.Y(n_2351)
);

AOI221xp5_ASAP7_75t_L g2352 ( 
.A1(n_2271),
.A2(n_767),
.B1(n_770),
.B2(n_769),
.C(n_765),
.Y(n_2352)
);

XNOR2xp5_ASAP7_75t_L g2353 ( 
.A(n_2192),
.B(n_772),
.Y(n_2353)
);

NAND3xp33_ASAP7_75t_L g2354 ( 
.A(n_2206),
.B(n_779),
.C(n_777),
.Y(n_2354)
);

AOI22x1_ASAP7_75t_L g2355 ( 
.A1(n_2193),
.A2(n_781),
.B1(n_787),
.B2(n_782),
.Y(n_2355)
);

OR2x2_ASAP7_75t_L g2356 ( 
.A(n_2277),
.B(n_4),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2284),
.B(n_795),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2250),
.Y(n_2358)
);

BUFx3_ASAP7_75t_L g2359 ( 
.A(n_2285),
.Y(n_2359)
);

OAI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2287),
.A2(n_1838),
.B1(n_812),
.B2(n_815),
.Y(n_2360)
);

OAI222xp33_ASAP7_75t_L g2361 ( 
.A1(n_2182),
.A2(n_1824),
.B1(n_1838),
.B2(n_821),
.C1(n_810),
.C2(n_823),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2253),
.Y(n_2362)
);

NOR3xp33_ASAP7_75t_L g2363 ( 
.A(n_2254),
.B(n_820),
.C(n_818),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2280),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2289),
.B(n_6),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2205),
.Y(n_2366)
);

INVx1_ASAP7_75t_SL g2367 ( 
.A(n_2288),
.Y(n_2367)
);

INVx1_ASAP7_75t_SL g2368 ( 
.A(n_2295),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2310),
.Y(n_2369)
);

NOR3xp33_ASAP7_75t_SL g2370 ( 
.A(n_2304),
.B(n_828),
.C(n_826),
.Y(n_2370)
);

AOI221xp5_ASAP7_75t_L g2371 ( 
.A1(n_2279),
.A2(n_831),
.B1(n_836),
.B2(n_833),
.C(n_832),
.Y(n_2371)
);

AOI221xp5_ASAP7_75t_L g2372 ( 
.A1(n_2179),
.A2(n_841),
.B1(n_853),
.B2(n_851),
.C(n_844),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2267),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2268),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_2197),
.B(n_855),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2306),
.B(n_858),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2278),
.B(n_860),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2307),
.B(n_6),
.Y(n_2378)
);

AOI211xp5_ASAP7_75t_L g2379 ( 
.A1(n_2187),
.A2(n_865),
.B(n_867),
.C(n_864),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2272),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_2235),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2315),
.B(n_870),
.Y(n_2382)
);

NAND3xp33_ASAP7_75t_L g2383 ( 
.A(n_2273),
.B(n_875),
.C(n_874),
.Y(n_2383)
);

NAND2x1p5_ASAP7_75t_L g2384 ( 
.A(n_2170),
.B(n_700),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2275),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_2225),
.B(n_876),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2222),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2211),
.B(n_880),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2270),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2213),
.B(n_881),
.Y(n_2390)
);

NAND2x1_ASAP7_75t_SL g2391 ( 
.A(n_2235),
.B(n_1731),
.Y(n_2391)
);

AOI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2221),
.A2(n_1765),
.B1(n_1838),
.B2(n_1829),
.Y(n_2392)
);

AOI211xp5_ASAP7_75t_L g2393 ( 
.A1(n_2269),
.A2(n_885),
.B(n_887),
.C(n_883),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2243),
.A2(n_1838),
.B1(n_891),
.B2(n_900),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2242),
.A2(n_901),
.B1(n_902),
.B2(n_888),
.Y(n_2395)
);

AOI31xp33_ASAP7_75t_SL g2396 ( 
.A1(n_2274),
.A2(n_9),
.A3(n_7),
.B(n_8),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2296),
.A2(n_2300),
.B(n_2225),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2199),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2247),
.Y(n_2399)
);

INVxp67_ASAP7_75t_L g2400 ( 
.A(n_2314),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_2316),
.B(n_808),
.Y(n_2401)
);

AOI211xp5_ASAP7_75t_L g2402 ( 
.A1(n_2228),
.A2(n_909),
.B(n_910),
.C(n_904),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2217),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2201),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2286),
.Y(n_2405)
);

INVx1_ASAP7_75t_SL g2406 ( 
.A(n_2297),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2185),
.Y(n_2407)
);

OAI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2233),
.A2(n_914),
.B(n_912),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_SL g2409 ( 
.A1(n_2241),
.A2(n_862),
.B(n_808),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2175),
.Y(n_2410)
);

OAI21xp33_ASAP7_75t_L g2411 ( 
.A1(n_2298),
.A2(n_922),
.B(n_921),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2230),
.Y(n_2412)
);

OAI22xp33_ASAP7_75t_L g2413 ( 
.A1(n_2191),
.A2(n_1823),
.B1(n_1828),
.B2(n_1826),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2168),
.B(n_923),
.Y(n_2414)
);

OR2x2_ASAP7_75t_L g2415 ( 
.A(n_2196),
.B(n_7),
.Y(n_2415)
);

OAI31xp33_ASAP7_75t_L g2416 ( 
.A1(n_2177),
.A2(n_1824),
.A3(n_1828),
.B(n_1823),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2281),
.B(n_2200),
.Y(n_2417)
);

AOI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2215),
.A2(n_1829),
.B1(n_929),
.B2(n_933),
.Y(n_2418)
);

AOI322xp5_ASAP7_75t_L g2419 ( 
.A1(n_2226),
.A2(n_1828),
.A3(n_1812),
.B1(n_1808),
.B2(n_942),
.C1(n_934),
.C2(n_935),
.Y(n_2419)
);

AOI32xp33_ASAP7_75t_L g2420 ( 
.A1(n_2203),
.A2(n_944),
.A3(n_948),
.B1(n_941),
.B2(n_927),
.Y(n_2420)
);

OAI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2234),
.A2(n_953),
.B(n_949),
.Y(n_2421)
);

AOI31xp33_ASAP7_75t_L g2422 ( 
.A1(n_2173),
.A2(n_956),
.A3(n_957),
.B(n_954),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2210),
.B(n_959),
.Y(n_2423)
);

OA21x2_ASAP7_75t_SL g2424 ( 
.A1(n_2263),
.A2(n_1727),
.B(n_1709),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_SL g2425 ( 
.A1(n_2184),
.A2(n_982),
.B1(n_1014),
.B2(n_965),
.Y(n_2425)
);

AOI21xp33_ASAP7_75t_SL g2426 ( 
.A1(n_2188),
.A2(n_988),
.B(n_966),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2219),
.B(n_961),
.Y(n_2427)
);

OAI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2180),
.A2(n_1780),
.B1(n_1812),
.B2(n_1808),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2273),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2204),
.B(n_964),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2223),
.B(n_969),
.Y(n_2431)
);

OAI221xp5_ASAP7_75t_L g2432 ( 
.A1(n_2236),
.A2(n_976),
.B1(n_977),
.B2(n_975),
.C(n_972),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2218),
.B(n_1709),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2239),
.Y(n_2434)
);

AOI221xp5_ASAP7_75t_L g2435 ( 
.A1(n_2244),
.A2(n_989),
.B1(n_992),
.B2(n_986),
.C(n_978),
.Y(n_2435)
);

AOI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_2422),
.A2(n_2262),
.B(n_2252),
.Y(n_2436)
);

OAI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2397),
.A2(n_2237),
.B(n_2231),
.Y(n_2437)
);

NAND4xp25_ASAP7_75t_SL g2438 ( 
.A(n_2406),
.B(n_2238),
.C(n_2294),
.D(n_2207),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2324),
.B(n_2239),
.Y(n_2439)
);

OAI211xp5_ASAP7_75t_SL g2440 ( 
.A1(n_2343),
.A2(n_2224),
.B(n_2303),
.C(n_2176),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2381),
.Y(n_2441)
);

OAI221xp5_ASAP7_75t_L g2442 ( 
.A1(n_2328),
.A2(n_2266),
.B1(n_2227),
.B2(n_2214),
.C(n_2209),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2327),
.B(n_2319),
.Y(n_2443)
);

OAI22xp33_ASAP7_75t_L g2444 ( 
.A1(n_2318),
.A2(n_2299),
.B1(n_2246),
.B2(n_2305),
.Y(n_2444)
);

NOR3xp33_ASAP7_75t_L g2445 ( 
.A(n_2317),
.B(n_2259),
.C(n_2292),
.Y(n_2445)
);

OAI211xp5_ASAP7_75t_L g2446 ( 
.A1(n_2319),
.A2(n_2313),
.B(n_2257),
.C(n_2186),
.Y(n_2446)
);

AOI221xp5_ASAP7_75t_L g2447 ( 
.A1(n_2400),
.A2(n_2244),
.B1(n_2208),
.B2(n_2229),
.C(n_2171),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2326),
.A2(n_2194),
.B(n_2178),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2381),
.B(n_2240),
.Y(n_2449)
);

NAND3xp33_ASAP7_75t_SL g2450 ( 
.A(n_2363),
.B(n_997),
.C(n_995),
.Y(n_2450)
);

AOI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2339),
.A2(n_1004),
.B(n_1000),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2405),
.B(n_1007),
.Y(n_2452)
);

HB1xp67_ASAP7_75t_L g2453 ( 
.A(n_2335),
.Y(n_2453)
);

OAI221xp5_ASAP7_75t_L g2454 ( 
.A1(n_2393),
.A2(n_1010),
.B1(n_1015),
.B2(n_1009),
.C(n_1008),
.Y(n_2454)
);

AOI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2425),
.A2(n_1017),
.B(n_1016),
.Y(n_2455)
);

NOR4xp25_ASAP7_75t_L g2456 ( 
.A(n_2320),
.B(n_11),
.C(n_8),
.D(n_10),
.Y(n_2456)
);

AOI21xp33_ASAP7_75t_L g2457 ( 
.A1(n_2340),
.A2(n_1021),
.B(n_862),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_L g2458 ( 
.A(n_2387),
.B(n_10),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2323),
.B(n_862),
.Y(n_2459)
);

OAI221xp5_ASAP7_75t_L g2460 ( 
.A1(n_2321),
.A2(n_898),
.B1(n_943),
.B2(n_862),
.C(n_808),
.Y(n_2460)
);

OAI221xp5_ASAP7_75t_L g2461 ( 
.A1(n_2367),
.A2(n_943),
.B1(n_1013),
.B2(n_898),
.C(n_808),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2359),
.B(n_898),
.Y(n_2462)
);

NAND3xp33_ASAP7_75t_L g2463 ( 
.A(n_2419),
.B(n_943),
.C(n_898),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2368),
.A2(n_1013),
.B1(n_943),
.B2(n_615),
.C(n_753),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2353),
.Y(n_2465)
);

NOR3xp33_ASAP7_75t_L g2466 ( 
.A(n_2361),
.B(n_753),
.C(n_712),
.Y(n_2466)
);

OAI311xp33_ASAP7_75t_L g2467 ( 
.A1(n_2331),
.A2(n_1731),
.A3(n_15),
.B1(n_12),
.C1(n_13),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2344),
.A2(n_1013),
.B(n_943),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_SL g2469 ( 
.A(n_2337),
.B(n_1013),
.Y(n_2469)
);

AOI221xp5_ASAP7_75t_L g2470 ( 
.A1(n_2412),
.A2(n_2395),
.B1(n_2394),
.B2(n_2351),
.C(n_2333),
.Y(n_2470)
);

OAI211xp5_ASAP7_75t_L g2471 ( 
.A1(n_2349),
.A2(n_1013),
.B(n_15),
.C(n_12),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2356),
.Y(n_2472)
);

AOI222xp33_ASAP7_75t_L g2473 ( 
.A1(n_2429),
.A2(n_890),
.B1(n_1808),
.B2(n_1812),
.C1(n_803),
.C2(n_1825),
.Y(n_2473)
);

NAND2x1p5_ASAP7_75t_L g2474 ( 
.A(n_2355),
.B(n_13),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2408),
.A2(n_1727),
.B(n_1709),
.Y(n_2475)
);

AOI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2364),
.A2(n_1727),
.B1(n_1785),
.B2(n_1833),
.Y(n_2476)
);

AOI221xp5_ASAP7_75t_L g2477 ( 
.A1(n_2426),
.A2(n_1827),
.B1(n_1830),
.B2(n_1825),
.C(n_1833),
.Y(n_2477)
);

AOI21xp5_ASAP7_75t_L g2478 ( 
.A1(n_2430),
.A2(n_1841),
.B(n_1728),
.Y(n_2478)
);

OAI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2377),
.A2(n_1740),
.B(n_1734),
.Y(n_2479)
);

AOI222xp33_ASAP7_75t_L g2480 ( 
.A1(n_2322),
.A2(n_1830),
.B1(n_1825),
.B2(n_1827),
.C1(n_1833),
.C2(n_588),
.Y(n_2480)
);

AOI21xp5_ASAP7_75t_L g2481 ( 
.A1(n_2330),
.A2(n_1841),
.B(n_1728),
.Y(n_2481)
);

AOI322xp5_ASAP7_75t_L g2482 ( 
.A1(n_2403),
.A2(n_1830),
.A3(n_1827),
.B1(n_1833),
.B2(n_1798),
.C1(n_1795),
.C2(n_1806),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2384),
.Y(n_2483)
);

AOI222xp33_ASAP7_75t_L g2484 ( 
.A1(n_2366),
.A2(n_2380),
.B1(n_2385),
.B2(n_2373),
.C1(n_2417),
.C2(n_2404),
.Y(n_2484)
);

NAND4xp25_ASAP7_75t_SL g2485 ( 
.A(n_2420),
.B(n_1792),
.C(n_18),
.D(n_16),
.Y(n_2485)
);

AOI22xp33_ASAP7_75t_SL g2486 ( 
.A1(n_2342),
.A2(n_1780),
.B1(n_1785),
.B2(n_1792),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2370),
.B(n_17),
.Y(n_2487)
);

AOI221xp5_ASAP7_75t_L g2488 ( 
.A1(n_2426),
.A2(n_588),
.B1(n_636),
.B2(n_656),
.C(n_608),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2365),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_L g2490 ( 
.A(n_2409),
.B(n_686),
.C(n_681),
.Y(n_2490)
);

AOI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2427),
.A2(n_1841),
.B(n_1728),
.Y(n_2491)
);

AOI311xp33_ASAP7_75t_L g2492 ( 
.A1(n_2357),
.A2(n_21),
.A3(n_18),
.B(n_20),
.C(n_23),
.Y(n_2492)
);

AOI21xp33_ASAP7_75t_SL g2493 ( 
.A1(n_2378),
.A2(n_2360),
.B(n_2376),
.Y(n_2493)
);

AOI211xp5_ASAP7_75t_L g2494 ( 
.A1(n_2396),
.A2(n_25),
.B(n_21),
.C(n_24),
.Y(n_2494)
);

OAI221xp5_ASAP7_75t_L g2495 ( 
.A1(n_2418),
.A2(n_1782),
.B1(n_1841),
.B2(n_1795),
.C(n_1798),
.Y(n_2495)
);

OAI221xp5_ASAP7_75t_L g2496 ( 
.A1(n_2391),
.A2(n_1782),
.B1(n_1841),
.B2(n_1795),
.C(n_1798),
.Y(n_2496)
);

NAND4xp25_ASAP7_75t_L g2497 ( 
.A(n_2424),
.B(n_2411),
.C(n_2325),
.D(n_2329),
.Y(n_2497)
);

OAI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_2433),
.A2(n_2382),
.B1(n_2414),
.B2(n_2431),
.Y(n_2498)
);

AOI221xp5_ASAP7_75t_L g2499 ( 
.A1(n_2358),
.A2(n_588),
.B1(n_738),
.B2(n_751),
.C(n_694),
.Y(n_2499)
);

AOI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2388),
.A2(n_1785),
.B1(n_1841),
.B2(n_1795),
.Y(n_2500)
);

OAI211xp5_ASAP7_75t_SL g2501 ( 
.A1(n_2371),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2501)
);

NAND5xp2_ASAP7_75t_L g2502 ( 
.A(n_2346),
.B(n_29),
.C(n_27),
.D(n_28),
.E(n_30),
.Y(n_2502)
);

OAI31xp33_ASAP7_75t_L g2503 ( 
.A1(n_2362),
.A2(n_1793),
.A3(n_1806),
.B(n_1798),
.Y(n_2503)
);

NAND3xp33_ASAP7_75t_L g2504 ( 
.A(n_2402),
.B(n_588),
.C(n_756),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_SL g2505 ( 
.A(n_2379),
.B(n_774),
.C(n_764),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2375),
.B(n_29),
.Y(n_2506)
);

AOI321xp33_ASAP7_75t_L g2507 ( 
.A1(n_2347),
.A2(n_2369),
.A3(n_2407),
.B1(n_2410),
.B2(n_2389),
.C(n_2434),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2390),
.A2(n_30),
.B(n_31),
.Y(n_2508)
);

A2O1A1Ixp33_ASAP7_75t_L g2509 ( 
.A1(n_2386),
.A2(n_1734),
.B(n_1806),
.C(n_1793),
.Y(n_2509)
);

AOI221xp5_ASAP7_75t_L g2510 ( 
.A1(n_2372),
.A2(n_588),
.B1(n_805),
.B2(n_837),
.C(n_804),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2415),
.Y(n_2511)
);

AOI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2423),
.A2(n_1793),
.B1(n_1806),
.B2(n_1648),
.Y(n_2512)
);

AOI32xp33_ASAP7_75t_L g2513 ( 
.A1(n_2433),
.A2(n_37),
.A3(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_2513)
);

AO22x1_ASAP7_75t_L g2514 ( 
.A1(n_2350),
.A2(n_1792),
.B1(n_40),
.B2(n_32),
.Y(n_2514)
);

NOR3xp33_ASAP7_75t_L g2515 ( 
.A(n_2383),
.B(n_856),
.C(n_845),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2401),
.A2(n_37),
.B(n_41),
.Y(n_2516)
);

AOI221xp5_ASAP7_75t_L g2517 ( 
.A1(n_2352),
.A2(n_962),
.B1(n_1002),
.B2(n_946),
.C(n_861),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2398),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2374),
.A2(n_1793),
.B1(n_1648),
.B2(n_1792),
.Y(n_2519)
);

BUFx12f_ASAP7_75t_L g2520 ( 
.A(n_2421),
.Y(n_2520)
);

AOI221xp5_ASAP7_75t_L g2521 ( 
.A1(n_2432),
.A2(n_1003),
.B1(n_43),
.B2(n_41),
.C(n_42),
.Y(n_2521)
);

NOR2x1_ASAP7_75t_L g2522 ( 
.A(n_2345),
.B(n_42),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2435),
.A2(n_43),
.B(n_44),
.Y(n_2523)
);

AOI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2341),
.A2(n_44),
.B(n_45),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2354),
.A2(n_46),
.B(n_47),
.Y(n_2525)
);

AOI21xp33_ASAP7_75t_SL g2526 ( 
.A1(n_2399),
.A2(n_46),
.B(n_47),
.Y(n_2526)
);

AOI221xp5_ASAP7_75t_L g2527 ( 
.A1(n_2413),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_2527)
);

AOI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2348),
.A2(n_1842),
.B1(n_1115),
.B2(n_51),
.Y(n_2528)
);

O2A1O1Ixp33_ASAP7_75t_L g2529 ( 
.A1(n_2336),
.A2(n_53),
.B(n_48),
.C(n_50),
.Y(n_2529)
);

AOI311xp33_ASAP7_75t_L g2530 ( 
.A1(n_2428),
.A2(n_56),
.A3(n_53),
.B(n_54),
.C(n_58),
.Y(n_2530)
);

OAI221xp5_ASAP7_75t_SL g2531 ( 
.A1(n_2416),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_2531)
);

NAND2x1p5_ASAP7_75t_L g2532 ( 
.A(n_2424),
.B(n_62),
.Y(n_2532)
);

AOI311xp33_ASAP7_75t_L g2533 ( 
.A1(n_2338),
.A2(n_65),
.A3(n_63),
.B(n_64),
.C(n_66),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2334),
.Y(n_2534)
);

AOI221xp5_ASAP7_75t_L g2535 ( 
.A1(n_2392),
.A2(n_66),
.B1(n_63),
.B2(n_64),
.C(n_67),
.Y(n_2535)
);

AOI22xp5_ASAP7_75t_SL g2536 ( 
.A1(n_2332),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2536)
);

OAI21xp33_ASAP7_75t_L g2537 ( 
.A1(n_2406),
.A2(n_69),
.B(n_70),
.Y(n_2537)
);

AOI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2422),
.A2(n_70),
.B(n_72),
.Y(n_2538)
);

NOR3xp33_ASAP7_75t_L g2539 ( 
.A(n_2328),
.B(n_73),
.C(n_74),
.Y(n_2539)
);

OAI21xp33_ASAP7_75t_L g2540 ( 
.A1(n_2406),
.A2(n_74),
.B(n_75),
.Y(n_2540)
);

OAI21xp33_ASAP7_75t_L g2541 ( 
.A1(n_2406),
.A2(n_75),
.B(n_76),
.Y(n_2541)
);

NOR3xp33_ASAP7_75t_L g2542 ( 
.A(n_2328),
.B(n_76),
.C(n_77),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_L g2543 ( 
.A(n_2324),
.B(n_78),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_2319),
.B(n_78),
.Y(n_2544)
);

OAI211xp5_ASAP7_75t_SL g2545 ( 
.A1(n_2343),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2319),
.B(n_79),
.Y(n_2546)
);

AOI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2422),
.A2(n_80),
.B(n_83),
.Y(n_2547)
);

OAI21xp33_ASAP7_75t_L g2548 ( 
.A1(n_2406),
.A2(n_83),
.B(n_84),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2324),
.B(n_85),
.Y(n_2549)
);

A2O1A1Ixp33_ASAP7_75t_L g2550 ( 
.A1(n_2343),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_L g2551 ( 
.A(n_2328),
.B(n_89),
.C(n_90),
.Y(n_2551)
);

NOR2x1_ASAP7_75t_L g2552 ( 
.A(n_2319),
.B(n_91),
.Y(n_2552)
);

NAND3xp33_ASAP7_75t_SL g2553 ( 
.A(n_2324),
.B(n_92),
.C(n_93),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2324),
.B(n_92),
.Y(n_2554)
);

AOI322xp5_ASAP7_75t_L g2555 ( 
.A1(n_2328),
.A2(n_104),
.A3(n_99),
.B1(n_96),
.B2(n_94),
.C1(n_95),
.C2(n_97),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2324),
.B(n_99),
.Y(n_2556)
);

A2O1A1Ixp33_ASAP7_75t_L g2557 ( 
.A1(n_2343),
.A2(n_108),
.B(n_105),
.C(n_107),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2366),
.A2(n_1842),
.B1(n_1115),
.B2(n_1712),
.Y(n_2558)
);

OAI221xp5_ASAP7_75t_L g2559 ( 
.A1(n_2343),
.A2(n_1842),
.B1(n_109),
.B2(n_105),
.C(n_107),
.Y(n_2559)
);

INVxp67_ASAP7_75t_L g2560 ( 
.A(n_2335),
.Y(n_2560)
);

AOI221xp5_ASAP7_75t_L g2561 ( 
.A1(n_2343),
.A2(n_113),
.B1(n_110),
.B2(n_111),
.C(n_114),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2324),
.B(n_110),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2324),
.B(n_113),
.Y(n_2563)
);

AOI211xp5_ASAP7_75t_L g2564 ( 
.A1(n_2406),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2564)
);

OAI221xp5_ASAP7_75t_L g2565 ( 
.A1(n_2343),
.A2(n_1842),
.B1(n_118),
.B2(n_115),
.C(n_116),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2351),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2319),
.B(n_118),
.Y(n_2567)
);

HB1xp67_ASAP7_75t_L g2568 ( 
.A(n_2381),
.Y(n_2568)
);

NOR3xp33_ASAP7_75t_L g2569 ( 
.A(n_2328),
.B(n_119),
.C(n_121),
.Y(n_2569)
);

O2A1O1Ixp5_ASAP7_75t_L g2570 ( 
.A1(n_2381),
.A2(n_123),
.B(n_119),
.C(n_122),
.Y(n_2570)
);

OAI21xp33_ASAP7_75t_L g2571 ( 
.A1(n_2406),
.A2(n_122),
.B(n_124),
.Y(n_2571)
);

AOI211xp5_ASAP7_75t_L g2572 ( 
.A1(n_2406),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_2572)
);

AOI221xp5_ASAP7_75t_L g2573 ( 
.A1(n_2343),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.C(n_130),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2319),
.B(n_128),
.Y(n_2574)
);

NOR3xp33_ASAP7_75t_L g2575 ( 
.A(n_2328),
.B(n_131),
.C(n_132),
.Y(n_2575)
);

AOI22xp33_ASAP7_75t_L g2576 ( 
.A1(n_2366),
.A2(n_1842),
.B1(n_1115),
.B2(n_1141),
.Y(n_2576)
);

OAI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2397),
.A2(n_131),
.B(n_133),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2381),
.Y(n_2578)
);

O2A1O1Ixp5_ASAP7_75t_L g2579 ( 
.A1(n_2381),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_2579)
);

AOI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2324),
.A2(n_1842),
.B1(n_1115),
.B2(n_138),
.Y(n_2580)
);

AOI221xp5_ASAP7_75t_L g2581 ( 
.A1(n_2343),
.A2(n_138),
.B1(n_134),
.B2(n_135),
.C(n_139),
.Y(n_2581)
);

A2O1A1Ixp33_ASAP7_75t_L g2582 ( 
.A1(n_2343),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_2582)
);

NAND3xp33_ASAP7_75t_SL g2583 ( 
.A(n_2324),
.B(n_143),
.C(n_144),
.Y(n_2583)
);

AOI221xp5_ASAP7_75t_L g2584 ( 
.A1(n_2343),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2453),
.Y(n_2585)
);

AOI21x1_ASAP7_75t_L g2586 ( 
.A1(n_2568),
.A2(n_146),
.B(n_147),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2546),
.Y(n_2587)
);

AOI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2544),
.A2(n_149),
.B(n_150),
.Y(n_2588)
);

NAND5xp2_ASAP7_75t_L g2589 ( 
.A(n_2507),
.B(n_152),
.C(n_150),
.D(n_151),
.E(n_153),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_SL g2590 ( 
.A(n_2543),
.B(n_151),
.Y(n_2590)
);

AOI211xp5_ASAP7_75t_L g2591 ( 
.A1(n_2559),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_2591)
);

AOI21xp33_ASAP7_75t_L g2592 ( 
.A1(n_2560),
.A2(n_155),
.B(n_156),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2567),
.Y(n_2593)
);

O2A1O1Ixp33_ASAP7_75t_L g2594 ( 
.A1(n_2550),
.A2(n_2582),
.B(n_2557),
.C(n_2545),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_SL g2595 ( 
.A1(n_2520),
.A2(n_160),
.B1(n_157),
.B2(n_158),
.Y(n_2595)
);

INVxp67_ASAP7_75t_L g2596 ( 
.A(n_2552),
.Y(n_2596)
);

A2O1A1Ixp33_ASAP7_75t_L g2597 ( 
.A1(n_2534),
.A2(n_161),
.B(n_158),
.C(n_160),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2574),
.B(n_161),
.Y(n_2598)
);

AOI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2443),
.A2(n_162),
.B(n_163),
.Y(n_2599)
);

OAI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2549),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_2600)
);

INVx2_ASAP7_75t_SL g2601 ( 
.A(n_2441),
.Y(n_2601)
);

INVx1_ASAP7_75t_SL g2602 ( 
.A(n_2474),
.Y(n_2602)
);

NOR2x1_ASAP7_75t_L g2603 ( 
.A(n_2578),
.B(n_164),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2553),
.B(n_166),
.Y(n_2604)
);

AOI211xp5_ASAP7_75t_SL g2605 ( 
.A1(n_2449),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_2605)
);

INVx1_ASAP7_75t_SL g2606 ( 
.A(n_2474),
.Y(n_2606)
);

INVx1_ASAP7_75t_SL g2607 ( 
.A(n_2487),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_SL g2608 ( 
.A(n_2563),
.B(n_167),
.Y(n_2608)
);

A2O1A1Ixp33_ASAP7_75t_L g2609 ( 
.A1(n_2584),
.A2(n_171),
.B(n_168),
.C(n_170),
.Y(n_2609)
);

OAI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2554),
.A2(n_174),
.B1(n_171),
.B2(n_173),
.Y(n_2610)
);

NAND2x1_ASAP7_75t_SL g2611 ( 
.A(n_2452),
.B(n_173),
.Y(n_2611)
);

CKINVDCx6p67_ASAP7_75t_R g2612 ( 
.A(n_2556),
.Y(n_2612)
);

OAI21xp5_ASAP7_75t_SL g2613 ( 
.A1(n_2440),
.A2(n_174),
.B(n_175),
.Y(n_2613)
);

OAI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2570),
.A2(n_175),
.B(n_176),
.Y(n_2614)
);

OAI322xp33_ASAP7_75t_L g2615 ( 
.A1(n_2565),
.A2(n_176),
.A3(n_177),
.B1(n_178),
.B2(n_179),
.C1(n_181),
.C2(n_182),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2439),
.Y(n_2616)
);

NOR2x1_ASAP7_75t_L g2617 ( 
.A(n_2450),
.B(n_177),
.Y(n_2617)
);

AOI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2561),
.A2(n_183),
.B1(n_178),
.B2(n_179),
.C(n_184),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2566),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_2619)
);

AOI32xp33_ASAP7_75t_L g2620 ( 
.A1(n_2573),
.A2(n_189),
.A3(n_185),
.B1(n_187),
.B2(n_191),
.Y(n_2620)
);

OAI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2579),
.A2(n_189),
.B(n_192),
.Y(n_2621)
);

OAI221xp5_ASAP7_75t_L g2622 ( 
.A1(n_2581),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.C(n_196),
.Y(n_2622)
);

AOI22xp5_ASAP7_75t_L g2623 ( 
.A1(n_2528),
.A2(n_197),
.B1(n_193),
.B2(n_196),
.Y(n_2623)
);

NAND4xp25_ASAP7_75t_L g2624 ( 
.A(n_2437),
.B(n_200),
.C(n_197),
.D(n_198),
.Y(n_2624)
);

AOI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2493),
.A2(n_203),
.B1(n_198),
.B2(n_202),
.C(n_204),
.Y(n_2625)
);

AOI221xp5_ASAP7_75t_L g2626 ( 
.A1(n_2498),
.A2(n_206),
.B1(n_203),
.B2(n_205),
.C(n_207),
.Y(n_2626)
);

AOI21xp5_ASAP7_75t_L g2627 ( 
.A1(n_2436),
.A2(n_205),
.B(n_206),
.Y(n_2627)
);

XNOR2x1_ASAP7_75t_L g2628 ( 
.A(n_2532),
.B(n_2522),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2494),
.B(n_207),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2456),
.B(n_208),
.Y(n_2630)
);

AOI22x1_ASAP7_75t_L g2631 ( 
.A1(n_2536),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_2631)
);

INVxp67_ASAP7_75t_SL g2632 ( 
.A(n_2562),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2472),
.Y(n_2633)
);

A2O1A1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2529),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_2634)
);

OAI221xp5_ASAP7_75t_L g2635 ( 
.A1(n_2577),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.C(n_216),
.Y(n_2635)
);

AOI221xp5_ASAP7_75t_SL g2636 ( 
.A1(n_2444),
.A2(n_217),
.B1(n_214),
.B2(n_215),
.C(n_218),
.Y(n_2636)
);

OAI21xp33_ASAP7_75t_L g2637 ( 
.A1(n_2519),
.A2(n_217),
.B(n_218),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2583),
.B(n_220),
.Y(n_2638)
);

OAI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2551),
.A2(n_224),
.B1(n_220),
.B2(n_221),
.Y(n_2639)
);

BUFx2_ASAP7_75t_L g2640 ( 
.A(n_2489),
.Y(n_2640)
);

AOI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_2470),
.A2(n_226),
.B1(n_221),
.B2(n_225),
.Y(n_2641)
);

OAI31xp33_ASAP7_75t_L g2642 ( 
.A1(n_2471),
.A2(n_228),
.A3(n_225),
.B(n_227),
.Y(n_2642)
);

AOI221xp5_ASAP7_75t_L g2643 ( 
.A1(n_2447),
.A2(n_232),
.B1(n_229),
.B2(n_231),
.C(n_233),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2564),
.A2(n_234),
.B1(n_229),
.B2(n_233),
.Y(n_2644)
);

O2A1O1Ixp5_ASAP7_75t_L g2645 ( 
.A1(n_2446),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_2645)
);

OAI32xp33_ASAP7_75t_L g2646 ( 
.A1(n_2518),
.A2(n_238),
.A3(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2526),
.B(n_238),
.Y(n_2647)
);

AOI221xp5_ASAP7_75t_L g2648 ( 
.A1(n_2438),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.C(n_242),
.Y(n_2648)
);

O2A1O1Ixp33_ASAP7_75t_SL g2649 ( 
.A1(n_2572),
.A2(n_243),
.B(n_240),
.C(n_241),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2511),
.Y(n_2650)
);

AOI322xp5_ASAP7_75t_L g2651 ( 
.A1(n_2465),
.A2(n_244),
.A3(n_245),
.B1(n_246),
.B2(n_247),
.C1(n_248),
.C2(n_250),
.Y(n_2651)
);

AOI221xp5_ASAP7_75t_L g2652 ( 
.A1(n_2467),
.A2(n_251),
.B1(n_247),
.B2(n_250),
.C(n_252),
.Y(n_2652)
);

AOI321xp33_ASAP7_75t_L g2653 ( 
.A1(n_2442),
.A2(n_252),
.A3(n_253),
.B1(n_254),
.B2(n_255),
.C(n_256),
.Y(n_2653)
);

AOI222xp33_ASAP7_75t_L g2654 ( 
.A1(n_2535),
.A2(n_253),
.B1(n_254),
.B2(n_257),
.C1(n_258),
.C2(n_259),
.Y(n_2654)
);

NAND2x1_ASAP7_75t_SL g2655 ( 
.A(n_2458),
.B(n_260),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2506),
.Y(n_2656)
);

AO22x1_ASAP7_75t_L g2657 ( 
.A1(n_2539),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_2657)
);

AOI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2485),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2532),
.Y(n_2659)
);

AOI21xp33_ASAP7_75t_SL g2660 ( 
.A1(n_2514),
.A2(n_265),
.B(n_266),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2469),
.Y(n_2661)
);

NAND2xp33_ASAP7_75t_L g2662 ( 
.A(n_2492),
.B(n_265),
.Y(n_2662)
);

AOI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2580),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_2663)
);

AOI222xp33_ASAP7_75t_L g2664 ( 
.A1(n_2469),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.C1(n_271),
.C2(n_272),
.Y(n_2664)
);

AOI221xp5_ASAP7_75t_L g2665 ( 
.A1(n_2531),
.A2(n_273),
.B1(n_269),
.B2(n_272),
.C(n_274),
.Y(n_2665)
);

OAI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2500),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_2666)
);

AOI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2542),
.A2(n_283),
.B1(n_279),
.B2(n_282),
.Y(n_2667)
);

AOI211xp5_ASAP7_75t_L g2668 ( 
.A1(n_2537),
.A2(n_286),
.B(n_279),
.C(n_285),
.Y(n_2668)
);

OAI22xp33_ASAP7_75t_L g2669 ( 
.A1(n_2497),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_2669)
);

AOI321xp33_ASAP7_75t_L g2670 ( 
.A1(n_2533),
.A2(n_287),
.A3(n_288),
.B1(n_290),
.B2(n_291),
.C(n_292),
.Y(n_2670)
);

A2O1A1Ixp33_ASAP7_75t_L g2671 ( 
.A1(n_2508),
.A2(n_295),
.B(n_288),
.C(n_291),
.Y(n_2671)
);

OAI32xp33_ASAP7_75t_L g2672 ( 
.A1(n_2569),
.A2(n_297),
.A3(n_295),
.B1(n_296),
.B2(n_298),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2655),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2586),
.Y(n_2674)
);

AOI211xp5_ASAP7_75t_L g2675 ( 
.A1(n_2585),
.A2(n_2540),
.B(n_2548),
.C(n_2541),
.Y(n_2675)
);

AOI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2662),
.A2(n_2571),
.B(n_2547),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2605),
.B(n_2538),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2640),
.A2(n_2486),
.B1(n_2454),
.B2(n_2476),
.Y(n_2678)
);

OAI211xp5_ASAP7_75t_SL g2679 ( 
.A1(n_2596),
.A2(n_2484),
.B(n_2576),
.C(n_2459),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_2589),
.Y(n_2680)
);

AOI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2632),
.A2(n_2612),
.B1(n_2606),
.B2(n_2602),
.Y(n_2681)
);

AOI21xp33_ASAP7_75t_L g2682 ( 
.A1(n_2659),
.A2(n_2480),
.B(n_2473),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2603),
.Y(n_2683)
);

CKINVDCx20_ASAP7_75t_R g2684 ( 
.A(n_2607),
.Y(n_2684)
);

HB1xp67_ASAP7_75t_L g2685 ( 
.A(n_2598),
.Y(n_2685)
);

AOI21xp33_ASAP7_75t_L g2686 ( 
.A1(n_2628),
.A2(n_2463),
.B(n_2460),
.Y(n_2686)
);

NAND2xp33_ASAP7_75t_SL g2687 ( 
.A(n_2601),
.B(n_2483),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_L g2688 ( 
.A(n_2624),
.B(n_2502),
.Y(n_2688)
);

AND3x4_ASAP7_75t_L g2689 ( 
.A(n_2617),
.B(n_2575),
.C(n_2445),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2630),
.Y(n_2690)
);

OAI22xp33_ASAP7_75t_R g2691 ( 
.A1(n_2650),
.A2(n_2633),
.B1(n_2616),
.B2(n_2593),
.Y(n_2691)
);

NOR2xp67_ASAP7_75t_L g2692 ( 
.A(n_2599),
.B(n_2505),
.Y(n_2692)
);

AOI221xp5_ASAP7_75t_L g2693 ( 
.A1(n_2597),
.A2(n_2613),
.B1(n_2660),
.B2(n_2648),
.C(n_2666),
.Y(n_2693)
);

AOI221xp5_ASAP7_75t_L g2694 ( 
.A1(n_2614),
.A2(n_2457),
.B1(n_2448),
.B2(n_2491),
.C(n_2478),
.Y(n_2694)
);

OAI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2670),
.A2(n_2530),
.B1(n_2527),
.B2(n_2479),
.C(n_2490),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2611),
.Y(n_2696)
);

OAI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2645),
.A2(n_2516),
.B(n_2523),
.Y(n_2697)
);

AOI221xp5_ASAP7_75t_L g2698 ( 
.A1(n_2621),
.A2(n_2481),
.B1(n_2495),
.B2(n_2509),
.C(n_2461),
.Y(n_2698)
);

XNOR2x1_ASAP7_75t_L g2699 ( 
.A(n_2657),
.B(n_2504),
.Y(n_2699)
);

AOI211xp5_ASAP7_75t_L g2700 ( 
.A1(n_2669),
.A2(n_2515),
.B(n_2488),
.C(n_2462),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2653),
.B(n_2636),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2631),
.Y(n_2702)
);

HB1xp67_ASAP7_75t_L g2703 ( 
.A(n_2587),
.Y(n_2703)
);

OAI211xp5_ASAP7_75t_SL g2704 ( 
.A1(n_2643),
.A2(n_2513),
.B(n_2555),
.C(n_2464),
.Y(n_2704)
);

XOR2x2_ASAP7_75t_L g2705 ( 
.A(n_2658),
.B(n_2525),
.Y(n_2705)
);

AOI221xp5_ASAP7_75t_L g2706 ( 
.A1(n_2656),
.A2(n_2594),
.B1(n_2652),
.B2(n_2649),
.C(n_2637),
.Y(n_2706)
);

AOI31xp33_ASAP7_75t_L g2707 ( 
.A1(n_2627),
.A2(n_2521),
.A3(n_2451),
.B(n_2510),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2647),
.Y(n_2708)
);

OAI22xp5_ASAP7_75t_L g2709 ( 
.A1(n_2663),
.A2(n_2496),
.B1(n_2524),
.B2(n_2512),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2604),
.A2(n_2501),
.B1(n_2466),
.B2(n_2499),
.Y(n_2710)
);

AOI22xp5_ASAP7_75t_SL g2711 ( 
.A1(n_2638),
.A2(n_2455),
.B1(n_2468),
.B2(n_2475),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_2588),
.B(n_2558),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2590),
.A2(n_2503),
.B1(n_2477),
.B2(n_2517),
.Y(n_2713)
);

AOI22xp33_ASAP7_75t_L g2714 ( 
.A1(n_2608),
.A2(n_2482),
.B1(n_1115),
.B2(n_1141),
.Y(n_2714)
);

OAI21xp33_ASAP7_75t_L g2715 ( 
.A1(n_2623),
.A2(n_300),
.B(n_301),
.Y(n_2715)
);

NAND2xp33_ASAP7_75t_SL g2716 ( 
.A(n_2629),
.B(n_301),
.Y(n_2716)
);

AOI221x1_ASAP7_75t_SL g2717 ( 
.A1(n_2591),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.C(n_306),
.Y(n_2717)
);

XNOR2xp5_ASAP7_75t_L g2718 ( 
.A(n_2668),
.B(n_302),
.Y(n_2718)
);

NOR2x1_ASAP7_75t_L g2719 ( 
.A(n_2635),
.B(n_2600),
.Y(n_2719)
);

OAI221xp5_ASAP7_75t_L g2720 ( 
.A1(n_2642),
.A2(n_307),
.B1(n_304),
.B2(n_306),
.C(n_308),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2595),
.B(n_307),
.Y(n_2721)
);

AOI221xp5_ASAP7_75t_L g2722 ( 
.A1(n_2615),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.C(n_312),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2619),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2667),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2672),
.Y(n_2725)
);

AOI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2639),
.A2(n_313),
.B(n_314),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2671),
.Y(n_2727)
);

A2O1A1Ixp33_ASAP7_75t_SL g2728 ( 
.A1(n_2661),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_2728)
);

OAI21xp5_ASAP7_75t_SL g2729 ( 
.A1(n_2641),
.A2(n_317),
.B(n_318),
.Y(n_2729)
);

AOI21xp33_ASAP7_75t_L g2730 ( 
.A1(n_2642),
.A2(n_318),
.B(n_319),
.Y(n_2730)
);

NAND4xp25_ASAP7_75t_L g2731 ( 
.A(n_2681),
.B(n_2665),
.C(n_2620),
.D(n_2618),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2685),
.Y(n_2732)
);

OAI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2684),
.A2(n_2622),
.B1(n_2609),
.B2(n_2634),
.Y(n_2733)
);

XNOR2xp5_ASAP7_75t_L g2734 ( 
.A(n_2689),
.B(n_2644),
.Y(n_2734)
);

XOR2xp5_ASAP7_75t_L g2735 ( 
.A(n_2718),
.B(n_2610),
.Y(n_2735)
);

AOI22xp5_ASAP7_75t_L g2736 ( 
.A1(n_2690),
.A2(n_2654),
.B1(n_2592),
.B2(n_2625),
.Y(n_2736)
);

OAI31xp33_ASAP7_75t_L g2737 ( 
.A1(n_2674),
.A2(n_2664),
.A3(n_2646),
.B(n_2651),
.Y(n_2737)
);

AOI211xp5_ASAP7_75t_L g2738 ( 
.A1(n_2691),
.A2(n_2626),
.B(n_321),
.C(n_319),
.Y(n_2738)
);

AOI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2680),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_2739)
);

AOI221xp5_ASAP7_75t_L g2740 ( 
.A1(n_2707),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.C(n_325),
.Y(n_2740)
);

AOI31xp33_ASAP7_75t_L g2741 ( 
.A1(n_2703),
.A2(n_326),
.A3(n_323),
.B(n_325),
.Y(n_2741)
);

AOI211xp5_ASAP7_75t_SL g2742 ( 
.A1(n_2675),
.A2(n_330),
.B(n_327),
.C(n_329),
.Y(n_2742)
);

NOR2x1p5_ASAP7_75t_L g2743 ( 
.A(n_2702),
.B(n_327),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2683),
.Y(n_2744)
);

OAI21xp5_ASAP7_75t_L g2745 ( 
.A1(n_2676),
.A2(n_329),
.B(n_330),
.Y(n_2745)
);

AOI321xp33_ASAP7_75t_L g2746 ( 
.A1(n_2673),
.A2(n_331),
.A3(n_332),
.B1(n_333),
.B2(n_334),
.C(n_336),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2708),
.A2(n_1115),
.B1(n_1141),
.B2(n_1121),
.Y(n_2747)
);

AO22x2_ASAP7_75t_L g2748 ( 
.A1(n_2696),
.A2(n_2725),
.B1(n_2699),
.B2(n_2727),
.Y(n_2748)
);

NAND2x1_ASAP7_75t_L g2749 ( 
.A(n_2692),
.B(n_331),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2693),
.B(n_332),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2701),
.B(n_333),
.Y(n_2751)
);

OAI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2695),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2677),
.Y(n_2753)
);

A2O1A1Ixp33_ASAP7_75t_L g2754 ( 
.A1(n_2688),
.A2(n_340),
.B(n_337),
.C(n_339),
.Y(n_2754)
);

NOR2x1p5_ASAP7_75t_L g2755 ( 
.A(n_2721),
.B(n_340),
.Y(n_2755)
);

OAI31xp33_ASAP7_75t_L g2756 ( 
.A1(n_2716),
.A2(n_344),
.A3(n_341),
.B(n_342),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2705),
.Y(n_2757)
);

AOI21xp5_ASAP7_75t_L g2758 ( 
.A1(n_2687),
.A2(n_342),
.B(n_345),
.Y(n_2758)
);

AO22x2_ASAP7_75t_L g2759 ( 
.A1(n_2724),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_2759)
);

AOI22xp33_ASAP7_75t_L g2760 ( 
.A1(n_2682),
.A2(n_1115),
.B1(n_1141),
.B2(n_1121),
.Y(n_2760)
);

OAI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2678),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_2761)
);

AOI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2709),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_2762)
);

NOR2xp67_ASAP7_75t_SL g2763 ( 
.A(n_2720),
.B(n_350),
.Y(n_2763)
);

INVxp67_ASAP7_75t_L g2764 ( 
.A(n_2719),
.Y(n_2764)
);

AOI221xp5_ASAP7_75t_L g2765 ( 
.A1(n_2730),
.A2(n_351),
.B1(n_353),
.B2(n_355),
.C(n_356),
.Y(n_2765)
);

OAI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2713),
.A2(n_359),
.B1(n_355),
.B2(n_357),
.Y(n_2766)
);

NOR2x1_ASAP7_75t_L g2767 ( 
.A(n_2732),
.B(n_2679),
.Y(n_2767)
);

NOR2xp67_ASAP7_75t_L g2768 ( 
.A(n_2744),
.B(n_2726),
.Y(n_2768)
);

OAI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2753),
.A2(n_2722),
.B1(n_2706),
.B2(n_2710),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2764),
.Y(n_2770)
);

NOR2x1_ASAP7_75t_L g2771 ( 
.A(n_2731),
.B(n_2729),
.Y(n_2771)
);

NOR2x1_ASAP7_75t_L g2772 ( 
.A(n_2745),
.B(n_2723),
.Y(n_2772)
);

INVxp67_ASAP7_75t_L g2773 ( 
.A(n_2759),
.Y(n_2773)
);

AO22x2_ASAP7_75t_L g2774 ( 
.A1(n_2749),
.A2(n_2697),
.B1(n_2712),
.B2(n_2717),
.Y(n_2774)
);

INVxp67_ASAP7_75t_L g2775 ( 
.A(n_2759),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2748),
.Y(n_2776)
);

AOI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2751),
.A2(n_2712),
.B1(n_2694),
.B2(n_2715),
.Y(n_2777)
);

NOR2x1_ASAP7_75t_L g2778 ( 
.A(n_2741),
.B(n_2704),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2743),
.B(n_2728),
.Y(n_2779)
);

INVx3_ASAP7_75t_L g2780 ( 
.A(n_2748),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2742),
.B(n_2700),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2735),
.B(n_2711),
.Y(n_2782)
);

AO22x1_ASAP7_75t_L g2783 ( 
.A1(n_2752),
.A2(n_2700),
.B1(n_2686),
.B2(n_2714),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2746),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2755),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2736),
.A2(n_2698),
.B1(n_361),
.B2(n_357),
.Y(n_2786)
);

OR2x2_ASAP7_75t_L g2787 ( 
.A(n_2780),
.B(n_2758),
.Y(n_2787)
);

AOI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2770),
.A2(n_2733),
.B1(n_2757),
.B2(n_2766),
.Y(n_2788)
);

INVx2_ASAP7_75t_SL g2789 ( 
.A(n_2774),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2774),
.Y(n_2790)
);

NOR2x1_ASAP7_75t_L g2791 ( 
.A(n_2767),
.B(n_2776),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2768),
.B(n_2738),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2779),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2778),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2781),
.Y(n_2795)
);

NOR2x1_ASAP7_75t_L g2796 ( 
.A(n_2769),
.B(n_2761),
.Y(n_2796)
);

NOR2x1_ASAP7_75t_SL g2797 ( 
.A(n_2784),
.B(n_2750),
.Y(n_2797)
);

XOR2x1_ASAP7_75t_L g2798 ( 
.A(n_2785),
.B(n_2734),
.Y(n_2798)
);

NAND4xp75_ASAP7_75t_L g2799 ( 
.A(n_2782),
.B(n_2737),
.C(n_2756),
.D(n_2765),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2773),
.B(n_2754),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2775),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2771),
.Y(n_2802)
);

OR2x2_ASAP7_75t_L g2803 ( 
.A(n_2786),
.B(n_2762),
.Y(n_2803)
);

OAI221xp5_ASAP7_75t_L g2804 ( 
.A1(n_2789),
.A2(n_2777),
.B1(n_2772),
.B2(n_2740),
.C(n_2747),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2793),
.A2(n_2763),
.B1(n_2739),
.B2(n_2783),
.Y(n_2805)
);

OAI221xp5_ASAP7_75t_L g2806 ( 
.A1(n_2794),
.A2(n_2760),
.B1(n_362),
.B2(n_363),
.C(n_364),
.Y(n_2806)
);

NAND4xp25_ASAP7_75t_L g2807 ( 
.A(n_2791),
.B(n_364),
.C(n_360),
.D(n_362),
.Y(n_2807)
);

OAI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2790),
.A2(n_365),
.B(n_367),
.Y(n_2808)
);

AND3x4_ASAP7_75t_L g2809 ( 
.A(n_2796),
.B(n_2795),
.C(n_2798),
.Y(n_2809)
);

AOI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2801),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_2810)
);

OAI221xp5_ASAP7_75t_L g2811 ( 
.A1(n_2802),
.A2(n_368),
.B1(n_371),
.B2(n_372),
.C(n_373),
.Y(n_2811)
);

NAND3xp33_ASAP7_75t_SL g2812 ( 
.A(n_2788),
.B(n_371),
.C(n_374),
.Y(n_2812)
);

OAI221xp5_ASAP7_75t_L g2813 ( 
.A1(n_2787),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.C(n_378),
.Y(n_2813)
);

AOI221xp5_ASAP7_75t_L g2814 ( 
.A1(n_2792),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.C(n_382),
.Y(n_2814)
);

OAI322xp33_ASAP7_75t_L g2815 ( 
.A1(n_2800),
.A2(n_380),
.A3(n_381),
.B1(n_382),
.B2(n_384),
.C1(n_385),
.C2(n_387),
.Y(n_2815)
);

AOI211xp5_ASAP7_75t_L g2816 ( 
.A1(n_2803),
.A2(n_384),
.B(n_387),
.C(n_389),
.Y(n_2816)
);

AO22x2_ASAP7_75t_L g2817 ( 
.A1(n_2799),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_2817)
);

OAI321xp33_ASAP7_75t_L g2818 ( 
.A1(n_2797),
.A2(n_391),
.A3(n_393),
.B1(n_394),
.B2(n_395),
.C(n_396),
.Y(n_2818)
);

AOI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2799),
.A2(n_394),
.B1(n_395),
.B2(n_397),
.Y(n_2819)
);

OAI221xp5_ASAP7_75t_L g2820 ( 
.A1(n_2789),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.C(n_400),
.Y(n_2820)
);

OAI221xp5_ASAP7_75t_L g2821 ( 
.A1(n_2789),
.A2(n_398),
.B1(n_400),
.B2(n_401),
.C(n_402),
.Y(n_2821)
);

NOR3xp33_ASAP7_75t_L g2822 ( 
.A(n_2791),
.B(n_401),
.C(n_402),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2817),
.Y(n_2823)
);

NAND3xp33_ASAP7_75t_L g2824 ( 
.A(n_2822),
.B(n_1115),
.C(n_403),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2818),
.B(n_403),
.Y(n_2825)
);

NAND2x1p5_ASAP7_75t_L g2826 ( 
.A(n_2805),
.B(n_405),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2817),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2809),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2819),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2816),
.B(n_406),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2820),
.Y(n_2831)
);

OAI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2808),
.A2(n_406),
.B(n_407),
.Y(n_2832)
);

HB1xp67_ASAP7_75t_L g2833 ( 
.A(n_2807),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2810),
.B(n_408),
.Y(n_2834)
);

NAND3xp33_ASAP7_75t_L g2835 ( 
.A(n_2804),
.B(n_409),
.C(n_410),
.Y(n_2835)
);

NOR2xp67_ASAP7_75t_L g2836 ( 
.A(n_2821),
.B(n_409),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2812),
.A2(n_1156),
.B1(n_1153),
.B2(n_1141),
.Y(n_2837)
);

OA22x2_ASAP7_75t_L g2838 ( 
.A1(n_2813),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2815),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2811),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2806),
.Y(n_2841)
);

OR2x2_ASAP7_75t_L g2842 ( 
.A(n_2814),
.B(n_411),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2817),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2828),
.A2(n_413),
.B1(n_414),
.B2(n_415),
.Y(n_2844)
);

AND2x2_ASAP7_75t_SL g2845 ( 
.A(n_2827),
.B(n_413),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2823),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2823),
.Y(n_2847)
);

INVx4_ASAP7_75t_L g2848 ( 
.A(n_2826),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2839),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2843),
.B(n_417),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2833),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2836),
.B(n_2837),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2838),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2829),
.B(n_420),
.Y(n_2854)
);

NOR2xp67_ASAP7_75t_L g2855 ( 
.A(n_2835),
.B(n_420),
.Y(n_2855)
);

XOR2xp5_ASAP7_75t_L g2856 ( 
.A(n_2841),
.B(n_421),
.Y(n_2856)
);

AND2x4_ASAP7_75t_L g2857 ( 
.A(n_2831),
.B(n_422),
.Y(n_2857)
);

NAND2xp33_ASAP7_75t_SL g2858 ( 
.A(n_2830),
.B(n_424),
.Y(n_2858)
);

AOI221xp5_ASAP7_75t_L g2859 ( 
.A1(n_2846),
.A2(n_2825),
.B1(n_2824),
.B2(n_2832),
.C(n_2840),
.Y(n_2859)
);

AOI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2851),
.A2(n_2834),
.B1(n_2842),
.B2(n_426),
.Y(n_2860)
);

AOI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2847),
.A2(n_424),
.B1(n_425),
.B2(n_427),
.Y(n_2861)
);

INVx3_ASAP7_75t_L g2862 ( 
.A(n_2848),
.Y(n_2862)
);

OAI21x1_ASAP7_75t_L g2863 ( 
.A1(n_2850),
.A2(n_425),
.B(n_428),
.Y(n_2863)
);

INVx4_ASAP7_75t_L g2864 ( 
.A(n_2857),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2845),
.Y(n_2865)
);

CKINVDCx20_ASAP7_75t_R g2866 ( 
.A(n_2858),
.Y(n_2866)
);

NOR2x1_ASAP7_75t_L g2867 ( 
.A(n_2854),
.B(n_428),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2856),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2853),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2855),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2852),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2849),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2862),
.B(n_2844),
.Y(n_2873)
);

AOI21xp33_ASAP7_75t_SL g2874 ( 
.A1(n_2869),
.A2(n_429),
.B(n_430),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2865),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2867),
.Y(n_2876)
);

OR2x2_ASAP7_75t_L g2877 ( 
.A(n_2864),
.B(n_430),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2863),
.Y(n_2878)
);

AO22x2_ASAP7_75t_L g2879 ( 
.A1(n_2870),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_2879)
);

OAI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2871),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_2880)
);

XNOR2x1_ASAP7_75t_SL g2881 ( 
.A(n_2868),
.B(n_434),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2866),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2872),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2860),
.B(n_434),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2859),
.B(n_435),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2861),
.B(n_435),
.Y(n_2886)
);

AOI21xp33_ASAP7_75t_L g2887 ( 
.A1(n_2871),
.A2(n_436),
.B(n_437),
.Y(n_2887)
);

OR2x6_ASAP7_75t_L g2888 ( 
.A(n_2864),
.B(n_438),
.Y(n_2888)
);

OAI22x1_ASAP7_75t_SL g2889 ( 
.A1(n_2876),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_2889)
);

OAI22xp5_ASAP7_75t_L g2890 ( 
.A1(n_2882),
.A2(n_441),
.B1(n_443),
.B2(n_444),
.Y(n_2890)
);

INVxp67_ASAP7_75t_SL g2891 ( 
.A(n_2881),
.Y(n_2891)
);

AOI22x1_ASAP7_75t_L g2892 ( 
.A1(n_2873),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.Y(n_2892)
);

CKINVDCx20_ASAP7_75t_R g2893 ( 
.A(n_2883),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2877),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2888),
.Y(n_2895)
);

HB1xp67_ASAP7_75t_L g2896 ( 
.A(n_2888),
.Y(n_2896)
);

AO22x2_ASAP7_75t_L g2897 ( 
.A1(n_2878),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2875),
.B(n_447),
.Y(n_2898)
);

OAI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2885),
.A2(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_2899)
);

OAI22x1_ASAP7_75t_SL g2900 ( 
.A1(n_2884),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_2900)
);

AOI22x1_ASAP7_75t_L g2901 ( 
.A1(n_2891),
.A2(n_2879),
.B1(n_2874),
.B2(n_2887),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2896),
.A2(n_2886),
.B(n_2880),
.Y(n_2902)
);

OAI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2893),
.A2(n_451),
.B(n_452),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2897),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2894),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2895),
.A2(n_2898),
.B(n_2899),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2892),
.Y(n_2907)
);

OAI21x1_ASAP7_75t_L g2908 ( 
.A1(n_2890),
.A2(n_452),
.B(n_454),
.Y(n_2908)
);

OAI21xp33_ASAP7_75t_L g2909 ( 
.A1(n_2900),
.A2(n_454),
.B(n_456),
.Y(n_2909)
);

OAI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2889),
.A2(n_457),
.B1(n_459),
.B2(n_460),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2891),
.B(n_459),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2905),
.A2(n_461),
.B(n_462),
.Y(n_2912)
);

INVxp67_ASAP7_75t_L g2913 ( 
.A(n_2904),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2902),
.A2(n_461),
.B(n_462),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2911),
.A2(n_464),
.B(n_466),
.Y(n_2915)
);

AOI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2910),
.A2(n_464),
.B1(n_468),
.B2(n_469),
.Y(n_2916)
);

OA21x2_ASAP7_75t_L g2917 ( 
.A1(n_2906),
.A2(n_468),
.B(n_469),
.Y(n_2917)
);

HB1xp67_ASAP7_75t_L g2918 ( 
.A(n_2901),
.Y(n_2918)
);

AO21x2_ASAP7_75t_L g2919 ( 
.A1(n_2909),
.A2(n_470),
.B(n_472),
.Y(n_2919)
);

AOI22xp33_ASAP7_75t_L g2920 ( 
.A1(n_2907),
.A2(n_470),
.B1(n_472),
.B2(n_474),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2903),
.A2(n_474),
.B(n_475),
.Y(n_2921)
);

OAI222xp33_ASAP7_75t_L g2922 ( 
.A1(n_2913),
.A2(n_2918),
.B1(n_2916),
.B2(n_2914),
.C1(n_2915),
.C2(n_2921),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2917),
.A2(n_2908),
.B1(n_477),
.B2(n_478),
.Y(n_2923)
);

AOI222xp33_ASAP7_75t_SL g2924 ( 
.A1(n_2919),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.C1(n_479),
.C2(n_481),
.Y(n_2924)
);

AOI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2912),
.A2(n_476),
.B1(n_479),
.B2(n_483),
.Y(n_2925)
);

AOI221xp5_ASAP7_75t_L g2926 ( 
.A1(n_2920),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.C(n_486),
.Y(n_2926)
);

AOI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2924),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_2927)
);

AOI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2923),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_2928)
);

AO22x2_ASAP7_75t_L g2929 ( 
.A1(n_2928),
.A2(n_2922),
.B1(n_2925),
.B2(n_2926),
.Y(n_2929)
);

O2A1O1Ixp33_ASAP7_75t_L g2930 ( 
.A1(n_2929),
.A2(n_2927),
.B(n_491),
.C(n_492),
.Y(n_2930)
);

AOI211xp5_ASAP7_75t_L g2931 ( 
.A1(n_2930),
.A2(n_490),
.B(n_491),
.C(n_492),
.Y(n_2931)
);


endmodule