module fake_jpeg_5223_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx14_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_8),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_30),
.B1(n_33),
.B2(n_18),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_21),
.B1(n_10),
.B2(n_12),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_21),
.B1(n_9),
.B2(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_40),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_20),
.B(n_11),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_36),
.B1(n_29),
.B2(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_39),
.B(n_44),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_46),
.B1(n_29),
.B2(n_38),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_35),
.B1(n_41),
.B2(n_13),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_47),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_50),
.B1(n_31),
.B2(n_17),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.C(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);


endmodule