module fake_netlist_6_127_n_6525 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_6525);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_6525;

wire n_5643;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_6441;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_6141;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_5653;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_677;
wire n_6126;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_2179;
wire n_5963;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_5950;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_3030;
wire n_830;
wire n_5838;
wire n_5725;
wire n_6324;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_6325;
wire n_4724;
wire n_945;
wire n_5598;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_5819;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_6280;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_5930;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_5908;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_6243;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_6374;
wire n_2843;
wire n_3760;
wire n_6015;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_5638;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_6323;
wire n_6110;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_6371;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_5684;
wire n_5729;
wire n_6404;
wire n_5680;
wire n_6148;
wire n_686;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_5902;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_6196;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_6485;
wire n_6107;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_1075;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_6282;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_6383;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_6151;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_6431;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_6055;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_5897;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3875;
wire n_3012;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_5922;
wire n_2641;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_5667;
wire n_780;
wire n_2624;
wire n_5865;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_6248;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_5795;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_5226;
wire n_687;
wire n_890;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_6010;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_6185;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_6042;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_5957;
wire n_4228;
wire n_3423;
wire n_6357;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_2767;
wire n_963;
wire n_6509;
wire n_4576;
wire n_5929;
wire n_4615;
wire n_5787;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_6033;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_6097;
wire n_6369;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_4310;
wire n_6359;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_5811;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_5901;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_648;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_6519;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_6402;
wire n_4551;
wire n_2857;
wire n_6195;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_6149;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_6414;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_6264;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_5741;
wire n_2773;
wire n_6205;
wire n_6380;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_6449;
wire n_2797;
wire n_6440;
wire n_4746;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_5952;
wire n_3964;
wire n_2416;
wire n_5947;
wire n_1877;
wire n_3944;
wire n_6124;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_5985;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_5761;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_6382;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_2146;
wire n_2131;
wire n_5472;
wire n_3547;
wire n_5679;
wire n_2575;
wire n_5100;
wire n_5973;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_6339;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_6417;
wire n_5740;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_858;
wire n_5182;
wire n_956;
wire n_5534;
wire n_663;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_664;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_6199;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_6471;
wire n_2448;
wire n_5949;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_6478;
wire n_3406;
wire n_820;
wire n_951;
wire n_6100;
wire n_6516;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_6522;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_5906;
wire n_1934;
wire n_628;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_6024;
wire n_807;
wire n_4761;
wire n_6270;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_5783;
wire n_6207;
wire n_3120;
wire n_5821;
wire n_6245;
wire n_6079;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_5556;
wire n_4932;
wire n_5456;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_6427;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_6412;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_6437;
wire n_3195;
wire n_2526;
wire n_6346;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_6059;
wire n_3042;
wire n_6065;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_6075;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_6117;
wire n_5618;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_6494;
wire n_6133;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_6453;
wire n_5978;
wire n_4996;
wire n_4990;
wire n_5247;
wire n_6127;
wire n_4398;
wire n_2498;
wire n_6217;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_6006;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_5689;
wire n_1043;
wire n_4090;
wire n_6115;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_6048;
wire n_4144;
wire n_6416;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_5931;
wire n_2371;
wire n_6139;
wire n_1361;
wire n_662;
wire n_6256;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_1642;
wire n_3210;
wire n_6361;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_6085;
wire n_5731;
wire n_6329;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_6370;
wire n_2518;
wire n_5883;
wire n_5754;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_6147;
wire n_2852;
wire n_1524;
wire n_6448;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_5934;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_6157;
wire n_4859;
wire n_2626;
wire n_5880;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_5960;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_6397;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_6073;
wire n_1484;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_6405;
wire n_5149;
wire n_5571;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_6206;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_6363;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_6290;
wire n_6025;
wire n_1337;
wire n_1477;
wire n_6455;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5607;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_5999;
wire n_4376;
wire n_6203;
wire n_1001;
wire n_6408;
wire n_2241;
wire n_6150;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_695;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_6401;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_5911;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_5577;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_6392;
wire n_1810;
wire n_5915;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_5779;
wire n_1643;
wire n_2020;
wire n_6260;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_6286;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_3617;
wire n_2076;
wire n_6019;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_6214;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_6036;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_1944;
wire n_6403;
wire n_1347;
wire n_795;
wire n_1221;
wire n_6013;
wire n_1245;
wire n_3215;
wire n_6491;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_6348;
wire n_1561;
wire n_1112;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_6293;
wire n_5847;
wire n_6049;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_668;
wire n_4166;
wire n_1821;
wire n_6136;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_5541;
wire n_5568;
wire n_6312;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_5723;
wire n_5918;
wire n_3468;
wire n_6388;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_5696;
wire n_4486;
wire n_1816;
wire n_6131;
wire n_5848;
wire n_3024;
wire n_4612;
wire n_6435;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_6351;
wire n_5163;
wire n_6212;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_5485;
wire n_5823;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_6334;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_3552;
wire n_941;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_6429;
wire n_6407;
wire n_4091;
wire n_1753;
wire n_6389;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_633;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_6113;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_3896;
wire n_3815;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_722;
wire n_5613;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_629;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_6278;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_5581;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_6200;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_6373;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_5601;
wire n_5784;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_6411;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_6381;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_6265;
wire n_2989;
wire n_5778;
wire n_3395;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_6135;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_2356;
wire n_1511;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_5788;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_641;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_6168;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_6450;
wire n_3261;
wire n_666;
wire n_4187;
wire n_6309;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_5942;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_6300;
wire n_3532;
wire n_5716;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_6179;
wire n_6395;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_659;
wire n_3351;
wire n_6171;
wire n_808;
wire n_5519;
wire n_4047;
wire n_6269;
wire n_5753;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_6083;
wire n_3164;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5808;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_6120;
wire n_6068;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_6423;
wire n_2850;
wire n_6342;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_3883;
wire n_5961;
wire n_5866;
wire n_3728;
wire n_6507;
wire n_2925;
wire n_4499;
wire n_6399;
wire n_5822;
wire n_5195;
wire n_6121;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_5533;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_5953;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_6459;
wire n_1663;
wire n_6505;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_6001;
wire n_3686;
wire n_4502;
wire n_5958;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_5792;
wire n_3581;
wire n_3069;
wire n_6183;
wire n_6023;
wire n_6258;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_5554;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_5553;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_5790;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_6186;
wire n_816;
wire n_6210;
wire n_6500;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_6163;
wire n_5972;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_5757;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_637;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_5488;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_5637;
wire n_1987;
wire n_6452;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_5843;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_6355;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_6227;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_6468;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_6442;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_6499;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_631;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_5887;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_6276;
wire n_5631;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_6008;
wire n_1022;
wire n_6420;
wire n_5854;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_5686;
wire n_5899;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_6447;
wire n_4264;
wire n_5981;
wire n_3788;
wire n_4891;
wire n_5937;
wire n_777;
wire n_6422;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_6040;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_6460;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_6160;
wire n_796;
wire n_1195;
wire n_6192;
wire n_1811;
wire n_6368;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_6039;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_5721;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_6012;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_6064;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_6275;
wire n_1564;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_5893;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_6277;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_1220;
wire n_6051;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_6487;
wire n_5121;
wire n_6026;
wire n_6070;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_5589;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_6481;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_6341;
wire n_6384;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_5475;
wire n_5807;
wire n_4448;
wire n_1096;
wire n_6233;
wire n_2227;
wire n_6377;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_6257;
wire n_2159;
wire n_688;
wire n_2315;
wire n_4132;
wire n_4386;
wire n_1077;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_5936;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_856;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_6069;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_5187;
wire n_5875;
wire n_4024;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_732;
wire n_2983;
wire n_6335;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_6252;
wire n_1871;
wire n_4860;
wire n_6211;
wire n_845;
wire n_5844;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_6164;
wire n_768;
wire n_6173;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_2598;
wire n_1916;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_6189;
wire n_1206;
wire n_4016;
wire n_5867;
wire n_750;
wire n_5508;
wire n_4656;
wire n_6479;
wire n_3839;
wire n_2823;
wire n_6410;
wire n_6158;
wire n_5597;
wire n_4915;
wire n_4328;
wire n_6413;
wire n_6090;
wire n_1057;
wire n_6506;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_5862;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_6234;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_5980;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_6430;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5987;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5988;
wire n_5585;
wire n_6058;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_6190;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_6249;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_624;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_936;
wire n_885;
wire n_6161;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_5904;
wire n_4739;
wire n_6062;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_6482;
wire n_4128;
wire n_6294;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_5503;
wire n_5845;
wire n_5945;
wire n_804;
wire n_2390;
wire n_6246;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_5755;
wire n_5600;
wire n_707;
wire n_1900;
wire n_5048;
wire n_6053;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_6123;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_5749;
wire n_1672;
wire n_6271;
wire n_6489;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_5993;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_6521;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_6162;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_6198;
wire n_4269;
wire n_5418;
wire n_6178;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_1019;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_6458;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_6315;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_6262;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_6319;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_6175;
wire n_3806;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_5909;
wire n_671;
wire n_6093;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_6099;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_6321;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_5890;
wire n_6415;
wire n_6465;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_676;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_5891;
wire n_3541;
wire n_6101;
wire n_3117;
wire n_5935;
wire n_4930;
wire n_5623;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_5990;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_6281;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_6311;
wire n_930;
wire n_2620;
wire n_5162;
wire n_6134;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_653;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_626;
wire n_990;
wire n_6231;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_6443;
wire n_5709;
wire n_1693;
wire n_6446;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_6337;
wire n_3643;
wire n_6181;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_5799;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_5266;
wire n_5580;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_6310;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_5764;
wire n_2282;
wire n_6365;
wire n_4628;
wire n_2047;
wire n_6229;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_635;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_6177;
wire n_1996;
wire n_6332;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_5982;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_5917;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_6116;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5561;
wire n_5410;
wire n_2215;
wire n_6167;
wire n_1884;
wire n_6170;
wire n_665;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_6307;
wire n_632;
wire n_6094;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_6155;
wire n_6267;
wire n_1833;
wire n_3903;
wire n_5998;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_6028;
wire n_1417;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_5916;
wire n_681;
wire n_4648;
wire n_3094;
wire n_6299;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_5691;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_6316;
wire n_6292;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_6220;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_1003;
wire n_5713;
wire n_5256;
wire n_6318;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_5550;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_6366;
wire n_6230;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_6391;
wire n_5659;
wire n_3619;
wire n_1415;
wire n_5881;
wire n_1370;
wire n_1786;
wire n_6473;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_6483;
wire n_1803;
wire n_4065;
wire n_5863;
wire n_2645;
wire n_3904;
wire n_1517;
wire n_1867;
wire n_1393;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_5955;
wire n_658;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_6076;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_758;
wire n_5851;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_6390;
wire n_5796;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_6297;
wire n_6523;
wire n_6096;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_638;
wire n_1404;
wire n_5492;
wire n_5995;
wire n_2378;
wire n_887;
wire n_5905;
wire n_2655;
wire n_4600;
wire n_6193;
wire n_6501;
wire n_1467;
wire n_4250;
wire n_5829;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_5525;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_6052;
wire n_2907;
wire n_5374;
wire n_5575;
wire n_1843;
wire n_5675;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_6240;
wire n_6347;
wire n_5020;
wire n_6511;
wire n_5297;
wire n_1309;
wire n_1123;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_1970;
wire n_6358;
wire n_630;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_5959;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_6396;
wire n_5642;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_6109;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_689;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_692;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_5885;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_1312;
wire n_5668;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_1165;
wire n_5892;
wire n_4773;
wire n_5654;
wire n_2008;
wire n_6009;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_5923;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_690;
wire n_5692;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_6066;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_696;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_6296;
wire n_4055;
wire n_2178;
wire n_5968;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_6497;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_6470;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_6187;
wire n_678;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_6409;
wire n_1634;
wire n_3252;
wire n_627;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_6130;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_5976;
wire n_3128;
wire n_1527;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_5690;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_5801;
wire n_6047;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_6354;
wire n_3608;
wire n_4540;
wire n_6344;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_3499;
wire n_4284;
wire n_6305;
wire n_1005;
wire n_1947;
wire n_6209;
wire n_3426;
wire n_4971;
wire n_5656;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_2650;
wire n_5652;
wire n_6457;
wire n_987;
wire n_5499;
wire n_720;
wire n_3348;
wire n_3229;
wire n_1707;
wire n_656;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_684;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_6466;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_5442;
wire n_6386;
wire n_5948;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_6208;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_6438;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_6291;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_5584;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_6469;
wire n_2682;
wire n_3032;
wire n_6223;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_5497;
wire n_880;
wire n_6464;
wire n_6356;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_5964;
wire n_6004;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_6272;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_5467;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_6222;
wire n_1093;
wire n_1783;
wire n_6268;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_6456;
wire n_651;
wire n_3407;
wire n_5992;
wire n_5313;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_6467;
wire n_5079;
wire n_1453;
wire n_6336;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_5592;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_5157;
wire n_2100;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_5708;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_6298;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_6421;
wire n_1905;
wire n_3466;
wire n_762;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_6328;
wire n_5956;
wire n_5287;
wire n_6236;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_6007;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_6144;
wire n_3338;
wire n_4217;
wire n_6197;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_6247;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_3572;
wire n_3886;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_6242;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_6285;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_5677;
wire n_4124;
wire n_5570;
wire n_6418;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5927;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_6400;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_6398;
wire n_5486;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_5889;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_5849;
wire n_4554;
wire n_6224;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_6092;
wire n_5951;
wire n_6241;
wire n_1692;
wire n_1084;
wire n_5912;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_650;
wire n_6165;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_5910;
wire n_5895;
wire n_1041;
wire n_5804;
wire n_3134;
wire n_5965;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5682;
wire n_5387;
wire n_654;
wire n_5557;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_5681;
wire n_6119;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4145;
wire n_4821;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_5703;
wire n_833;
wire n_6320;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_6202;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_652;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_5979;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_6044;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_6125;
wire n_655;
wire n_4726;
wire n_1045;
wire n_5907;
wire n_786;
wire n_1559;
wire n_6045;
wire n_1872;
wire n_5040;
wire n_6063;
wire n_1325;
wire n_6504;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_6154;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_5977;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_6003;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_6031;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_6060;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_680;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_1953;
wire n_6191;
wire n_4741;
wire n_6172;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_643;
wire n_5842;
wire n_5814;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_6215;
wire n_3231;
wire n_789;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_6517;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_6088;
wire n_5777;
wire n_4225;
wire n_747;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_6393;
wire n_5064;
wire n_5610;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_6035;
wire n_957;
wire n_1994;
wire n_2566;
wire n_6364;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_6114;
wire n_4568;
wire n_1205;
wire n_6061;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_6253;
wire n_2914;
wire n_5786;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_1016;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_6419;
wire n_1083;
wire n_5768;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_1721;
wire n_3494;
wire n_6244;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_5872;
wire n_5858;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_6338;
wire n_5700;
wire n_1500;
wire n_6037;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_5874;
wire n_6266;
wire n_6488;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_5873;
wire n_1085;
wire n_2042;
wire n_771;
wire n_6317;
wire n_924;
wire n_1582;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_6480;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_4845;
wire n_2033;
wire n_4104;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_6176;
wire n_2174;
wire n_6367;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_6080;
wire n_4865;
wire n_1039;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_6056;
wire n_5832;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_4522;
wire n_967;
wire n_2001;
wire n_4341;
wire n_679;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_5971;
wire n_6327;
wire n_812;
wire n_6145;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_5933;
wire n_1888;
wire n_6204;
wire n_1311;
wire n_4780;
wire n_670;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_6451;
wire n_3039;
wire n_1226;
wire n_6514;
wire n_3740;
wire n_5996;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_640;
wire n_1322;
wire n_1958;
wire n_5903;
wire n_5986;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_6345;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_5782;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_649;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_6050;
wire n_625;
wire n_6444;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_6379;
wire n_798;
wire n_2324;
wire n_5563;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_2647;
wire n_883;
wire n_6232;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_6017;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_6362;
wire n_4777;
wire n_5720;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_1285;
wire n_1985;
wire n_6326;
wire n_5898;
wire n_1172;
wire n_6283;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_6213;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_6239;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_5896;
wire n_1649;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_1344;
wire n_6174;
wire n_2730;
wire n_2495;
wire n_6087;
wire n_5249;
wire n_2603;
wire n_2090;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_5969;
wire n_3655;
wire n_3825;
wire n_3225;
wire n_2880;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_6454;
wire n_5022;
wire n_5670;
wire n_1280;
wire n_6041;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_6472;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_5879;
wire n_4403;
wire n_5238;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_3531;
wire n_6375;
wire n_6352;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_6238;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_6081;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_5535;
wire n_645;
wire n_3910;
wire n_3812;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_6002;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_6289;
wire n_3748;
wire n_3272;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_5640;
wire n_2831;
wire n_4318;
wire n_932;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_2123;
wire n_1697;
wire n_6512;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_6108;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_6086;
wire n_1396;
wire n_634;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_5941;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_6340;
wire n_3092;
wire n_1289;
wire n_6219;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1014;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_6067;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_674;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5970;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_3861;
wire n_675;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_6011;
wire n_1886;
wire n_4371;
wire n_6225;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_877;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_6182;
wire n_4041;
wire n_2947;
wire n_6520;
wire n_3918;
wire n_5876;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_697;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_5856;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_2663;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_5596;
wire n_6074;
wire n_2684;
wire n_5983;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_5604;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_673;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_5815;
wire n_4191;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_6306;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_6095;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_5565;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_5520;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_5800;
wire n_5984;
wire n_1838;
wire n_6287;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_5772;
wire n_4775;
wire n_2208;
wire n_5884;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_6308;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_5603;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_6128;
wire n_2489;
wire n_6029;
wire n_1087;
wire n_657;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_5924;
wire n_1505;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_2403;
wire n_1070;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_6005;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_6169;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_5926;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_2589;
wire n_4535;
wire n_755;
wire n_6302;
wire n_2442;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_5919;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_6343;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_6098;
wire n_6014;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2357;
wire n_2025;
wire n_5583;
wire n_4654;
wire n_6433;
wire n_3640;
wire n_642;
wire n_1159;
wire n_3481;
wire n_995;
wire n_2250;
wire n_3033;
wire n_6142;
wire n_5775;
wire n_6462;
wire n_2374;
wire n_1681;
wire n_6034;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_6221;
wire n_6279;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_6071;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_6295;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_6385;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_6143;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_793;
wire n_5967;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_6084;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_5966;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_5735;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_5360;
wire n_6104;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_667;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5877;
wire n_6018;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_1216;
wire n_2716;
wire n_6032;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_6122;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_5454;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_6439;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_5913;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_6406;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_6474;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_4888;
wire n_776;
wire n_1823;
wire n_3350;
wire n_2479;
wire n_6000;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_6425;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_6502;
wire n_6250;
wire n_6288;
wire n_5974;
wire n_6492;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_6046;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_6118;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_5991;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_6251;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_5914;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_6146;
wire n_5813;
wire n_790;
wire n_5833;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_5616;
wire n_5805;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_672;
wire n_6228;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_6102;
wire n_636;
wire n_6274;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_6072;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_6353;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_646;
wire n_1329;
wire n_6322;
wire n_5167;
wire n_5661;
wire n_5830;
wire n_5932;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_6498;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_5558;
wire n_1826;
wire n_5687;
wire n_6378;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5587;
wire n_6304;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_661;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_5651;
wire n_4630;
wire n_1217;
wire n_5645;
wire n_3990;
wire n_1628;
wire n_5766;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_5878;
wire n_5671;
wire n_4534;
wire n_1536;
wire n_6301;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_669;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_6259;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_3774;
wire n_863;
wire n_5733;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_6333;
wire n_5791;
wire n_5727;
wire n_761;
wire n_5946;
wire n_5997;
wire n_2492;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_5657;
wire n_1173;
wire n_4974;
wire n_5975;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_6510;
wire n_3334;
wire n_5938;
wire n_6237;
wire n_5602;
wire n_647;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_3114;
wire n_2741;
wire n_888;
wire n_6360;
wire n_2203;
wire n_2255;
wire n_5246;
wire n_3584;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_6475;
wire n_3982;
wire n_6314;
wire n_6103;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_3796;
wire n_6394;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_5994;
wire n_6495;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_6426;
wire n_2600;
wire n_984;
wire n_5626;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_6350;
wire n_4787;
wire n_5633;
wire n_5664;
wire n_1218;
wire n_5921;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_6159;
wire n_2429;
wire n_985;
wire n_2440;
wire n_6054;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_6235;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_6496;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_6513;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_5925;
wire n_2909;
wire n_754;
wire n_6138;
wire n_5369;
wire n_975;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_6330;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_6477;
wire n_6263;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_6490;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_6184;
wire n_730;
wire n_5817;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_6038;
wire n_5861;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_6313;
wire n_784;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_3965;
wire n_5859;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_5776;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_2091;
wire n_5920;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_6180;
wire n_5683;
wire n_6349;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_6476;
wire n_1742;
wire n_4030;

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_505),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_601),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_426),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_88),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_454),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_22),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_527),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_111),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_244),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_378),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_153),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_470),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_262),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_523),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_267),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_179),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_440),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_555),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_299),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_184),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_444),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_284),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_491),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_478),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_177),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_575),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_623),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_252),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_69),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_501),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_371),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_478),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_579),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_312),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_531),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_520),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_502),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_419),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_587),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_284),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_302),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_464),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_209),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_63),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_350),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_49),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_133),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_209),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_613),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_572),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_78),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_414),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_312),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_331),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_512),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_551),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_599),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_117),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_507),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_418),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_567),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_568),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_370),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_18),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_448),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_494),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_432),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_354),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_169),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_453),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_419),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_619),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_287),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_477),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_483),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_425),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_598),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_134),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_508),
.Y(n_703)
);

CKINVDCx14_ASAP7_75t_R g704 ( 
.A(n_504),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_511),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_32),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_255),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_580),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_112),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_109),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_79),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_525),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_433),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_363),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_358),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_481),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_621),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_12),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_320),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_532),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_138),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_502),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_31),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_56),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_368),
.B(n_249),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_477),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_204),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_463),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_524),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_500),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_169),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_190),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_413),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_473),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_83),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_155),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_606),
.Y(n_738)
);

CKINVDCx16_ASAP7_75t_R g739 ( 
.A(n_602),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_604),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_592),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_608),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_190),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_16),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_383),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_232),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_594),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_268),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_221),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_569),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_129),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_298),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_466),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_196),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_584),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_441),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_580),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_220),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_273),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_549),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_517),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_556),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_144),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_536),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_513),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_75),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_245),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_95),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_357),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_576),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_100),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_107),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_238),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_620),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_447),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_271),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_588),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_133),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_59),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_545),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_330),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_213),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_382),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_385),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_96),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_313),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_303),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_433),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_557),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_516),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_174),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_8),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_341),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_448),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_106),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_498),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_378),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_294),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_309),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_392),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_160),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_576),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_154),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_566),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_476),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_357),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_213),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_613),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_554),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_401),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_236),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_586),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_30),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_260),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_407),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_65),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_180),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_323),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_475),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_568),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_541),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_560),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_217),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_440),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_313),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_615),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_281),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_386),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_425),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_111),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_44),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_462),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_410),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_242),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_512),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_495),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_376),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_180),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_622),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_590),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_593),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_29),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_510),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_435),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_561),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_305),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_562),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_522),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_73),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_311),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_581),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_3),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_390),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_205),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_204),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_143),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_230),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_601),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_184),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_207),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_403),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_94),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_224),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_578),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_559),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_517),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_212),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_97),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_90),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_147),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_366),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_465),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_368),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_201),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_497),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_577),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_197),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_612),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_551),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_452),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_329),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_212),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_338),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_113),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_25),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_582),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_595),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_163),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_439),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_109),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_330),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_15),
.Y(n_892)
);

BUFx10_ASAP7_75t_L g893 ( 
.A(n_417),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_103),
.Y(n_894)
);

BUFx10_ASAP7_75t_L g895 ( 
.A(n_110),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_254),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_318),
.Y(n_897)
);

CKINVDCx16_ASAP7_75t_R g898 ( 
.A(n_119),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_615),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_362),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_567),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_285),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_179),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_333),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_320),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_293),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_427),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_423),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_272),
.Y(n_909)
);

CKINVDCx14_ASAP7_75t_R g910 ( 
.A(n_65),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_581),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_150),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_290),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_455),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_452),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_584),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_480),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_340),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_123),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_229),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_202),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_345),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_409),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_504),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_118),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_356),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_186),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_610),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_607),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_561),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_66),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_206),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_265),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_565),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_88),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_251),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_1),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_605),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_458),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_273),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_353),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_614),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_304),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_408),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_574),
.Y(n_945)
);

INVxp33_ASAP7_75t_R g946 ( 
.A(n_294),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_96),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_67),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_423),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_139),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_76),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_393),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_81),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_269),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_85),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_537),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_236),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_247),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_304),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_143),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_47),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_621),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_401),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_316),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_26),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_223),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_445),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_611),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_506),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_323),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_249),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_418),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_545),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_600),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_33),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_437),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_585),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_397),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_528),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_56),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_410),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_306),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_121),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_492),
.Y(n_984)
);

BUFx8_ASAP7_75t_SL g985 ( 
.A(n_549),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_591),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_324),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_287),
.Y(n_988)
);

CKINVDCx16_ASAP7_75t_R g989 ( 
.A(n_291),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_407),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_583),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_540),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_168),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_1),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_571),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_511),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_104),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_442),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_319),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_10),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_26),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_274),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_579),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_339),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_539),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_530),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_68),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_219),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_91),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_519),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_107),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_620),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_0),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_181),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_18),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_609),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_285),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_76),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_334),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_22),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_128),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_358),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_550),
.Y(n_1023)
);

BUFx5_ASAP7_75t_L g1024 ( 
.A(n_591),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_289),
.Y(n_1025)
);

CKINVDCx16_ASAP7_75t_R g1026 ( 
.A(n_611),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_322),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_333),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_29),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_3),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_165),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_388),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_344),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_31),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_71),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_392),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_496),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_117),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_299),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_603),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_271),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_522),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_274),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_150),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_394),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_37),
.Y(n_1046)
);

CKINVDCx16_ASAP7_75t_R g1047 ( 
.A(n_71),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_443),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_489),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_519),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_569),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_524),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_426),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_94),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_521),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_503),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_495),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_4),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_347),
.Y(n_1059)
);

BUFx10_ASAP7_75t_L g1060 ( 
.A(n_520),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_91),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_160),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_505),
.Y(n_1063)
);

CKINVDCx16_ASAP7_75t_R g1064 ( 
.A(n_39),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_50),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_493),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_441),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_242),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_388),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_360),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_112),
.Y(n_1071)
);

BUFx10_ASAP7_75t_L g1072 ( 
.A(n_366),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_231),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_344),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_553),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_489),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_571),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_514),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_455),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_37),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_206),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_575),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_529),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_421),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_526),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_589),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_985),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1024),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1024),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_985),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_704),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_704),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_688),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_910),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_625),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1024),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1024),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1024),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1024),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_688),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_910),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_671),
.B(n_1),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1024),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1024),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_629),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1024),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_706),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_625),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1024),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_636),
.Y(n_1110)
);

BUFx5_ASAP7_75t_L g1111 ( 
.A(n_636),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_632),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_650),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_632),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_650),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_639),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_635),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_671),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_635),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_739),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_739),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_639),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_650),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_694),
.Y(n_1124)
);

CKINVDCx16_ASAP7_75t_R g1125 ( 
.A(n_898),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_650),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_624),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_898),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_624),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_644),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_644),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_644),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_748),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_748),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_989),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_989),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_650),
.Y(n_1137)
);

BUFx5_ASAP7_75t_L g1138 ( 
.A(n_748),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_766),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_650),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_766),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1026),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1026),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1047),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_726),
.B(n_0),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_682),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1047),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_766),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1080),
.Y(n_1149)
);

INVxp33_ASAP7_75t_SL g1150 ( 
.A(n_743),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_782),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1064),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1080),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_743),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_682),
.Y(n_1155)
);

BUFx2_ASAP7_75t_R g1156 ( 
.A(n_1025),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1064),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_626),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_782),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_694),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_782),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_627),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_784),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_784),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_784),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_628),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_630),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_650),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_634),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_638),
.Y(n_1170)
);

INVxp33_ASAP7_75t_SL g1171 ( 
.A(n_808),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_857),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_640),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1080),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_857),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1080),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_713),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_857),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_876),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_641),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_642),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_876),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_876),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_643),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_925),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_645),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_648),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_925),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_925),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_808),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_927),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_649),
.Y(n_1192)
);

CKINVDCx6p67_ASAP7_75t_R g1193 ( 
.A(n_674),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_927),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_724),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_813),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_927),
.Y(n_1197)
);

CKINVDCx16_ASAP7_75t_R g1198 ( 
.A(n_674),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_713),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_955),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_955),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_790),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_955),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_852),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_892),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_965),
.Y(n_1206)
);

CKINVDCx16_ASAP7_75t_R g1207 ( 
.A(n_674),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_747),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_975),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_957),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_994),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_957),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_957),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1015),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1010),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1020),
.Y(n_1216)
);

NOR2xp67_ASAP7_75t_L g1217 ( 
.A(n_726),
.B(n_0),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1010),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_L g1219 ( 
.A(n_956),
.B(n_2),
.Y(n_1219)
);

INVxp33_ASAP7_75t_L g1220 ( 
.A(n_956),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_691),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1058),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1010),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1017),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1017),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_651),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_652),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_747),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_790),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_655),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1017),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_719),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_656),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_719),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_657),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_691),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_744),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_659),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_744),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_660),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_691),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_662),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_664),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_666),
.Y(n_1244)
);

CKINVDCx14_ASAP7_75t_R g1245 ( 
.A(n_674),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_792),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_792),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_842),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_691),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_842),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_753),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_668),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_669),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_885),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_676),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_885),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_937),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_937),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1000),
.Y(n_1259)
);

XNOR2xp5_ASAP7_75t_L g1260 ( 
.A(n_753),
.B(n_2),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1000),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1013),
.Y(n_1262)
);

BUFx8_ASAP7_75t_SL g1263 ( 
.A(n_816),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1013),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1030),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1030),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_670),
.Y(n_1267)
);

BUFx5_ASAP7_75t_L g1268 ( 
.A(n_631),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1034),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_691),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1034),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_672),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_677),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_679),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_691),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_691),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1001),
.B(n_3),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_685),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_745),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_687),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_745),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_745),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_745),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_745),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_745),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_692),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_745),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_850),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_850),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_693),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_695),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_850),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_696),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_850),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_850),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_850),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_850),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_864),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_864),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_816),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_864),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_697),
.Y(n_1302)
);

CKINVDCx14_ASAP7_75t_R g1303 ( 
.A(n_676),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_864),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_864),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_864),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_864),
.Y(n_1307)
);

CKINVDCx16_ASAP7_75t_R g1308 ( 
.A(n_676),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_879),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_879),
.Y(n_1310)
);

BUFx5_ASAP7_75t_L g1311 ( 
.A(n_631),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_879),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_698),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_879),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_879),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_700),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_879),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_919),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_919),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_919),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_701),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_702),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_919),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_834),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_919),
.Y(n_1325)
);

BUFx5_ASAP7_75t_L g1326 ( 
.A(n_646),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_821),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_919),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1054),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1054),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_703),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_705),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_707),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1054),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_L g1335 ( 
.A(n_740),
.B(n_2),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1054),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1054),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1054),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1056),
.Y(n_1339)
);

BUFx10_ASAP7_75t_L g1340 ( 
.A(n_1056),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_708),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_710),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1056),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1056),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_821),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1056),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1056),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1069),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_711),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_716),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1069),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_717),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_720),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1069),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1069),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1069),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_721),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1069),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_722),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_723),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_731),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_732),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1080),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_676),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1080),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1080),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_735),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_646),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_654),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_736),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_654),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_740),
.B(n_4),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_658),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_738),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_741),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_658),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_661),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_742),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_661),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_831),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_804),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_633),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_746),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_665),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_665),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_730),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_730),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_633),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_667),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_749),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_831),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_730),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_667),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_673),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_750),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_751),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_678),
.B(n_5),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_754),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_924),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_633),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_730),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_673),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_757),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_762),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_869),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_763),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_675),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_675),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_647),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_893),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_765),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_680),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_680),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_647),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_647),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_767),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_653),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_653),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_769),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_771),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_681),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_772),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_681),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_653),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_773),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_684),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_774),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_684),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_776),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_779),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_781),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_783),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_663),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_686),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_686),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_689),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_689),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_893),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_785),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_690),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_893),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_690),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_699),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_834),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_787),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_699),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_869),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_788),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_663),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_791),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_793),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_795),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_796),
.Y(n_1453)
);

INVxp33_ASAP7_75t_SL g1454 ( 
.A(n_797),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_798),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_663),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_709),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_712),
.Y(n_1458)
);

BUFx10_ASAP7_75t_L g1459 ( 
.A(n_678),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_712),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_709),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_893),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_714),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_714),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_709),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_718),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_799),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_801),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_802),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_803),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_805),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_806),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_807),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_886),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_715),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_715),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_718),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_811),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_727),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_886),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_900),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_950),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_812),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_814),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_900),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_815),
.Y(n_1486)
);

BUFx10_ASAP7_75t_L g1487 ( 
.A(n_678),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_715),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_817),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_727),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_752),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_728),
.Y(n_1492)
);

BUFx2_ASAP7_75t_SL g1493 ( 
.A(n_895),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_818),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_752),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_822),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_729),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_752),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_729),
.Y(n_1499)
);

CKINVDCx16_ASAP7_75t_R g1500 ( 
.A(n_895),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_733),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_895),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_914),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_823),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1001),
.B(n_6),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_914),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_794),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_824),
.Y(n_1508)
);

NOR2xp67_ASAP7_75t_L g1509 ( 
.A(n_870),
.B(n_5),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_825),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_737),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_983),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_983),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_737),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_829),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_794),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_832),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_836),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_837),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_840),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_755),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_755),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_758),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_758),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_759),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_759),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1021),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_760),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_794),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_841),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_843),
.Y(n_1531)
);

CKINVDCx14_ASAP7_75t_R g1532 ( 
.A(n_895),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_760),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1127),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1461),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1110),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1226),
.Y(n_1537)
);

BUFx2_ASAP7_75t_SL g1538 ( 
.A(n_1087),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1116),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1227),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1230),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1233),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1127),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1235),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1122),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1129),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1129),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1146),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1238),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1240),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1493),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1242),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1108),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1130),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1146),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1131),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1302),
.Y(n_1557)
);

BUFx2_ASAP7_75t_SL g1558 ( 
.A(n_1087),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1324),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1155),
.Y(n_1560)
);

CKINVDCx14_ASAP7_75t_R g1561 ( 
.A(n_1245),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_1444),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1115),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1132),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1133),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1134),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1131),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1139),
.Y(n_1568)
);

INVxp33_ASAP7_75t_SL g1569 ( 
.A(n_1091),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_1155),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1141),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1151),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1243),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1244),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1164),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1159),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1161),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1448),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1163),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1165),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1252),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1172),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1108),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1178),
.Y(n_1584)
);

BUFx2_ASAP7_75t_SL g1585 ( 
.A(n_1364),
.Y(n_1585)
);

INVxp33_ASAP7_75t_L g1586 ( 
.A(n_1263),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1253),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1267),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1179),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1182),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1164),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1272),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1483),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1183),
.Y(n_1594)
);

INVxp67_ASAP7_75t_SL g1595 ( 
.A(n_1175),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1095),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1185),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1177),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1188),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1189),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1191),
.Y(n_1601)
);

INVxp33_ASAP7_75t_SL g1602 ( 
.A(n_1092),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_1177),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1199),
.Y(n_1604)
);

INVxp67_ASAP7_75t_SL g1605 ( 
.A(n_1175),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1194),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1197),
.Y(n_1607)
);

CKINVDCx16_ASAP7_75t_R g1608 ( 
.A(n_1125),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1273),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1112),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1200),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1201),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_1199),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1203),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1210),
.Y(n_1615)
);

CKINVDCx16_ASAP7_75t_R g1616 ( 
.A(n_1303),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1212),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1215),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1213),
.Y(n_1619)
);

INVxp33_ASAP7_75t_SL g1620 ( 
.A(n_1094),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1218),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1223),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1224),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1225),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1341),
.Y(n_1625)
);

CKINVDCx20_ASAP7_75t_R g1626 ( 
.A(n_1208),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1231),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1208),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1213),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1342),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1275),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1115),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1228),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1276),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1228),
.Y(n_1635)
);

INVxp33_ASAP7_75t_SL g1636 ( 
.A(n_1101),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1349),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1114),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1386),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1114),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1386),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1279),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1350),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1281),
.Y(n_1644)
);

CKINVDCx20_ASAP7_75t_R g1645 ( 
.A(n_1251),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1282),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1352),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1353),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1283),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1357),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1111),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1111),
.Y(n_1652)
);

CKINVDCx16_ASAP7_75t_R g1653 ( 
.A(n_1532),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1359),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1360),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1251),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1361),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1285),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1287),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1362),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1292),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1294),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1300),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1140),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1295),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1296),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1300),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1367),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1297),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1327),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1298),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1299),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1301),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1370),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1305),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1306),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1309),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1374),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1312),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1315),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_1327),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1317),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1319),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1117),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1323),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1328),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1375),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1345),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1329),
.Y(n_1689)
);

INVxp33_ASAP7_75t_SL g1690 ( 
.A(n_1090),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1330),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1334),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1336),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1337),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1343),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1378),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1345),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1380),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1344),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1347),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1348),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1356),
.Y(n_1702)
);

INVxp67_ASAP7_75t_SL g1703 ( 
.A(n_1392),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1392),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1358),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1365),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1459),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1304),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1304),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1123),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_1380),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1339),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1339),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1363),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1117),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1363),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1088),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1089),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1383),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1096),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1097),
.Y(n_1721)
);

CKINVDCx20_ASAP7_75t_R g1722 ( 
.A(n_1391),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1119),
.Y(n_1723)
);

INVxp33_ASAP7_75t_SL g1724 ( 
.A(n_1090),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1429),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_1391),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1390),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1098),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1401),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1119),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1395),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1099),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1103),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1396),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1111),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1104),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1401),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1106),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1398),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1120),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1123),
.Y(n_1741)
);

INVxp33_ASAP7_75t_L g1742 ( 
.A(n_1263),
.Y(n_1742)
);

CKINVDCx16_ASAP7_75t_R g1743 ( 
.A(n_1198),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1382),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1403),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1382),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1120),
.Y(n_1747)
);

INVxp33_ASAP7_75t_SL g1748 ( 
.A(n_1121),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1382),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1404),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1382),
.Y(n_1751)
);

INVxp33_ASAP7_75t_SL g1752 ( 
.A(n_1121),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1128),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1111),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1128),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1406),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1381),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1399),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1405),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1409),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1405),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1472),
.Y(n_1762)
);

INVxp33_ASAP7_75t_L g1763 ( 
.A(n_1154),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1409),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1447),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1126),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1409),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1411),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1409),
.Y(n_1769)
);

CKINVDCx14_ASAP7_75t_R g1770 ( 
.A(n_1193),
.Y(n_1770)
);

CKINVDCx16_ASAP7_75t_R g1771 ( 
.A(n_1207),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1484),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1415),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1415),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1416),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1447),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1419),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1415),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1420),
.Y(n_1779)
);

INVxp33_ASAP7_75t_SL g1780 ( 
.A(n_1135),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1415),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1449),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1474),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1449),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1449),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1422),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1457),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1474),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1425),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1457),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1135),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1457),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1427),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1515),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1457),
.Y(n_1795)
);

INVxp33_ASAP7_75t_SL g1796 ( 
.A(n_1136),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1465),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1465),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1465),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1465),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1475),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1475),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1517),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1480),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1518),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1475),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1475),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1519),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1476),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1476),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1476),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1520),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_1480),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1476),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1126),
.Y(n_1815)
);

CKINVDCx16_ASAP7_75t_R g1816 ( 
.A(n_1255),
.Y(n_1816)
);

INVxp67_ASAP7_75t_SL g1817 ( 
.A(n_1441),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1105),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1441),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1137),
.Y(n_1820)
);

INVxp33_ASAP7_75t_SL g1821 ( 
.A(n_1136),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1107),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1495),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1495),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1137),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1495),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1149),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1495),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1142),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1498),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_1481),
.Y(n_1831)
);

CKINVDCx16_ASAP7_75t_R g1832 ( 
.A(n_1308),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1498),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1498),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1462),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1498),
.Y(n_1836)
);

INVxp33_ASAP7_75t_L g1837 ( 
.A(n_1220),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1232),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1234),
.Y(n_1839)
);

CKINVDCx16_ASAP7_75t_R g1840 ( 
.A(n_1500),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1237),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_1481),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1239),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1246),
.Y(n_1844)
);

INVxp33_ASAP7_75t_SL g1845 ( 
.A(n_1142),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1195),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1247),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1248),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1196),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1204),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1140),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1250),
.Y(n_1852)
);

INVxp33_ASAP7_75t_L g1853 ( 
.A(n_1118),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1254),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1257),
.Y(n_1855)
);

CKINVDCx20_ASAP7_75t_R g1856 ( 
.A(n_1485),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1258),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1259),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1261),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1262),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1264),
.Y(n_1861)
);

CKINVDCx14_ASAP7_75t_R g1862 ( 
.A(n_1193),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1205),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1265),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1206),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1266),
.Y(n_1866)
);

INVxp67_ASAP7_75t_SL g1867 ( 
.A(n_1462),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1269),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1143),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1364),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1271),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1111),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1209),
.Y(n_1873)
);

CKINVDCx20_ASAP7_75t_R g1874 ( 
.A(n_1485),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1503),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1111),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1503),
.Y(n_1877)
);

CKINVDCx16_ASAP7_75t_R g1878 ( 
.A(n_1482),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1149),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1111),
.Y(n_1880)
);

INVxp67_ASAP7_75t_L g1881 ( 
.A(n_1387),
.Y(n_1881)
);

CKINVDCx16_ASAP7_75t_R g1882 ( 
.A(n_1506),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1138),
.Y(n_1883)
);

CKINVDCx20_ASAP7_75t_R g1884 ( 
.A(n_1506),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1211),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1138),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1138),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1138),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1138),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1138),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1214),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1138),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1368),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1369),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1216),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1371),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1373),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1387),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1148),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1222),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1148),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1158),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1153),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1512),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1143),
.Y(n_1905)
);

INVxp67_ASAP7_75t_SL g1906 ( 
.A(n_1113),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1899),
.B(n_1388),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1563),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1708),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1585),
.A2(n_1021),
.B1(n_1040),
.B2(n_1027),
.Y(n_1910)
);

BUFx12f_ASAP7_75t_L g1911 ( 
.A(n_1818),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1901),
.B(n_1113),
.Y(n_1912)
);

AND2x6_ASAP7_75t_L g1913 ( 
.A(n_1651),
.B(n_800),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1536),
.Y(n_1914)
);

NOR2x1_ASAP7_75t_L g1915 ( 
.A(n_1899),
.B(n_1145),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1664),
.Y(n_1916)
);

OA21x2_ASAP7_75t_L g1917 ( 
.A1(n_1631),
.A2(n_1168),
.B(n_1153),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1709),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1878),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1563),
.Y(n_1920)
);

CKINVDCx11_ASAP7_75t_R g1921 ( 
.A(n_1534),
.Y(n_1921)
);

AND2x6_ASAP7_75t_L g1922 ( 
.A(n_1651),
.B(n_800),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1632),
.Y(n_1923)
);

AND2x2_ASAP7_75t_SL g1924 ( 
.A(n_1583),
.B(n_1102),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1539),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1664),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1632),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1664),
.Y(n_1928)
);

AND2x6_ASAP7_75t_L g1929 ( 
.A(n_1652),
.B(n_800),
.Y(n_1929)
);

OA21x2_ASAP7_75t_L g1930 ( 
.A1(n_1634),
.A2(n_1174),
.B(n_1168),
.Y(n_1930)
);

OAI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1872),
.A2(n_1109),
.B(n_1174),
.Y(n_1931)
);

OA21x2_ASAP7_75t_L g1932 ( 
.A1(n_1642),
.A2(n_1241),
.B(n_1176),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1712),
.Y(n_1933)
);

CKINVDCx11_ASAP7_75t_R g1934 ( 
.A(n_1534),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1906),
.B(n_1113),
.Y(n_1935)
);

BUFx8_ASAP7_75t_L g1936 ( 
.A(n_1610),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1710),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1851),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1870),
.B(n_1454),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1713),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1851),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1851),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1559),
.A2(n_1217),
.B1(n_1171),
.B2(n_1150),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1567),
.B(n_1388),
.Y(n_1944)
);

AO22x1_ASAP7_75t_L g1945 ( 
.A1(n_1562),
.A2(n_1397),
.B1(n_1171),
.B2(n_1150),
.Y(n_1945)
);

NOR2x1_ASAP7_75t_L g1946 ( 
.A(n_1556),
.B(n_1219),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1710),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1652),
.Y(n_1948)
);

OAI21x1_ASAP7_75t_L g1949 ( 
.A1(n_1876),
.A2(n_1109),
.B(n_1176),
.Y(n_1949)
);

INVx4_ASAP7_75t_L g1950 ( 
.A(n_1735),
.Y(n_1950)
);

OA21x2_ASAP7_75t_L g1951 ( 
.A1(n_1644),
.A2(n_1249),
.B(n_1241),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1629),
.B(n_1545),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1741),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1575),
.B(n_1249),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1595),
.B(n_1284),
.Y(n_1955)
);

BUFx8_ASAP7_75t_L g1956 ( 
.A(n_1638),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1735),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1714),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1716),
.Y(n_1959)
);

OA21x2_ASAP7_75t_L g1960 ( 
.A1(n_1646),
.A2(n_1658),
.B(n_1649),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1717),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1561),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1718),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1554),
.B(n_1400),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1741),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1720),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1754),
.Y(n_1967)
);

INVx5_ASAP7_75t_L g1968 ( 
.A(n_1754),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1556),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1605),
.B(n_1400),
.Y(n_1970)
);

BUFx12f_ASAP7_75t_L g1971 ( 
.A(n_1818),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1619),
.B(n_1414),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1766),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1564),
.Y(n_1974)
);

NAND2xp33_ASAP7_75t_L g1975 ( 
.A(n_1721),
.B(n_1268),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1766),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1815),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1815),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1557),
.A2(n_1454),
.B1(n_1144),
.B2(n_1152),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1820),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1565),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1820),
.Y(n_1982)
);

OAI21x1_ASAP7_75t_L g1983 ( 
.A1(n_1880),
.A2(n_1310),
.B(n_1284),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1825),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1566),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1616),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1881),
.B(n_1158),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1825),
.Y(n_1988)
);

OA21x2_ASAP7_75t_L g1989 ( 
.A1(n_1659),
.A2(n_1314),
.B(n_1310),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1728),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1591),
.B(n_1414),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1568),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1591),
.B(n_1417),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1707),
.B(n_1162),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1571),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1572),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1827),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1827),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1732),
.Y(n_1999)
);

OA21x2_ASAP7_75t_L g2000 ( 
.A1(n_1661),
.A2(n_1320),
.B(n_1314),
.Y(n_2000)
);

INVx5_ASAP7_75t_L g2001 ( 
.A(n_1879),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1733),
.B(n_1320),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1736),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1879),
.Y(n_2004)
);

OAI22x1_ASAP7_75t_L g2005 ( 
.A1(n_1757),
.A2(n_1260),
.B1(n_1124),
.B2(n_1229),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1576),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1903),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1577),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1744),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1579),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1580),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1662),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1665),
.Y(n_2013)
);

OA21x2_ASAP7_75t_L g2014 ( 
.A1(n_1666),
.A2(n_1351),
.B(n_1346),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1582),
.B(n_1584),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1738),
.Y(n_2016)
);

OA21x2_ASAP7_75t_L g2017 ( 
.A1(n_1669),
.A2(n_1351),
.B(n_1346),
.Y(n_2017)
);

OAI21x1_ASAP7_75t_L g2018 ( 
.A1(n_1883),
.A2(n_1366),
.B(n_1529),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1758),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1671),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1886),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1535),
.B(n_1366),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1672),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1898),
.B(n_1162),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1673),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1653),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1675),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1589),
.B(n_1417),
.Y(n_2028)
);

OAI22x1_ASAP7_75t_SL g2029 ( 
.A1(n_1543),
.A2(n_1100),
.B1(n_1093),
.B2(n_1512),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_1543),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1746),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1749),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1751),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1590),
.B(n_1424),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1760),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1594),
.B(n_1424),
.Y(n_2036)
);

OAI21x1_ASAP7_75t_L g2037 ( 
.A1(n_1887),
.A2(n_1529),
.B(n_1456),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1764),
.B(n_1166),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1767),
.Y(n_2039)
);

BUFx8_ASAP7_75t_SL g2040 ( 
.A(n_1546),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1676),
.Y(n_2041)
);

OA21x2_ASAP7_75t_L g2042 ( 
.A1(n_1677),
.A2(n_1680),
.B(n_1679),
.Y(n_2042)
);

INVx4_ASAP7_75t_L g2043 ( 
.A(n_1888),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1769),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1707),
.B(n_1551),
.Y(n_2045)
);

CKINVDCx20_ASAP7_75t_R g2046 ( 
.A(n_1546),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1773),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1682),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1578),
.B(n_1166),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1683),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_1593),
.A2(n_1147),
.B1(n_1152),
.B2(n_1144),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1597),
.B(n_1433),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1889),
.A2(n_1892),
.B(n_1890),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1685),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1686),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1689),
.Y(n_2056)
);

INVx5_ASAP7_75t_L g2057 ( 
.A(n_1596),
.Y(n_2057)
);

OAI21x1_ASAP7_75t_L g2058 ( 
.A1(n_1691),
.A2(n_1516),
.B(n_1456),
.Y(n_2058)
);

CKINVDCx16_ASAP7_75t_R g2059 ( 
.A(n_1608),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1692),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1837),
.B(n_1725),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1693),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1694),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1774),
.Y(n_2064)
);

INVx4_ASAP7_75t_L g2065 ( 
.A(n_1778),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_1755),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1781),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1782),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_1762),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1695),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1699),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1599),
.B(n_1433),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1770),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1772),
.A2(n_1157),
.B1(n_1169),
.B2(n_1167),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1600),
.Y(n_2075)
);

BUFx2_ASAP7_75t_L g2076 ( 
.A(n_1869),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1601),
.Y(n_2077)
);

BUFx12f_ASAP7_75t_L g2078 ( 
.A(n_1822),
.Y(n_2078)
);

INVxp33_ASAP7_75t_L g2079 ( 
.A(n_1853),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1606),
.Y(n_2080)
);

CKINVDCx8_ASAP7_75t_R g2081 ( 
.A(n_1538),
.Y(n_2081)
);

OA21x2_ASAP7_75t_L g2082 ( 
.A1(n_1700),
.A2(n_1491),
.B(n_1488),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_1701),
.Y(n_2083)
);

INVxp33_ASAP7_75t_SL g2084 ( 
.A(n_1822),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1862),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1607),
.Y(n_2086)
);

CKINVDCx6p67_ASAP7_75t_R g2087 ( 
.A(n_1743),
.Y(n_2087)
);

BUFx8_ASAP7_75t_SL g2088 ( 
.A(n_1547),
.Y(n_2088)
);

BUFx8_ASAP7_75t_SL g2089 ( 
.A(n_1547),
.Y(n_2089)
);

BUFx6f_ASAP7_75t_L g2090 ( 
.A(n_1784),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1639),
.A2(n_1641),
.B1(n_1704),
.B2(n_1703),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1702),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1705),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1611),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1612),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1614),
.Y(n_2096)
);

BUFx8_ASAP7_75t_L g2097 ( 
.A(n_1838),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_1729),
.A2(n_1160),
.B1(n_1170),
.B2(n_1169),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1785),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1787),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1615),
.B(n_1488),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1617),
.Y(n_2102)
);

OA21x2_ASAP7_75t_L g2103 ( 
.A1(n_1706),
.A2(n_1792),
.B(n_1790),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1795),
.B(n_1170),
.Y(n_2104)
);

INVxp33_ASAP7_75t_SL g2105 ( 
.A(n_1873),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_1553),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1797),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1618),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1798),
.B(n_1173),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1621),
.Y(n_2110)
);

AOI22x1_ASAP7_75t_SL g2111 ( 
.A1(n_1548),
.A2(n_1100),
.B1(n_1093),
.B2(n_1027),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1622),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1799),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1800),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1801),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1623),
.B(n_1491),
.Y(n_2116)
);

AND2x6_ASAP7_75t_L g2117 ( 
.A(n_1624),
.B(n_839),
.Y(n_2117)
);

OAI21x1_ASAP7_75t_L g2118 ( 
.A1(n_1802),
.A2(n_1516),
.B(n_1507),
.Y(n_2118)
);

CKINVDCx20_ASAP7_75t_R g2119 ( 
.A(n_1548),
.Y(n_2119)
);

OA21x2_ASAP7_75t_L g2120 ( 
.A1(n_1806),
.A2(n_1507),
.B(n_1377),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1807),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_L g2122 ( 
.A1(n_1809),
.A2(n_1418),
.B(n_872),
.Y(n_2122)
);

OAI21x1_ASAP7_75t_L g2123 ( 
.A1(n_1810),
.A2(n_1418),
.B(n_872),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1811),
.Y(n_2124)
);

CKINVDCx6p67_ASAP7_75t_R g2125 ( 
.A(n_1771),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1627),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1839),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1814),
.B(n_1173),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1823),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1841),
.Y(n_2130)
);

CKINVDCx8_ASAP7_75t_R g2131 ( 
.A(n_1558),
.Y(n_2131)
);

OAI22x1_ASAP7_75t_SL g2132 ( 
.A1(n_1555),
.A2(n_1527),
.B1(n_1513),
.B2(n_1040),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1824),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1826),
.Y(n_2134)
);

INVx6_ASAP7_75t_L g2135 ( 
.A(n_1816),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_1843),
.B(n_1376),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1828),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1830),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_1737),
.A2(n_1181),
.B1(n_1184),
.B2(n_1180),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1833),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1552),
.B(n_1180),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1834),
.B(n_1181),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1836),
.B(n_1184),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1844),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1893),
.Y(n_2145)
);

BUFx8_ASAP7_75t_SL g2146 ( 
.A(n_1555),
.Y(n_2146)
);

INVx5_ASAP7_75t_L g2147 ( 
.A(n_1817),
.Y(n_2147)
);

CKINVDCx20_ASAP7_75t_R g2148 ( 
.A(n_1560),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1873),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1894),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1847),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1896),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1848),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1852),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1854),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1855),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1897),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1857),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1819),
.B(n_1186),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1858),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1859),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_1860),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_1835),
.A2(n_1867),
.B1(n_1752),
.B2(n_1780),
.Y(n_2163)
);

OA21x2_ASAP7_75t_L g2164 ( 
.A1(n_1861),
.A2(n_1384),
.B(n_1379),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_1864),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_1866),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1868),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1871),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1625),
.B(n_1186),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1630),
.Y(n_2170)
);

AOI22x1_ASAP7_75t_SL g2171 ( 
.A1(n_1570),
.A2(n_1051),
.B1(n_1068),
.B2(n_1059),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1637),
.B(n_1187),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1643),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1647),
.B(n_1187),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_1846),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1849),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1640),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1850),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1648),
.B(n_1192),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_1684),
.B(n_1385),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1650),
.B(n_1192),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_1668),
.B(n_1274),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1715),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1674),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1678),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1723),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1730),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1895),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1687),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_L g2190 ( 
.A1(n_1740),
.A2(n_1418),
.B(n_872),
.Y(n_2190)
);

BUFx6f_ASAP7_75t_L g2191 ( 
.A(n_1863),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1747),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_1696),
.B(n_1274),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1763),
.B(n_1459),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1719),
.B(n_1459),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1753),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1791),
.Y(n_2197)
);

OAI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_1569),
.A2(n_1280),
.B1(n_1286),
.B2(n_1278),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1829),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1905),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1865),
.Y(n_2201)
);

INVxp67_ASAP7_75t_L g2202 ( 
.A(n_1902),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1885),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_1882),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1727),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1731),
.Y(n_2206)
);

OAI22xp33_ASAP7_75t_SL g2207 ( 
.A1(n_1569),
.A2(n_1190),
.B1(n_1505),
.B2(n_1277),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_1734),
.B(n_1389),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1739),
.Y(n_2209)
);

INVx4_ASAP7_75t_L g2210 ( 
.A(n_1745),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_1895),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_1900),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1750),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1891),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_1537),
.Y(n_2215)
);

OA21x2_ASAP7_75t_L g2216 ( 
.A1(n_1537),
.A2(n_1394),
.B(n_1393),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_1540),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_1602),
.A2(n_1286),
.B1(n_1290),
.B2(n_1280),
.Y(n_2218)
);

OAI22x1_ASAP7_75t_L g2219 ( 
.A1(n_1900),
.A2(n_1202),
.B1(n_1438),
.B2(n_1410),
.Y(n_2219)
);

AND2x6_ASAP7_75t_L g2220 ( 
.A(n_1602),
.B(n_839),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_1620),
.A2(n_1291),
.B1(n_1293),
.B2(n_1290),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1540),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_1541),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_1620),
.A2(n_1293),
.B1(n_1313),
.B2(n_1291),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1541),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1542),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_1542),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1544),
.B(n_1313),
.Y(n_2228)
);

INVxp33_ASAP7_75t_SL g2229 ( 
.A(n_1544),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1549),
.Y(n_2230)
);

OA21x2_ASAP7_75t_L g2231 ( 
.A1(n_1549),
.A2(n_1407),
.B(n_1402),
.Y(n_2231)
);

OA21x2_ASAP7_75t_L g2232 ( 
.A1(n_1550),
.A2(n_1412),
.B(n_1408),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1550),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1573),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1573),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_1748),
.A2(n_1321),
.B1(n_1322),
.B2(n_1316),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1574),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1574),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1581),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_1581),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1587),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1587),
.B(n_1316),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1588),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1588),
.B(n_1413),
.Y(n_2244)
);

INVxp67_ASAP7_75t_L g2245 ( 
.A(n_1592),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1592),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1609),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1609),
.Y(n_2248)
);

INVx5_ASAP7_75t_L g2249 ( 
.A(n_1832),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_1654),
.Y(n_2250)
);

BUFx6f_ASAP7_75t_L g2251 ( 
.A(n_1654),
.Y(n_2251)
);

AND2x6_ASAP7_75t_L g2252 ( 
.A(n_1636),
.B(n_839),
.Y(n_2252)
);

BUFx2_ASAP7_75t_L g2253 ( 
.A(n_1655),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1655),
.B(n_1487),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1657),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_1657),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1660),
.Y(n_2257)
);

OA21x2_ASAP7_75t_L g2258 ( 
.A1(n_1660),
.A2(n_1423),
.B(n_1421),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1756),
.Y(n_2259)
);

INVx4_ASAP7_75t_L g2260 ( 
.A(n_1756),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1768),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_1768),
.Y(n_2262)
);

OAI22x1_ASAP7_75t_SL g2263 ( 
.A1(n_1570),
.A2(n_1527),
.B1(n_1513),
.B2(n_1051),
.Y(n_2263)
);

BUFx8_ASAP7_75t_L g2264 ( 
.A(n_1840),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1775),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1777),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1777),
.B(n_1487),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1779),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1779),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_1636),
.B(n_1321),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1786),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_1748),
.A2(n_1331),
.B1(n_1332),
.B2(n_1322),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1786),
.B(n_1487),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1789),
.B(n_1410),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1789),
.Y(n_2275)
);

BUFx2_ASAP7_75t_L g2276 ( 
.A(n_1793),
.Y(n_2276)
);

INVx5_ASAP7_75t_L g2277 ( 
.A(n_1793),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1794),
.Y(n_2278)
);

OA21x2_ASAP7_75t_L g2279 ( 
.A1(n_1794),
.A2(n_1428),
.B(n_1426),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1803),
.Y(n_2280)
);

BUFx8_ASAP7_75t_SL g2281 ( 
.A(n_1598),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_1803),
.B(n_1438),
.Y(n_2282)
);

BUFx2_ASAP7_75t_L g2283 ( 
.A(n_1805),
.Y(n_2283)
);

OA21x2_ASAP7_75t_L g2284 ( 
.A1(n_1805),
.A2(n_1435),
.B(n_1434),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1808),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_1808),
.B(n_1502),
.Y(n_2286)
);

HB1xp67_ASAP7_75t_L g2287 ( 
.A(n_1812),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_1812),
.B(n_1331),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_1752),
.A2(n_1333),
.B1(n_1430),
.B2(n_1332),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_1603),
.B(n_1436),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_1780),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_1796),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1603),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1904),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_1604),
.B(n_1437),
.Y(n_2295)
);

BUFx6f_ASAP7_75t_L g2296 ( 
.A(n_1796),
.Y(n_2296)
);

BUFx12f_ASAP7_75t_L g2297 ( 
.A(n_1690),
.Y(n_2297)
);

INVx3_ASAP7_75t_L g2298 ( 
.A(n_1821),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1821),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1845),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_1586),
.B(n_1502),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1845),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_1604),
.B(n_1440),
.Y(n_2303)
);

AOI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_1690),
.A2(n_1430),
.B1(n_1431),
.B2(n_1333),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_1742),
.B(n_1268),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_1724),
.Y(n_2306)
);

BUFx2_ASAP7_75t_L g2307 ( 
.A(n_1613),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_1724),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1904),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1613),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1884),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1884),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1626),
.B(n_1431),
.Y(n_2313)
);

BUFx3_ASAP7_75t_L g2314 ( 
.A(n_1626),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1877),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_1877),
.Y(n_2316)
);

BUFx6f_ASAP7_75t_L g2317 ( 
.A(n_1628),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_1628),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1875),
.Y(n_2319)
);

INVx3_ASAP7_75t_L g2320 ( 
.A(n_1633),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_1633),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_1635),
.B(n_1432),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_1635),
.B(n_1432),
.Y(n_2323)
);

INVx4_ASAP7_75t_L g2324 ( 
.A(n_1645),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_1645),
.B(n_1442),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1656),
.B(n_1439),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1656),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_1663),
.Y(n_2328)
);

BUFx12f_ASAP7_75t_L g2329 ( 
.A(n_1663),
.Y(n_2329)
);

CKINVDCx20_ASAP7_75t_R g2330 ( 
.A(n_1667),
.Y(n_2330)
);

OA21x2_ASAP7_75t_L g2331 ( 
.A1(n_1667),
.A2(n_1446),
.B(n_1443),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_1670),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_1670),
.B(n_1458),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_1681),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_1681),
.B(n_1439),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_1688),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1697),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1991),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1991),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2120),
.Y(n_2340)
);

HB1xp67_ASAP7_75t_L g2341 ( 
.A(n_2019),
.Y(n_2341)
);

CKINVDCx20_ASAP7_75t_R g2342 ( 
.A(n_2030),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_2040),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_2040),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_2120),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_2088),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2082),
.Y(n_2347)
);

BUFx3_ASAP7_75t_L g2348 ( 
.A(n_1969),
.Y(n_2348)
);

BUFx10_ASAP7_75t_L g2349 ( 
.A(n_2288),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1991),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_2149),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2082),
.Y(n_2352)
);

CKINVDCx8_ASAP7_75t_R g2353 ( 
.A(n_2059),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_2149),
.Y(n_2354)
);

CKINVDCx20_ASAP7_75t_R g2355 ( 
.A(n_2030),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1993),
.Y(n_2356)
);

BUFx2_ASAP7_75t_L g2357 ( 
.A(n_2307),
.Y(n_2357)
);

XOR2xp5_ASAP7_75t_L g2358 ( 
.A(n_2204),
.B(n_1697),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1944),
.B(n_1445),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_1969),
.B(n_1460),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_2088),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1993),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_2089),
.Y(n_2363)
);

CKINVDCx20_ASAP7_75t_R g2364 ( 
.A(n_2046),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2194),
.B(n_1445),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_SL g2366 ( 
.A(n_2210),
.B(n_1156),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2079),
.Y(n_2367)
);

CKINVDCx20_ASAP7_75t_R g2368 ( 
.A(n_2046),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_1944),
.B(n_1970),
.Y(n_2369)
);

CKINVDCx20_ASAP7_75t_R g2370 ( 
.A(n_2119),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_1944),
.B(n_1450),
.Y(n_2371)
);

CKINVDCx20_ASAP7_75t_R g2372 ( 
.A(n_2119),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_2146),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_2146),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_1993),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1909),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2281),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_L g2378 ( 
.A(n_2120),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1918),
.Y(n_2379)
);

BUFx6f_ASAP7_75t_L g2380 ( 
.A(n_1948),
.Y(n_2380)
);

NAND2xp33_ASAP7_75t_SL g2381 ( 
.A(n_2219),
.B(n_2274),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2082),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2194),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2144),
.B(n_1463),
.Y(n_2384)
);

HB1xp67_ASAP7_75t_L g2385 ( 
.A(n_2317),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1918),
.Y(n_2386)
);

BUFx2_ASAP7_75t_L g2387 ( 
.A(n_2307),
.Y(n_2387)
);

CKINVDCx20_ASAP7_75t_R g2388 ( 
.A(n_2148),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1933),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_1948),
.Y(n_2390)
);

CKINVDCx5p33_ASAP7_75t_R g2391 ( 
.A(n_2281),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1933),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_1948),
.Y(n_2393)
);

CKINVDCx20_ASAP7_75t_R g2394 ( 
.A(n_2148),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1940),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_2244),
.B(n_1450),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2082),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_1919),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1958),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_1959),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2150),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_1919),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_1921),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_1934),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2150),
.Y(n_2405)
);

NAND2xp33_ASAP7_75t_R g2406 ( 
.A(n_2076),
.B(n_1451),
.Y(n_2406)
);

INVx4_ASAP7_75t_L g2407 ( 
.A(n_1948),
.Y(n_2407)
);

OR2x6_ASAP7_75t_L g2408 ( 
.A(n_2175),
.B(n_725),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_1948),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1970),
.B(n_1451),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2157),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_1970),
.B(n_1452),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2144),
.B(n_1464),
.Y(n_2413)
);

HB1xp67_ASAP7_75t_L g2414 ( 
.A(n_2317),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_1957),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2157),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2151),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_1911),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2037),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_2188),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2037),
.Y(n_2421)
);

AND2x6_ASAP7_75t_L g2422 ( 
.A(n_2305),
.B(n_882),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2151),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2153),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2153),
.Y(n_2425)
);

AND2x6_ASAP7_75t_L g2426 ( 
.A(n_2305),
.B(n_882),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2154),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2155),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2155),
.Y(n_2429)
);

AND2x4_ASAP7_75t_L g2430 ( 
.A(n_1972),
.B(n_1466),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_1972),
.B(n_1952),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2118),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2118),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2156),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2274),
.B(n_1453),
.Y(n_2435)
);

NAND2xp33_ASAP7_75t_L g2436 ( 
.A(n_1913),
.B(n_1268),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2058),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2156),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2058),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_1972),
.B(n_1453),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2158),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2158),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2167),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2167),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_1917),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_2018),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2168),
.Y(n_2447)
);

NAND2xp33_ASAP7_75t_L g2448 ( 
.A(n_1913),
.B(n_1922),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2168),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_2188),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2282),
.B(n_1455),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_2212),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_2212),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_2225),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_2225),
.Y(n_2455)
);

BUFx6f_ASAP7_75t_L g2456 ( 
.A(n_1957),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1964),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_2261),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1964),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_1971),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_1971),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_1917),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2018),
.Y(n_2463)
);

CKINVDCx20_ASAP7_75t_R g2464 ( 
.A(n_2330),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_2078),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_1917),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1917),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_1930),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1961),
.B(n_1467),
.Y(n_2469)
);

CKINVDCx20_ASAP7_75t_R g2470 ( 
.A(n_2330),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_1952),
.B(n_1477),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_1930),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2034),
.Y(n_2473)
);

CKINVDCx20_ASAP7_75t_R g2474 ( 
.A(n_2328),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2034),
.Y(n_2475)
);

INVx3_ASAP7_75t_L g2476 ( 
.A(n_1983),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2052),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2052),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2078),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2072),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_1930),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2061),
.B(n_1467),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_1961),
.B(n_1468),
.Y(n_2483)
);

INVxp67_ASAP7_75t_L g2484 ( 
.A(n_1939),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_1930),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2317),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_1932),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_1932),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2286),
.B(n_2195),
.Y(n_2489)
);

BUFx2_ASAP7_75t_L g2490 ( 
.A(n_2076),
.Y(n_2490)
);

HB1xp67_ASAP7_75t_L g2491 ( 
.A(n_2317),
.Y(n_2491)
);

BUFx3_ASAP7_75t_L g2492 ( 
.A(n_2135),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_2228),
.B(n_1468),
.Y(n_2493)
);

INVx4_ASAP7_75t_L g2494 ( 
.A(n_1957),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2073),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_2242),
.B(n_1469),
.Y(n_2496)
);

BUFx2_ASAP7_75t_L g2497 ( 
.A(n_2314),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2073),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2072),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2116),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2116),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_2085),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2286),
.B(n_1469),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_1957),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2085),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_1932),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2317),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_1963),
.B(n_1470),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_1907),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2015),
.B(n_1907),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2127),
.Y(n_2511)
);

CKINVDCx20_ASAP7_75t_R g2512 ( 
.A(n_2328),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_1957),
.Y(n_2513)
);

OAI22xp5_ASAP7_75t_SL g2514 ( 
.A1(n_1910),
.A2(n_1698),
.B1(n_1722),
.B2(n_1711),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_1932),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_1963),
.B(n_1471),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2130),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_1962),
.Y(n_2518)
);

CKINVDCx20_ASAP7_75t_R g2519 ( 
.A(n_2314),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2254),
.B(n_1473),
.Y(n_2520)
);

BUFx6f_ASAP7_75t_L g2521 ( 
.A(n_1967),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2161),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1914),
.Y(n_2523)
);

CKINVDCx20_ASAP7_75t_R g2524 ( 
.A(n_2316),
.Y(n_2524)
);

CKINVDCx20_ASAP7_75t_R g2525 ( 
.A(n_2316),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_1925),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_1974),
.Y(n_2527)
);

HB1xp67_ASAP7_75t_L g2528 ( 
.A(n_2318),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1981),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_1985),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_1992),
.Y(n_2531)
);

CKINVDCx20_ASAP7_75t_R g2532 ( 
.A(n_2087),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_1962),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1966),
.B(n_1990),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_R g2535 ( 
.A(n_2261),
.B(n_1783),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_1995),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_1986),
.Y(n_2537)
);

CKINVDCx16_ASAP7_75t_R g2538 ( 
.A(n_2329),
.Y(n_2538)
);

CKINVDCx20_ASAP7_75t_R g2539 ( 
.A(n_2087),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_1986),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_2026),
.Y(n_2541)
);

INVxp67_ASAP7_75t_L g2542 ( 
.A(n_1987),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_1951),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_1951),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2015),
.B(n_1490),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_1996),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_1966),
.B(n_1473),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2318),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_2026),
.Y(n_2549)
);

AND2x4_ASAP7_75t_L g2550 ( 
.A(n_2015),
.B(n_1492),
.Y(n_2550)
);

BUFx2_ASAP7_75t_L g2551 ( 
.A(n_2318),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2254),
.B(n_1478),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2006),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2008),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2135),
.Y(n_2555)
);

NOR2xp67_ASAP7_75t_L g2556 ( 
.A(n_2057),
.B(n_2249),
.Y(n_2556)
);

INVx1_ASAP7_75t_SL g2557 ( 
.A(n_2267),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_1989),
.Y(n_2558)
);

INVx4_ASAP7_75t_L g2559 ( 
.A(n_1967),
.Y(n_2559)
);

INVx3_ASAP7_75t_L g2560 ( 
.A(n_1983),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2125),
.Y(n_2561)
);

CKINVDCx20_ASAP7_75t_R g2562 ( 
.A(n_2125),
.Y(n_2562)
);

INVx3_ASAP7_75t_L g2563 ( 
.A(n_1931),
.Y(n_2563)
);

AND2x6_ASAP7_75t_L g2564 ( 
.A(n_1915),
.B(n_882),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2010),
.Y(n_2565)
);

INVx3_ASAP7_75t_L g2566 ( 
.A(n_1931),
.Y(n_2566)
);

INVxp67_ASAP7_75t_L g2567 ( 
.A(n_2024),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_1967),
.Y(n_2568)
);

INVx1_ASAP7_75t_SL g2569 ( 
.A(n_2267),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2011),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_1990),
.B(n_1486),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2003),
.B(n_1486),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2297),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2075),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2077),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2080),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2003),
.B(n_1489),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2329),
.Y(n_2578)
);

INVx4_ASAP7_75t_L g2579 ( 
.A(n_1967),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_1967),
.Y(n_2580)
);

BUFx2_ASAP7_75t_L g2581 ( 
.A(n_2318),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2086),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_1989),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2094),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2264),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_2264),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2000),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2000),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2000),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2095),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2096),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_2084),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2102),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2273),
.B(n_1489),
.Y(n_2594)
);

CKINVDCx20_ASAP7_75t_R g2595 ( 
.A(n_2111),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_1954),
.B(n_1494),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2084),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2108),
.Y(n_2598)
);

BUFx2_ASAP7_75t_L g2599 ( 
.A(n_2318),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_1949),
.Y(n_2600)
);

NAND2x1p5_ASAP7_75t_L g2601 ( 
.A(n_2147),
.B(n_1140),
.Y(n_2601)
);

CKINVDCx20_ASAP7_75t_R g2602 ( 
.A(n_2111),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2110),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_1955),
.B(n_1494),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2273),
.B(n_1496),
.Y(n_2605)
);

CKINVDCx20_ASAP7_75t_R g2606 ( 
.A(n_1936),
.Y(n_2606)
);

OAI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2163),
.A2(n_1504),
.B1(n_1508),
.B2(n_1496),
.Y(n_2607)
);

NOR2xp67_ASAP7_75t_L g2608 ( 
.A(n_2057),
.B(n_1504),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_R g2609 ( 
.A(n_2081),
.B(n_1726),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2014),
.Y(n_2610)
);

OR2x2_ASAP7_75t_L g2611 ( 
.A(n_2293),
.B(n_1508),
.Y(n_2611)
);

CKINVDCx20_ASAP7_75t_R g2612 ( 
.A(n_1936),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2112),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2208),
.B(n_1510),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2014),
.Y(n_2615)
);

BUFx6f_ASAP7_75t_L g2616 ( 
.A(n_1949),
.Y(n_2616)
);

INVxp33_ASAP7_75t_L g2617 ( 
.A(n_2313),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2014),
.Y(n_2618)
);

CKINVDCx20_ASAP7_75t_R g2619 ( 
.A(n_1936),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2126),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2105),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2152),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2152),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2229),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2229),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2152),
.Y(n_2626)
);

XOR2xp5_ASAP7_75t_L g2627 ( 
.A(n_2029),
.B(n_1698),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2162),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2081),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2332),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2162),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2162),
.B(n_1530),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2166),
.Y(n_2633)
);

HB1xp67_ASAP7_75t_L g2634 ( 
.A(n_2332),
.Y(n_2634)
);

NAND2xp33_ASAP7_75t_R g2635 ( 
.A(n_2331),
.B(n_1530),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2166),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_1924),
.B(n_1531),
.Y(n_2637)
);

BUFx2_ASAP7_75t_L g2638 ( 
.A(n_2332),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2131),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2166),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2016),
.B(n_1531),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2016),
.B(n_1268),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_2131),
.Y(n_2643)
);

BUFx6f_ASAP7_75t_L g2644 ( 
.A(n_1999),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2017),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2028),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2028),
.Y(n_2647)
);

CKINVDCx20_ASAP7_75t_R g2648 ( 
.A(n_1956),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2017),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2136),
.B(n_1999),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2215),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2036),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2036),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2215),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_R g2655 ( 
.A(n_2217),
.B(n_1783),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2017),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2017),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_2215),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_2215),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2016),
.B(n_1268),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2215),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_1924),
.B(n_1479),
.Y(n_2662)
);

NAND2xp33_ASAP7_75t_L g2663 ( 
.A(n_1913),
.B(n_1268),
.Y(n_2663)
);

HB1xp67_ASAP7_75t_L g2664 ( 
.A(n_2332),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_2145),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2332),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2036),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2223),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_2103),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2101),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2101),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_2223),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_1923),
.Y(n_2673)
);

CKINVDCx20_ASAP7_75t_R g2674 ( 
.A(n_1956),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2223),
.Y(n_2675)
);

BUFx6f_ASAP7_75t_L g2676 ( 
.A(n_2145),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2277),
.B(n_1335),
.Y(n_2677)
);

BUFx6f_ASAP7_75t_L g2678 ( 
.A(n_2145),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2136),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2023),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_1923),
.Y(n_2681)
);

CKINVDCx20_ASAP7_75t_R g2682 ( 
.A(n_1956),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2023),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2041),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2041),
.Y(n_2685)
);

BUFx6f_ASAP7_75t_L g2686 ( 
.A(n_2145),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_1927),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2223),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2223),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2277),
.B(n_1372),
.Y(n_2690)
);

AND2x4_ASAP7_75t_L g2691 ( 
.A(n_2147),
.B(n_1497),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_1912),
.B(n_1268),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2226),
.Y(n_2693)
);

BUFx6f_ASAP7_75t_L g2694 ( 
.A(n_2145),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2226),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2226),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2226),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_R g2698 ( 
.A(n_2217),
.B(n_1856),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2049),
.B(n_946),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2055),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2055),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2056),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2180),
.B(n_1256),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2056),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2060),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_2226),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2238),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2060),
.Y(n_2708)
);

INVxp67_ASAP7_75t_L g2709 ( 
.A(n_2069),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2063),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_2336),
.Y(n_2711)
);

XNOR2x2_ASAP7_75t_L g2712 ( 
.A(n_2005),
.B(n_946),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2160),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2238),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2063),
.Y(n_2715)
);

CKINVDCx20_ASAP7_75t_R g2716 ( 
.A(n_2336),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_1927),
.Y(n_2717)
);

INVx3_ASAP7_75t_L g2718 ( 
.A(n_2103),
.Y(n_2718)
);

INVx3_ASAP7_75t_L g2719 ( 
.A(n_2103),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2114),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_1937),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_1937),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2114),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_1947),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2137),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_1947),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_1965),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2137),
.Y(n_2728)
);

HB1xp67_ASAP7_75t_L g2729 ( 
.A(n_2336),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_1965),
.Y(n_2730)
);

INVxp33_ASAP7_75t_SL g2731 ( 
.A(n_2211),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2238),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_2238),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2238),
.Y(n_2734)
);

INVx3_ASAP7_75t_L g2735 ( 
.A(n_2103),
.Y(n_2735)
);

INVx3_ASAP7_75t_L g2736 ( 
.A(n_2122),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2180),
.B(n_1509),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2147),
.B(n_1311),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2147),
.B(n_1499),
.Y(n_2739)
);

CKINVDCx20_ASAP7_75t_R g2740 ( 
.A(n_2336),
.Y(n_2740)
);

BUFx6f_ASAP7_75t_L g2741 ( 
.A(n_2160),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_1976),
.Y(n_2742)
);

AND2x2_ASAP7_75t_SL g2743 ( 
.A(n_2216),
.B(n_891),
.Y(n_2743)
);

BUFx6f_ASAP7_75t_L g2744 ( 
.A(n_2160),
.Y(n_2744)
);

INVx3_ASAP7_75t_L g2745 ( 
.A(n_2122),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2240),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_1976),
.Y(n_2747)
);

CKINVDCx20_ASAP7_75t_R g2748 ( 
.A(n_2337),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2138),
.Y(n_2749)
);

BUFx6f_ASAP7_75t_L g2750 ( 
.A(n_2160),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_1935),
.Y(n_2751)
);

CKINVDCx20_ASAP7_75t_R g2752 ( 
.A(n_2337),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2164),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2240),
.Y(n_2754)
);

INVx6_ASAP7_75t_L g2755 ( 
.A(n_2057),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_1978),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2160),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2175),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2164),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_2123),
.Y(n_2760)
);

BUFx2_ASAP7_75t_L g2761 ( 
.A(n_2337),
.Y(n_2761)
);

CKINVDCx20_ASAP7_75t_R g2762 ( 
.A(n_2337),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_1978),
.Y(n_2763)
);

BUFx2_ASAP7_75t_L g2764 ( 
.A(n_2337),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2169),
.B(n_1711),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_1982),
.Y(n_2766)
);

AND2x4_ASAP7_75t_L g2767 ( 
.A(n_2147),
.B(n_1501),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2164),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_1982),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2164),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2240),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2020),
.B(n_1311),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_2240),
.Y(n_2773)
);

CKINVDCx5p33_ASAP7_75t_R g2774 ( 
.A(n_2240),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2012),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2251),
.Y(n_2776)
);

INVx2_ASAP7_75t_SL g2777 ( 
.A(n_2431),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2673),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_2535),
.Y(n_2779)
);

INVx3_ASAP7_75t_L g2780 ( 
.A(n_2600),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2751),
.B(n_2216),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2673),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2681),
.Y(n_2783)
);

INVxp33_ASAP7_75t_L g2784 ( 
.A(n_2341),
.Y(n_2784)
);

NOR2x1p5_ASAP7_75t_L g2785 ( 
.A(n_2492),
.B(n_2291),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_SL g2786 ( 
.A(n_2651),
.B(n_2654),
.Y(n_2786)
);

INVx3_ASAP7_75t_L g2787 ( 
.A(n_2600),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2681),
.Y(n_2788)
);

INVx3_ASAP7_75t_L g2789 ( 
.A(n_2600),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2687),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2687),
.Y(n_2791)
);

INVx4_ASAP7_75t_L g2792 ( 
.A(n_2380),
.Y(n_2792)
);

BUFx6f_ASAP7_75t_L g2793 ( 
.A(n_2380),
.Y(n_2793)
);

OAI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2651),
.A2(n_2277),
.B1(n_2256),
.B2(n_2262),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2717),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2431),
.B(n_2216),
.Y(n_2796)
);

INVx8_ASAP7_75t_L g2797 ( 
.A(n_2422),
.Y(n_2797)
);

INVx3_ASAP7_75t_L g2798 ( 
.A(n_2600),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2721),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2721),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2722),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_SL g2802 ( 
.A(n_2351),
.B(n_2210),
.Y(n_2802)
);

AOI22xp5_ASAP7_75t_L g2803 ( 
.A1(n_2422),
.A2(n_2426),
.B1(n_2489),
.B2(n_2510),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2722),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2354),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2724),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_SL g2807 ( 
.A(n_2492),
.Y(n_2807)
);

INVx3_ASAP7_75t_L g2808 ( 
.A(n_2616),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2484),
.B(n_2182),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2724),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_2431),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2726),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_L g2813 ( 
.A(n_2542),
.B(n_2193),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2726),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2727),
.Y(n_2815)
);

BUFx10_ASAP7_75t_L g2816 ( 
.A(n_2420),
.Y(n_2816)
);

BUFx2_ASAP7_75t_L g2817 ( 
.A(n_2711),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2367),
.Y(n_2818)
);

BUFx4f_ASAP7_75t_L g2819 ( 
.A(n_2755),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2727),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2730),
.Y(n_2821)
);

OAI22xp33_ASAP7_75t_L g2822 ( 
.A1(n_2654),
.A2(n_2277),
.B1(n_2256),
.B2(n_2262),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2658),
.B(n_2277),
.Y(n_2823)
);

NAND2xp33_ASAP7_75t_SL g2824 ( 
.A(n_2658),
.B(n_2251),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2730),
.Y(n_2825)
);

INVxp67_ASAP7_75t_SL g2826 ( 
.A(n_2369),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2659),
.B(n_2251),
.Y(n_2827)
);

OR2x2_ASAP7_75t_L g2828 ( 
.A(n_2490),
.B(n_2326),
.Y(n_2828)
);

AOI22xp33_ASAP7_75t_L g2829 ( 
.A1(n_2422),
.A2(n_2220),
.B1(n_2252),
.B2(n_2231),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2567),
.B(n_2216),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2742),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2659),
.B(n_2251),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_SL g2833 ( 
.A(n_2661),
.B(n_2251),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_SL g2834 ( 
.A(n_2661),
.B(n_2256),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2401),
.B(n_2405),
.Y(n_2835)
);

OAI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_2668),
.A2(n_2262),
.B1(n_2256),
.B2(n_2234),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_SL g2837 ( 
.A(n_2668),
.B(n_2256),
.Y(n_2837)
);

INVx5_ASAP7_75t_L g2838 ( 
.A(n_2340),
.Y(n_2838)
);

INVx3_ASAP7_75t_L g2839 ( 
.A(n_2616),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2747),
.Y(n_2840)
);

BUFx6f_ASAP7_75t_L g2841 ( 
.A(n_2380),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2411),
.B(n_2231),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2756),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2416),
.B(n_2231),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2482),
.B(n_2172),
.Y(n_2845)
);

NAND2xp33_ASAP7_75t_L g2846 ( 
.A(n_2672),
.B(n_2220),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2756),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2763),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2617),
.B(n_2179),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2763),
.Y(n_2850)
);

AOI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2422),
.A2(n_2220),
.B1(n_2252),
.B2(n_2091),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2422),
.A2(n_2220),
.B1(n_2252),
.B2(n_2232),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2766),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2766),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2509),
.B(n_2231),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2617),
.B(n_2493),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2672),
.B(n_2262),
.Y(n_2857)
);

INVx2_ASAP7_75t_SL g2858 ( 
.A(n_2510),
.Y(n_2858)
);

NAND2xp33_ASAP7_75t_SL g2859 ( 
.A(n_2675),
.B(n_2262),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2680),
.B(n_2232),
.Y(n_2860)
);

INVx3_ASAP7_75t_L g2861 ( 
.A(n_2616),
.Y(n_2861)
);

INVx4_ASAP7_75t_L g2862 ( 
.A(n_2380),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2769),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2769),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2496),
.B(n_2181),
.Y(n_2865)
);

INVx2_ASAP7_75t_SL g2866 ( 
.A(n_2510),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2622),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_2675),
.B(n_2175),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2623),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2555),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2437),
.Y(n_2871)
);

CKINVDCx5p33_ASAP7_75t_R g2872 ( 
.A(n_2450),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2683),
.B(n_2232),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2390),
.Y(n_2874)
);

BUFx6f_ASAP7_75t_SL g2875 ( 
.A(n_2555),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2437),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2699),
.B(n_2217),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2626),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_2616),
.Y(n_2879)
);

INVx2_ASAP7_75t_SL g2880 ( 
.A(n_2360),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2684),
.B(n_2232),
.Y(n_2881)
);

INVxp33_ASAP7_75t_L g2882 ( 
.A(n_2358),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2457),
.B(n_2258),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2628),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2631),
.Y(n_2885)
);

NOR2xp33_ASAP7_75t_L g2886 ( 
.A(n_2709),
.B(n_2248),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2435),
.B(n_2248),
.Y(n_2887)
);

AO22x2_ASAP7_75t_L g2888 ( 
.A1(n_2662),
.A2(n_2171),
.B1(n_1943),
.B2(n_2293),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2422),
.A2(n_2252),
.B1(n_2220),
.B2(n_2258),
.Y(n_2889)
);

AND3x2_ASAP7_75t_L g2890 ( 
.A(n_2366),
.B(n_2276),
.C(n_2253),
.Y(n_2890)
);

INVx4_ASAP7_75t_L g2891 ( 
.A(n_2390),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2633),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2636),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_SL g2894 ( 
.A(n_2452),
.B(n_2210),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2640),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2439),
.Y(n_2896)
);

AOI21x1_ASAP7_75t_L g2897 ( 
.A1(n_2753),
.A2(n_2002),
.B(n_2022),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2340),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2439),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2347),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2347),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_L g2902 ( 
.A(n_2451),
.B(n_2248),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2419),
.Y(n_2903)
);

OR2x6_ASAP7_75t_L g2904 ( 
.A(n_2755),
.B(n_2175),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2685),
.B(n_2258),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2352),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2352),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2382),
.Y(n_2908)
);

BUFx2_ASAP7_75t_L g2909 ( 
.A(n_2711),
.Y(n_2909)
);

AND3x2_ASAP7_75t_L g2910 ( 
.A(n_2551),
.B(n_2276),
.C(n_2253),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_SL g2911 ( 
.A(n_2453),
.B(n_2260),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2419),
.Y(n_2912)
);

CKINVDCx6p67_ASAP7_75t_R g2913 ( 
.A(n_2532),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2421),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2421),
.Y(n_2915)
);

NAND2xp33_ASAP7_75t_L g2916 ( 
.A(n_2688),
.B(n_2220),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2432),
.Y(n_2917)
);

BUFx10_ASAP7_75t_L g2918 ( 
.A(n_2454),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2382),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2397),
.Y(n_2920)
);

INVx8_ASAP7_75t_L g2921 ( 
.A(n_2426),
.Y(n_2921)
);

AND2x4_ASAP7_75t_L g2922 ( 
.A(n_2650),
.B(n_2057),
.Y(n_2922)
);

AOI22xp33_ASAP7_75t_L g2923 ( 
.A1(n_2426),
.A2(n_2252),
.B1(n_2279),
.B2(n_2258),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2432),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2688),
.B(n_2175),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2689),
.B(n_2176),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2397),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2433),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2433),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2445),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2445),
.Y(n_2931)
);

NOR2x1p5_ASAP7_75t_L g2932 ( 
.A(n_2629),
.B(n_2291),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2689),
.B(n_2176),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2462),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2462),
.Y(n_2935)
);

BUFx10_ASAP7_75t_L g2936 ( 
.A(n_2455),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2466),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2466),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2467),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2467),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2693),
.B(n_2176),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2468),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2472),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2472),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2481),
.Y(n_2945)
);

INVx5_ASAP7_75t_L g2946 ( 
.A(n_2340),
.Y(n_2946)
);

INVx3_ASAP7_75t_L g2947 ( 
.A(n_2340),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2481),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_L g2949 ( 
.A(n_2503),
.B(n_2270),
.Y(n_2949)
);

AND2x2_ASAP7_75t_SL g2950 ( 
.A(n_2743),
.B(n_2279),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2485),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2487),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2487),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_SL g2954 ( 
.A(n_2349),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2488),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2488),
.Y(n_2956)
);

AOI22xp33_ASAP7_75t_L g2957 ( 
.A1(n_2426),
.A2(n_2284),
.B1(n_2279),
.B2(n_1913),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2345),
.Y(n_2958)
);

INVx2_ASAP7_75t_SL g2959 ( 
.A(n_2360),
.Y(n_2959)
);

OAI22xp33_ASAP7_75t_SL g2960 ( 
.A1(n_2758),
.A2(n_2278),
.B1(n_2280),
.B2(n_2271),
.Y(n_2960)
);

INVxp67_ASAP7_75t_SL g2961 ( 
.A(n_2390),
.Y(n_2961)
);

OR2x6_ASAP7_75t_L g2962 ( 
.A(n_2755),
.B(n_2650),
.Y(n_2962)
);

XNOR2xp5_ASAP7_75t_L g2963 ( 
.A(n_2627),
.B(n_2132),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2506),
.Y(n_2964)
);

BUFx10_ASAP7_75t_L g2965 ( 
.A(n_2458),
.Y(n_2965)
);

INVx4_ASAP7_75t_L g2966 ( 
.A(n_2390),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2693),
.B(n_2176),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2557),
.B(n_2291),
.Y(n_2968)
);

INVx6_ASAP7_75t_L g2969 ( 
.A(n_2644),
.Y(n_2969)
);

AND2x2_ASAP7_75t_SL g2970 ( 
.A(n_2743),
.B(n_2284),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2515),
.Y(n_2971)
);

AOI21x1_ASAP7_75t_L g2972 ( 
.A1(n_2759),
.A2(n_2053),
.B(n_2107),
.Y(n_2972)
);

BUFx3_ASAP7_75t_L g2973 ( 
.A(n_2581),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2426),
.A2(n_2284),
.B1(n_1913),
.B2(n_1929),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2543),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2543),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2544),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2544),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2345),
.Y(n_2979)
);

NAND2xp33_ASAP7_75t_L g2980 ( 
.A(n_2695),
.B(n_2176),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2345),
.Y(n_2981)
);

INVx3_ASAP7_75t_L g2982 ( 
.A(n_2345),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2558),
.Y(n_2983)
);

INVx4_ASAP7_75t_L g2984 ( 
.A(n_2393),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2583),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2695),
.B(n_2191),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2583),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_2696),
.B(n_2191),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2587),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_SL g2990 ( 
.A(n_2696),
.B(n_2191),
.Y(n_2990)
);

INVx6_ASAP7_75t_L g2991 ( 
.A(n_2644),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2587),
.Y(n_2992)
);

INVxp67_ASAP7_75t_SL g2993 ( 
.A(n_2393),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2588),
.Y(n_2994)
);

AOI22xp33_ASAP7_75t_L g2995 ( 
.A1(n_2459),
.A2(n_2473),
.B1(n_2477),
.B2(n_2475),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2588),
.Y(n_2996)
);

INVxp33_ASAP7_75t_L g2997 ( 
.A(n_2655),
.Y(n_2997)
);

INVx2_ASAP7_75t_SL g2998 ( 
.A(n_2360),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2589),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2393),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_SL g3001 ( 
.A(n_2398),
.B(n_2260),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2478),
.B(n_2331),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2378),
.Y(n_3003)
);

CKINVDCx5p33_ASAP7_75t_R g3004 ( 
.A(n_2609),
.Y(n_3004)
);

CKINVDCx5p33_ASAP7_75t_R g3005 ( 
.A(n_2403),
.Y(n_3005)
);

NAND3xp33_ASAP7_75t_L g3006 ( 
.A(n_2765),
.B(n_2098),
.C(n_2139),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_2697),
.B(n_2191),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2610),
.Y(n_3008)
);

OR2x6_ASAP7_75t_L g3009 ( 
.A(n_2650),
.B(n_2191),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2610),
.Y(n_3010)
);

NAND2xp33_ASAP7_75t_L g3011 ( 
.A(n_2697),
.B(n_2201),
.Y(n_3011)
);

INVx3_ASAP7_75t_L g3012 ( 
.A(n_2378),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2480),
.B(n_2331),
.Y(n_3013)
);

INVx3_ASAP7_75t_L g3014 ( 
.A(n_2378),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2615),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_SL g3016 ( 
.A(n_2706),
.B(n_2707),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2618),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2691),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2618),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2645),
.Y(n_3020)
);

CKINVDCx5p33_ASAP7_75t_R g3021 ( 
.A(n_2403),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2700),
.B(n_2165),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2649),
.Y(n_3023)
);

INVx2_ASAP7_75t_SL g3024 ( 
.A(n_2691),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2499),
.B(n_2331),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2649),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2656),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2500),
.B(n_2292),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_2501),
.A2(n_1913),
.B1(n_1929),
.B2(n_1922),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2656),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2701),
.B(n_2702),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2703),
.B(n_2292),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2657),
.Y(n_3033)
);

INVx2_ASAP7_75t_SL g3034 ( 
.A(n_2691),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2338),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_SL g3036 ( 
.A(n_2706),
.B(n_2201),
.Y(n_3036)
);

BUFx3_ASAP7_75t_L g3037 ( 
.A(n_2599),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2704),
.B(n_2705),
.Y(n_3038)
);

OAI22xp33_ASAP7_75t_L g3039 ( 
.A1(n_2707),
.A2(n_2234),
.B1(n_2235),
.B2(n_2222),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2339),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2350),
.Y(n_3041)
);

BUFx3_ASAP7_75t_L g3042 ( 
.A(n_2638),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2356),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2362),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2708),
.B(n_2165),
.Y(n_3045)
);

BUFx10_ASAP7_75t_L g3046 ( 
.A(n_2597),
.Y(n_3046)
);

INVx1_ASAP7_75t_SL g3047 ( 
.A(n_2357),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2569),
.B(n_2292),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2375),
.Y(n_3049)
);

INVx5_ASAP7_75t_L g3050 ( 
.A(n_2378),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2417),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2669),
.Y(n_3052)
);

INVx4_ASAP7_75t_SL g3053 ( 
.A(n_2564),
.Y(n_3053)
);

BUFx6f_ASAP7_75t_SL g3054 ( 
.A(n_2349),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_2596),
.B(n_2298),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2423),
.Y(n_3056)
);

XNOR2x2_ASAP7_75t_SL g3057 ( 
.A(n_2637),
.B(n_2309),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2424),
.Y(n_3058)
);

OR2x6_ASAP7_75t_L g3059 ( 
.A(n_2761),
.B(n_2201),
.Y(n_3059)
);

INVx2_ASAP7_75t_SL g3060 ( 
.A(n_2739),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_SL g3061 ( 
.A(n_2714),
.B(n_2201),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2714),
.B(n_2201),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2425),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2427),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2428),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_L g3066 ( 
.A(n_2604),
.B(n_2298),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2429),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2365),
.B(n_2298),
.Y(n_3068)
);

OAI21xp33_ASAP7_75t_SL g3069 ( 
.A1(n_2534),
.A2(n_2190),
.B(n_2053),
.Y(n_3069)
);

BUFx6f_ASAP7_75t_L g3070 ( 
.A(n_2393),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2669),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2434),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2438),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2669),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2732),
.B(n_2203),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2710),
.B(n_2165),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2718),
.Y(n_3077)
);

INVx2_ASAP7_75t_SL g3078 ( 
.A(n_2739),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2441),
.Y(n_3079)
);

HB1xp67_ASAP7_75t_L g3080 ( 
.A(n_2387),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2718),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2715),
.B(n_2159),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2718),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2719),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2442),
.Y(n_3085)
);

INVx6_ASAP7_75t_L g3086 ( 
.A(n_2644),
.Y(n_3086)
);

INVxp33_ASAP7_75t_L g3087 ( 
.A(n_2698),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2443),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2719),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_SL g3090 ( 
.A(n_2733),
.B(n_2734),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_SL g3091 ( 
.A(n_2733),
.B(n_2203),
.Y(n_3091)
);

INVx4_ASAP7_75t_L g3092 ( 
.A(n_2409),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2735),
.Y(n_3093)
);

OAI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2734),
.A2(n_2302),
.B1(n_2299),
.B2(n_2235),
.Y(n_3094)
);

INVxp33_ASAP7_75t_L g3095 ( 
.A(n_2514),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_SL g3096 ( 
.A(n_2746),
.B(n_2203),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2735),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2746),
.B(n_2203),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2735),
.Y(n_3099)
);

AOI21x1_ASAP7_75t_L g3100 ( 
.A1(n_2768),
.A2(n_2113),
.B(n_2107),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2444),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2447),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2348),
.B(n_2012),
.Y(n_3103)
);

OAI21xp33_ASAP7_75t_SL g3104 ( 
.A1(n_2376),
.A2(n_2190),
.B(n_2045),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2770),
.Y(n_3105)
);

BUFx8_ASAP7_75t_SL g3106 ( 
.A(n_2342),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2449),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2563),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2563),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2775),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2646),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2754),
.B(n_2275),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2647),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2652),
.Y(n_3114)
);

INVx5_ASAP7_75t_L g3115 ( 
.A(n_2409),
.Y(n_3115)
);

NAND3xp33_ASAP7_75t_L g3116 ( 
.A(n_2359),
.B(n_2272),
.C(n_2236),
.Y(n_3116)
);

INVx4_ASAP7_75t_L g3117 ( 
.A(n_2415),
.Y(n_3117)
);

AND2x6_ASAP7_75t_L g3118 ( 
.A(n_2563),
.B(n_2296),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2764),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2653),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2667),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2348),
.B(n_2013),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2566),
.Y(n_3123)
);

OAI22x1_ASAP7_75t_L g3124 ( 
.A1(n_2398),
.A2(n_2310),
.B1(n_2315),
.B2(n_2294),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2566),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2670),
.Y(n_3126)
);

NAND2xp33_ASAP7_75t_L g3127 ( 
.A(n_2754),
.B(n_2771),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2415),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2566),
.Y(n_3129)
);

BUFx6f_ASAP7_75t_L g3130 ( 
.A(n_2415),
.Y(n_3130)
);

AO22x2_ASAP7_75t_L g3131 ( 
.A1(n_2607),
.A2(n_2171),
.B1(n_2635),
.B2(n_2310),
.Y(n_3131)
);

AND2x6_ASAP7_75t_L g3132 ( 
.A(n_2446),
.B(n_2296),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2731),
.B(n_2243),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2671),
.Y(n_3134)
);

CKINVDCx5p33_ASAP7_75t_R g3135 ( 
.A(n_2404),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2446),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2446),
.Y(n_3137)
);

INVx5_ASAP7_75t_L g3138 ( 
.A(n_2415),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2463),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_SL g3140 ( 
.A(n_2402),
.B(n_2260),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2463),
.Y(n_3141)
);

AOI21x1_ASAP7_75t_L g3142 ( 
.A1(n_2642),
.A2(n_2115),
.B(n_2113),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2463),
.Y(n_3143)
);

INVx5_ASAP7_75t_L g3144 ( 
.A(n_2456),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2476),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2476),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_2771),
.B(n_2243),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2720),
.Y(n_3148)
);

INVx6_ASAP7_75t_L g3149 ( 
.A(n_2644),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2723),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2476),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2725),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2737),
.B(n_2296),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_2383),
.B(n_2246),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2728),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2560),
.Y(n_3156)
);

BUFx3_ASAP7_75t_L g3157 ( 
.A(n_2716),
.Y(n_3157)
);

NAND3xp33_ASAP7_75t_L g3158 ( 
.A(n_2371),
.B(n_2289),
.C(n_2074),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2430),
.B(n_2027),
.Y(n_3159)
);

AOI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_2632),
.A2(n_2259),
.B1(n_2265),
.B2(n_2246),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2560),
.Y(n_3161)
);

NOR2xp33_ASAP7_75t_R g3162 ( 
.A(n_2776),
.B(n_1722),
.Y(n_3162)
);

CKINVDCx5p33_ASAP7_75t_R g3163 ( 
.A(n_2404),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_2471),
.B(n_2296),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2560),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2749),
.Y(n_3166)
);

INVx1_ASAP7_75t_SL g3167 ( 
.A(n_2519),
.Y(n_3167)
);

BUFx2_ASAP7_75t_L g3168 ( 
.A(n_2716),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2379),
.Y(n_3169)
);

INVx2_ASAP7_75t_SL g3170 ( 
.A(n_2739),
.Y(n_3170)
);

BUFx6f_ASAP7_75t_L g3171 ( 
.A(n_2456),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2386),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2389),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2392),
.Y(n_3174)
);

OR2x6_ASAP7_75t_L g3175 ( 
.A(n_2408),
.B(n_2170),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2395),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_SL g3177 ( 
.A1(n_2773),
.A2(n_2774),
.B1(n_2776),
.B2(n_2178),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2399),
.Y(n_3178)
);

NOR2x1p5_ASAP7_75t_L g3179 ( 
.A(n_2629),
.B(n_2178),
.Y(n_3179)
);

NOR3xp33_ASAP7_75t_L g3180 ( 
.A(n_2396),
.B(n_2335),
.C(n_2322),
.Y(n_3180)
);

BUFx2_ASAP7_75t_L g3181 ( 
.A(n_2740),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2400),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2641),
.B(n_2048),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2736),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2773),
.B(n_2259),
.Y(n_3185)
);

XNOR2xp5_ASAP7_75t_L g3186 ( 
.A(n_2355),
.B(n_2263),
.Y(n_3186)
);

NAND3xp33_ASAP7_75t_L g3187 ( 
.A(n_2410),
.B(n_2304),
.C(n_1979),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2511),
.B(n_2050),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2517),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2522),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2523),
.Y(n_3191)
);

BUFx2_ASAP7_75t_L g3192 ( 
.A(n_2740),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2526),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2736),
.Y(n_3194)
);

BUFx3_ASAP7_75t_L g3195 ( 
.A(n_2748),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2527),
.B(n_2050),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2736),
.Y(n_3197)
);

INVx1_ASAP7_75t_SL g3198 ( 
.A(n_2524),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2529),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2745),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2745),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2471),
.B(n_2300),
.Y(n_3202)
);

NAND3xp33_ASAP7_75t_L g3203 ( 
.A(n_2412),
.B(n_2051),
.C(n_2198),
.Y(n_3203)
);

NOR2x1p5_ASAP7_75t_L g3204 ( 
.A(n_2639),
.B(n_2178),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2530),
.Y(n_3205)
);

NOR2xp33_ASAP7_75t_L g3206 ( 
.A(n_2349),
.B(n_2265),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2531),
.B(n_2054),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_2774),
.B(n_2275),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2536),
.Y(n_3209)
);

INVx2_ASAP7_75t_SL g3210 ( 
.A(n_2767),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2745),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2546),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2553),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_2760),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_L g3215 ( 
.A(n_2611),
.B(n_2227),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2554),
.B(n_2054),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_SL g3217 ( 
.A(n_2440),
.B(n_2300),
.Y(n_3217)
);

INVx2_ASAP7_75t_SL g3218 ( 
.A(n_2767),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2565),
.B(n_2062),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2570),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2760),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_2520),
.B(n_2227),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_SL g3223 ( 
.A(n_2469),
.B(n_2300),
.Y(n_3223)
);

INVx2_ASAP7_75t_SL g3224 ( 
.A(n_2384),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2574),
.Y(n_3225)
);

INVxp33_ASAP7_75t_SL g3226 ( 
.A(n_2402),
.Y(n_3226)
);

NAND2xp33_ASAP7_75t_L g3227 ( 
.A(n_2665),
.B(n_2300),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_2483),
.B(n_2300),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2760),
.Y(n_3229)
);

NAND2xp33_ASAP7_75t_L g3230 ( 
.A(n_2665),
.B(n_2306),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2575),
.B(n_2576),
.Y(n_3231)
);

OAI21xp5_ASAP7_75t_L g3232 ( 
.A1(n_3069),
.A2(n_2772),
.B(n_2660),
.Y(n_3232)
);

XOR2x2_ASAP7_75t_L g3233 ( 
.A(n_2963),
.B(n_2712),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3111),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3111),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_SL g3236 ( 
.A(n_2805),
.B(n_2621),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3113),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3113),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3114),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2949),
.B(n_2245),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3114),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2845),
.B(n_2471),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3120),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3120),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3121),
.Y(n_3245)
);

NOR2xp33_ASAP7_75t_L g3246 ( 
.A(n_2856),
.B(n_2283),
.Y(n_3246)
);

BUFx3_ASAP7_75t_L g3247 ( 
.A(n_3157),
.Y(n_3247)
);

XOR2x2_ASAP7_75t_L g3248 ( 
.A(n_2963),
.B(n_2323),
.Y(n_3248)
);

NAND2xp33_ASAP7_75t_R g3249 ( 
.A(n_3162),
.B(n_2592),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3121),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_2809),
.B(n_2283),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3126),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2865),
.B(n_2582),
.Y(n_3253)
);

BUFx6f_ASAP7_75t_L g3254 ( 
.A(n_2793),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3126),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3134),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_2778),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3134),
.Y(n_3258)
);

NAND2x1p5_ASAP7_75t_L g3259 ( 
.A(n_2838),
.B(n_2407),
.Y(n_3259)
);

AND2x4_ASAP7_75t_L g3260 ( 
.A(n_2922),
.B(n_2729),
.Y(n_3260)
);

XOR2xp5_ASAP7_75t_L g3261 ( 
.A(n_3186),
.B(n_1759),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_2783),
.Y(n_3262)
);

CKINVDCx20_ASAP7_75t_R g3263 ( 
.A(n_3106),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_L g3264 ( 
.A(n_2813),
.B(n_2202),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3032),
.B(n_2552),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3035),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_2846),
.A2(n_2448),
.B(n_2436),
.Y(n_3267)
);

BUFx3_ASAP7_75t_L g3268 ( 
.A(n_3157),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3040),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3040),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3041),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2790),
.Y(n_3272)
);

AND2x2_ASAP7_75t_SL g3273 ( 
.A(n_2980),
.B(n_2448),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_3222),
.B(n_2594),
.Y(n_3274)
);

INVxp33_ASAP7_75t_SL g3275 ( 
.A(n_2805),
.Y(n_3275)
);

XNOR2xp5_ASAP7_75t_L g3276 ( 
.A(n_2882),
.B(n_1761),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3043),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3043),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3044),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3044),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3049),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3049),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3174),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3215),
.B(n_2605),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3174),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3176),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3176),
.Y(n_3287)
);

INVxp67_ASAP7_75t_L g3288 ( 
.A(n_3080),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_2916),
.A2(n_2663),
.B(n_2436),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2795),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3148),
.Y(n_3291)
);

INVxp67_ASAP7_75t_L g3292 ( 
.A(n_2968),
.Y(n_3292)
);

NOR2xp33_ASAP7_75t_L g3293 ( 
.A(n_2849),
.B(n_2299),
.Y(n_3293)
);

INVx4_ASAP7_75t_SL g3294 ( 
.A(n_3118),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3133),
.B(n_2614),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2877),
.B(n_2302),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3150),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3150),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3152),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3152),
.Y(n_3300)
);

XNOR2xp5_ASAP7_75t_L g3301 ( 
.A(n_3005),
.B(n_1761),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3155),
.Y(n_3302)
);

INVx2_ASAP7_75t_SL g3303 ( 
.A(n_2818),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2795),
.Y(n_3304)
);

NAND2xp33_ASAP7_75t_R g3305 ( 
.A(n_2817),
.B(n_2592),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3166),
.Y(n_3306)
);

BUFx6f_ASAP7_75t_L g3307 ( 
.A(n_2793),
.Y(n_3307)
);

CKINVDCx20_ASAP7_75t_R g3308 ( 
.A(n_2872),
.Y(n_3308)
);

NOR2xp67_ASAP7_75t_L g3309 ( 
.A(n_3116),
.B(n_2057),
.Y(n_3309)
);

AOI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2826),
.A2(n_2663),
.B(n_1975),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_3055),
.B(n_3066),
.Y(n_3311)
);

CKINVDCx5p33_ASAP7_75t_R g3312 ( 
.A(n_3021),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3169),
.Y(n_3313)
);

XOR2xp5_ASAP7_75t_L g3314 ( 
.A(n_3135),
.B(n_1765),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3172),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_2799),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3172),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3173),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3173),
.Y(n_3319)
);

OR2x2_ASAP7_75t_L g3320 ( 
.A(n_2828),
.B(n_2294),
.Y(n_3320)
);

AND2x4_ASAP7_75t_L g3321 ( 
.A(n_2922),
.B(n_2385),
.Y(n_3321)
);

CKINVDCx20_ASAP7_75t_R g3322 ( 
.A(n_2913),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3178),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3178),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_2828),
.B(n_2315),
.Y(n_3325)
);

BUFx5_ASAP7_75t_L g3326 ( 
.A(n_3118),
.Y(n_3326)
);

OAI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2781),
.A2(n_2692),
.B(n_2123),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3182),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3182),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3189),
.Y(n_3330)
);

NOR2xp33_ASAP7_75t_L g3331 ( 
.A(n_3095),
.B(n_2271),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3068),
.B(n_2278),
.Y(n_3332)
);

AOI21x1_ASAP7_75t_L g3333 ( 
.A1(n_3100),
.A2(n_2738),
.B(n_2690),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3190),
.Y(n_3334)
);

XNOR2x2_ASAP7_75t_L g3335 ( 
.A(n_3131),
.B(n_2005),
.Y(n_3335)
);

INVxp33_ASAP7_75t_L g3336 ( 
.A(n_3154),
.Y(n_3336)
);

XNOR2x2_ASAP7_75t_L g3337 ( 
.A(n_3131),
.B(n_1029),
.Y(n_3337)
);

INVx1_ASAP7_75t_SL g3338 ( 
.A(n_3047),
.Y(n_3338)
);

XOR2xp5_ASAP7_75t_L g3339 ( 
.A(n_3135),
.B(n_1776),
.Y(n_3339)
);

XOR2x2_ASAP7_75t_L g3340 ( 
.A(n_3180),
.B(n_1945),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3191),
.Y(n_3341)
);

NOR2xp33_ASAP7_75t_L g3342 ( 
.A(n_3082),
.B(n_2887),
.Y(n_3342)
);

BUFx5_ASAP7_75t_L g3343 ( 
.A(n_3118),
.Y(n_3343)
);

INVxp33_ASAP7_75t_L g3344 ( 
.A(n_2784),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3193),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_2902),
.B(n_2280),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3199),
.Y(n_3347)
);

XOR2x2_ASAP7_75t_L g3348 ( 
.A(n_3006),
.B(n_1945),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3205),
.Y(n_3349)
);

XOR2xp5_ASAP7_75t_L g3350 ( 
.A(n_3163),
.B(n_1776),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3205),
.Y(n_3351)
);

XNOR2x2_ASAP7_75t_L g3352 ( 
.A(n_3131),
.B(n_1029),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3209),
.Y(n_3353)
);

CKINVDCx16_ASAP7_75t_R g3354 ( 
.A(n_2816),
.Y(n_3354)
);

INVx2_ASAP7_75t_SL g3355 ( 
.A(n_2818),
.Y(n_3355)
);

XOR2x2_ASAP7_75t_L g3356 ( 
.A(n_2890),
.B(n_2141),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3212),
.Y(n_3357)
);

INVx2_ASAP7_75t_SL g3358 ( 
.A(n_3195),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2804),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3212),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3213),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_3048),
.B(n_2285),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_2804),
.Y(n_3363)
);

CKINVDCx16_ASAP7_75t_R g3364 ( 
.A(n_2816),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3220),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3220),
.Y(n_3366)
);

XNOR2x2_ASAP7_75t_L g3367 ( 
.A(n_3131),
.B(n_637),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3225),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_2836),
.B(n_2170),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3225),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_2782),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_3028),
.B(n_2285),
.Y(n_3372)
);

CKINVDCx20_ASAP7_75t_R g3373 ( 
.A(n_3004),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2788),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_2788),
.Y(n_3375)
);

INVxp67_ASAP7_75t_SL g3376 ( 
.A(n_2930),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3028),
.B(n_2250),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2791),
.Y(n_3378)
);

XOR2x2_ASAP7_75t_L g3379 ( 
.A(n_3158),
.B(n_2174),
.Y(n_3379)
);

AND2x4_ASAP7_75t_L g3380 ( 
.A(n_3164),
.B(n_2414),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2791),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_2810),
.Y(n_3382)
);

INVxp33_ASAP7_75t_L g3383 ( 
.A(n_2817),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_2810),
.Y(n_3384)
);

XOR2xp5_ASAP7_75t_L g3385 ( 
.A(n_3163),
.B(n_1788),
.Y(n_3385)
);

CKINVDCx5p33_ASAP7_75t_R g3386 ( 
.A(n_3004),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2800),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2812),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_2830),
.B(n_2584),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_2801),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_2801),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_2806),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2806),
.Y(n_3393)
);

OR2x6_ASAP7_75t_L g3394 ( 
.A(n_2962),
.B(n_2135),
.Y(n_3394)
);

INVx4_ASAP7_75t_SL g3395 ( 
.A(n_3118),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2815),
.Y(n_3396)
);

OR2x2_ASAP7_75t_L g3397 ( 
.A(n_3167),
.B(n_2327),
.Y(n_3397)
);

NOR2xp33_ASAP7_75t_L g3398 ( 
.A(n_3187),
.B(n_2066),
.Y(n_3398)
);

AND2x6_ASAP7_75t_L g3399 ( 
.A(n_2852),
.B(n_2679),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2930),
.B(n_2590),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_2815),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_2821),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_2812),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2821),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2825),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2934),
.B(n_2591),
.Y(n_3406)
);

INVx2_ASAP7_75t_SL g3407 ( 
.A(n_2909),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2825),
.Y(n_3408)
);

AND2x2_ASAP7_75t_SL g3409 ( 
.A(n_3011),
.B(n_2486),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_SL g3410 ( 
.A(n_3226),
.B(n_2624),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_3206),
.B(n_2287),
.Y(n_3411)
);

CKINVDCx20_ASAP7_75t_R g3412 ( 
.A(n_2913),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_2814),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2934),
.B(n_2593),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2831),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_2814),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_2847),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_2935),
.B(n_2598),
.Y(n_3418)
);

OR2x2_ASAP7_75t_SL g3419 ( 
.A(n_3203),
.B(n_2538),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2848),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2848),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_2820),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_2853),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_2853),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_2864),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_2864),
.Y(n_3426)
);

CKINVDCx5p33_ASAP7_75t_R g3427 ( 
.A(n_2779),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3051),
.Y(n_3428)
);

INVxp67_ASAP7_75t_L g3429 ( 
.A(n_3153),
.Y(n_3429)
);

AND2x2_ASAP7_75t_SL g3430 ( 
.A(n_2950),
.B(n_2970),
.Y(n_3430)
);

AND2x4_ASAP7_75t_L g3431 ( 
.A(n_3164),
.B(n_2491),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3056),
.Y(n_3432)
);

NOR2xp33_ASAP7_75t_L g3433 ( 
.A(n_3112),
.B(n_2508),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3056),
.Y(n_3434)
);

INVxp33_ASAP7_75t_L g3435 ( 
.A(n_3168),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3058),
.Y(n_3436)
);

INVx4_ASAP7_75t_L g3437 ( 
.A(n_2962),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_3147),
.B(n_2516),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_L g3439 ( 
.A(n_3185),
.B(n_2547),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3063),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3063),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_L g3442 ( 
.A(n_3208),
.B(n_2571),
.Y(n_3442)
);

INVx2_ASAP7_75t_SL g3443 ( 
.A(n_3168),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_2786),
.B(n_2572),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3064),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3183),
.A2(n_1975),
.B(n_2407),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3064),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3202),
.B(n_2507),
.Y(n_3448)
);

INVxp33_ASAP7_75t_L g3449 ( 
.A(n_3181),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3065),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3067),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3072),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3072),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_2935),
.B(n_2603),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_3226),
.Y(n_3455)
);

CKINVDCx5p33_ASAP7_75t_R g3456 ( 
.A(n_2816),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3202),
.B(n_2528),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_2886),
.B(n_2548),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3073),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3073),
.Y(n_3460)
);

XNOR2xp5_ASAP7_75t_L g3461 ( 
.A(n_3057),
.B(n_1804),
.Y(n_3461)
);

CKINVDCx16_ASAP7_75t_R g3462 ( 
.A(n_2918),
.Y(n_3462)
);

XOR2xp5_ASAP7_75t_L g3463 ( 
.A(n_2997),
.B(n_1804),
.Y(n_3463)
);

AND2x2_ASAP7_75t_L g3464 ( 
.A(n_2973),
.B(n_2630),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3079),
.Y(n_3465)
);

AOI21x1_ASAP7_75t_L g3466 ( 
.A1(n_3100),
.A2(n_2677),
.B(n_2121),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_2973),
.B(n_2634),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3079),
.Y(n_3468)
);

AND2x4_ASAP7_75t_L g3469 ( 
.A(n_3037),
.B(n_2664),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3085),
.Y(n_3470)
);

INVx4_ASAP7_75t_L g3471 ( 
.A(n_2962),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_L g3472 ( 
.A(n_3016),
.B(n_2577),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3090),
.B(n_2106),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_2937),
.B(n_2613),
.Y(n_3474)
);

AND2x2_ASAP7_75t_SL g3475 ( 
.A(n_2950),
.B(n_2666),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3085),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_3087),
.B(n_2308),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_SL g3478 ( 
.A(n_3177),
.B(n_2173),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3088),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3088),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_3039),
.B(n_2639),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3101),
.Y(n_3482)
);

BUFx8_ASAP7_75t_L g3483 ( 
.A(n_2954),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2838),
.A2(n_2494),
.B(n_2407),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_2840),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3101),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_2843),
.Y(n_3487)
);

INVxp33_ASAP7_75t_L g3488 ( 
.A(n_3181),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3102),
.Y(n_3489)
);

INVx4_ASAP7_75t_L g3490 ( 
.A(n_2962),
.Y(n_3490)
);

INVx3_ASAP7_75t_L g3491 ( 
.A(n_2792),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3102),
.Y(n_3492)
);

INVxp67_ASAP7_75t_SL g3493 ( 
.A(n_2937),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3107),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3107),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3110),
.Y(n_3496)
);

INVxp67_ASAP7_75t_SL g3497 ( 
.A(n_2938),
.Y(n_3497)
);

AND2x4_ASAP7_75t_L g3498 ( 
.A(n_3037),
.B(n_2545),
.Y(n_3498)
);

NOR2xp33_ASAP7_75t_L g3499 ( 
.A(n_2880),
.B(n_2643),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3110),
.Y(n_3500)
);

XOR2xp5_ASAP7_75t_L g3501 ( 
.A(n_3192),
.B(n_1813),
.Y(n_3501)
);

AOI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_2838),
.A2(n_2559),
.B(n_2494),
.Y(n_3502)
);

INVxp33_ASAP7_75t_L g3503 ( 
.A(n_3192),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_2867),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_2869),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_2938),
.B(n_2620),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_2942),
.B(n_2545),
.Y(n_3507)
);

NAND2xp33_ASAP7_75t_R g3508 ( 
.A(n_2796),
.B(n_2537),
.Y(n_3508)
);

NOR2xp33_ASAP7_75t_SL g3509 ( 
.A(n_2802),
.B(n_2625),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2878),
.Y(n_3510)
);

CKINVDCx20_ASAP7_75t_R g3511 ( 
.A(n_2918),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_2850),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_2884),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_2884),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_2885),
.Y(n_3515)
);

XNOR2x2_ASAP7_75t_L g3516 ( 
.A(n_2888),
.B(n_637),
.Y(n_3516)
);

AND2x4_ASAP7_75t_L g3517 ( 
.A(n_3042),
.B(n_2545),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_2885),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_2892),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_2850),
.Y(n_3520)
);

CKINVDCx20_ASAP7_75t_R g3521 ( 
.A(n_2936),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_2880),
.B(n_2643),
.Y(n_3522)
);

OAI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_2842),
.A2(n_2860),
.B(n_2844),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_2893),
.Y(n_3524)
);

NAND2x1p5_ASAP7_75t_L g3525 ( 
.A(n_2838),
.B(n_2494),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_2895),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_2895),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_2854),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_2854),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_2863),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2863),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_2942),
.B(n_2550),
.Y(n_3532)
);

NOR2xp67_ASAP7_75t_L g3533 ( 
.A(n_3160),
.B(n_2249),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_2835),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_2943),
.B(n_2550),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3031),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3038),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_2943),
.Y(n_3538)
);

NOR2xp67_ASAP7_75t_L g3539 ( 
.A(n_3094),
.B(n_2249),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_2944),
.B(n_2550),
.Y(n_3540)
);

OAI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_2873),
.A2(n_2413),
.B(n_2384),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3052),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_2944),
.Y(n_3543)
);

AND2x4_ASAP7_75t_L g3544 ( 
.A(n_3119),
.B(n_2384),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_2945),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_2794),
.B(n_2184),
.Y(n_3546)
);

INVxp33_ASAP7_75t_L g3547 ( 
.A(n_2894),
.Y(n_3547)
);

OR2x2_ASAP7_75t_L g3548 ( 
.A(n_3198),
.B(n_2309),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_2945),
.Y(n_3549)
);

AOI21x1_ASAP7_75t_L g3550 ( 
.A1(n_2972),
.A2(n_2121),
.B(n_2115),
.Y(n_3550)
);

NAND2xp33_ASAP7_75t_R g3551 ( 
.A(n_2796),
.B(n_2537),
.Y(n_3551)
);

AND2x6_ASAP7_75t_L g3552 ( 
.A(n_2851),
.B(n_2780),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_2948),
.Y(n_3553)
);

AND2x2_ASAP7_75t_L g3554 ( 
.A(n_3119),
.B(n_2184),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_2995),
.B(n_2185),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_2948),
.Y(n_3556)
);

OR2x6_ASAP7_75t_L g3557 ( 
.A(n_3009),
.B(n_2135),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3052),
.Y(n_3558)
);

OR2x2_ASAP7_75t_L g3559 ( 
.A(n_3231),
.B(n_2311),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_2951),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_2951),
.Y(n_3561)
);

INVx1_ASAP7_75t_SL g3562 ( 
.A(n_2936),
.Y(n_3562)
);

AND2x4_ASAP7_75t_L g3563 ( 
.A(n_3009),
.B(n_2413),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_2953),
.Y(n_3564)
);

XOR2x2_ASAP7_75t_L g3565 ( 
.A(n_2910),
.B(n_2324),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_2953),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_2956),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_2956),
.Y(n_3568)
);

XOR2xp5_ASAP7_75t_L g3569 ( 
.A(n_2888),
.B(n_1831),
.Y(n_3569)
);

INVx3_ASAP7_75t_L g3570 ( 
.A(n_2792),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_2964),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_2971),
.Y(n_3572)
);

AND2x4_ASAP7_75t_L g3573 ( 
.A(n_3009),
.B(n_2413),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_2971),
.B(n_2021),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_2975),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3224),
.B(n_2185),
.Y(n_3576)
);

NAND2xp33_ASAP7_75t_R g3577 ( 
.A(n_2898),
.B(n_2540),
.Y(n_3577)
);

AND2x2_ASAP7_75t_L g3578 ( 
.A(n_3224),
.B(n_2189),
.Y(n_3578)
);

BUFx6f_ASAP7_75t_L g3579 ( 
.A(n_2793),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_2975),
.Y(n_3580)
);

AND2x4_ASAP7_75t_L g3581 ( 
.A(n_3009),
.B(n_2748),
.Y(n_3581)
);

NAND2xp33_ASAP7_75t_SL g3582 ( 
.A(n_2785),
.B(n_2306),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_2976),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_2976),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_2838),
.A2(n_2579),
.B(n_2559),
.Y(n_3585)
);

XNOR2x2_ASAP7_75t_L g3586 ( 
.A(n_2888),
.B(n_683),
.Y(n_3586)
);

NOR2xp33_ASAP7_75t_L g3587 ( 
.A(n_2959),
.B(n_2230),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_2977),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_2998),
.B(n_2233),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_2998),
.B(n_2209),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_2978),
.Y(n_3591)
);

INVx3_ASAP7_75t_R g3592 ( 
.A(n_2965),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_2978),
.Y(n_3593)
);

AND2x2_ASAP7_75t_L g3594 ( 
.A(n_2932),
.B(n_2209),
.Y(n_3594)
);

INVxp33_ASAP7_75t_L g3595 ( 
.A(n_2911),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_2983),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_2838),
.A2(n_2579),
.B(n_2559),
.Y(n_3597)
);

XOR2xp5_ASAP7_75t_L g3598 ( 
.A(n_2888),
.B(n_1842),
.Y(n_3598)
);

XNOR2xp5_ASAP7_75t_L g3599 ( 
.A(n_3179),
.B(n_1842),
.Y(n_3599)
);

CKINVDCx20_ASAP7_75t_R g3600 ( 
.A(n_2965),
.Y(n_3600)
);

OR2x2_ASAP7_75t_L g3601 ( 
.A(n_3188),
.B(n_2311),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_2983),
.Y(n_3602)
);

INVxp67_ASAP7_75t_SL g3603 ( 
.A(n_2985),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_2985),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3179),
.B(n_2213),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_2987),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_2987),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_L g3608 ( 
.A(n_3223),
.B(n_2237),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_3228),
.B(n_2239),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_2989),
.Y(n_3610)
);

INVx4_ASAP7_75t_SL g3611 ( 
.A(n_3118),
.Y(n_3611)
);

OR2x2_ASAP7_75t_L g3612 ( 
.A(n_3196),
.B(n_2312),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3204),
.B(n_2214),
.Y(n_3613)
);

CKINVDCx20_ASAP7_75t_R g3614 ( 
.A(n_2965),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_2989),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_SL g3616 ( 
.A(n_3242),
.B(n_2822),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3330),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_L g3618 ( 
.A1(n_3348),
.A2(n_2381),
.B1(n_3013),
.B2(n_3002),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3542),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3342),
.B(n_3127),
.Y(n_3620)
);

INVx3_ASAP7_75t_L g3621 ( 
.A(n_3437),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3558),
.Y(n_3622)
);

INVx2_ASAP7_75t_SL g3623 ( 
.A(n_3247),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3342),
.B(n_3013),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3242),
.B(n_2960),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3334),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3311),
.B(n_3002),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3311),
.B(n_3025),
.Y(n_3628)
);

INVx2_ASAP7_75t_SL g3629 ( 
.A(n_3268),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3534),
.B(n_3025),
.Y(n_3630)
);

NOR2xp33_ASAP7_75t_L g3631 ( 
.A(n_3336),
.B(n_2312),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_SL g3632 ( 
.A(n_3444),
.B(n_2824),
.Y(n_3632)
);

INVx5_ASAP7_75t_L g3633 ( 
.A(n_3254),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3341),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3536),
.B(n_2883),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_L g3636 ( 
.A(n_3336),
.B(n_2319),
.Y(n_3636)
);

BUFx8_ASAP7_75t_L g3637 ( 
.A(n_3407),
.Y(n_3637)
);

BUFx2_ASAP7_75t_L g3638 ( 
.A(n_3338),
.Y(n_3638)
);

INVx2_ASAP7_75t_SL g3639 ( 
.A(n_3303),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_L g3640 ( 
.A(n_3251),
.B(n_2319),
.Y(n_3640)
);

INVxp67_ASAP7_75t_SL g3641 ( 
.A(n_3376),
.Y(n_3641)
);

NOR2xp67_ASAP7_75t_L g3642 ( 
.A(n_3386),
.B(n_2249),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3537),
.B(n_3253),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3253),
.B(n_2883),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_L g3645 ( 
.A(n_3251),
.B(n_2324),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3289),
.A2(n_3310),
.B(n_3050),
.Y(n_3646)
);

AND2x4_ASAP7_75t_SL g3647 ( 
.A(n_3308),
.B(n_3046),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_SL g3648 ( 
.A(n_3331),
.B(n_2306),
.Y(n_3648)
);

INVx2_ASAP7_75t_SL g3649 ( 
.A(n_3355),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3296),
.B(n_3103),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3257),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3296),
.B(n_3122),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3264),
.A2(n_2525),
.B1(n_2541),
.B2(n_2540),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3346),
.B(n_2777),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_3246),
.B(n_2324),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3262),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3346),
.B(n_2777),
.Y(n_3657)
);

O2A1O1Ixp5_ASAP7_75t_L g3658 ( 
.A1(n_3546),
.A2(n_3369),
.B(n_3478),
.C(n_3232),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3293),
.B(n_2811),
.Y(n_3659)
);

NOR2xp33_ASAP7_75t_L g3660 ( 
.A(n_3246),
.B(n_2320),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3293),
.B(n_2320),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3240),
.B(n_2811),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3272),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3379),
.A2(n_2381),
.B1(n_3124),
.B2(n_2855),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3332),
.B(n_2868),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3444),
.B(n_2859),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3264),
.B(n_2925),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3362),
.B(n_2926),
.Y(n_3668)
);

INVx3_ASAP7_75t_L g3669 ( 
.A(n_3437),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3265),
.B(n_2933),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3295),
.B(n_2941),
.Y(n_3671)
);

NOR2xp33_ASAP7_75t_L g3672 ( 
.A(n_3331),
.B(n_2321),
.Y(n_3672)
);

AND2x2_ASAP7_75t_SL g3673 ( 
.A(n_3430),
.B(n_2970),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3284),
.B(n_2967),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3290),
.Y(n_3675)
);

AOI22xp33_ASAP7_75t_L g3676 ( 
.A1(n_3516),
.A2(n_3124),
.B1(n_2855),
.B2(n_3217),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3304),
.Y(n_3677)
);

INVx2_ASAP7_75t_SL g3678 ( 
.A(n_3554),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3316),
.Y(n_3679)
);

NOR2xp33_ASAP7_75t_L g3680 ( 
.A(n_3292),
.B(n_2321),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_L g3681 ( 
.A1(n_3586),
.A2(n_2905),
.B1(n_2881),
.B2(n_2832),
.Y(n_3681)
);

O2A1O1Ixp33_ASAP7_75t_L g3682 ( 
.A1(n_3478),
.A2(n_2218),
.B(n_2224),
.C(n_2221),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3274),
.B(n_2986),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3472),
.B(n_2988),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3472),
.B(n_2990),
.Y(n_3685)
);

AOI22xp33_ASAP7_75t_L g3686 ( 
.A1(n_3367),
.A2(n_2833),
.B1(n_2834),
.B2(n_2827),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3359),
.Y(n_3687)
);

OAI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3475),
.A2(n_3059),
.B1(n_2819),
.B2(n_2904),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_3411),
.B(n_2306),
.Y(n_3689)
);

OAI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3475),
.A2(n_3059),
.B1(n_2819),
.B2(n_2904),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_SL g3691 ( 
.A(n_3411),
.B(n_2306),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3433),
.B(n_3007),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_SL g3693 ( 
.A(n_3509),
.B(n_3001),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3433),
.B(n_3036),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3438),
.B(n_3439),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3438),
.B(n_2334),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3439),
.B(n_3442),
.Y(n_3697)
);

AO221x1_ASAP7_75t_L g3698 ( 
.A1(n_3337),
.A2(n_2219),
.B1(n_2334),
.B2(n_2247),
.C(n_2255),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3442),
.B(n_3061),
.Y(n_3699)
);

OAI22xp5_ASAP7_75t_SL g3700 ( 
.A1(n_3461),
.A2(n_2602),
.B1(n_2595),
.B2(n_1856),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3345),
.Y(n_3701)
);

INVx8_ASAP7_75t_L g3702 ( 
.A(n_3394),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3363),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3372),
.B(n_3062),
.Y(n_3704)
);

BUFx6f_ASAP7_75t_L g3705 ( 
.A(n_3254),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3382),
.Y(n_3706)
);

A2O1A1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_3398),
.A2(n_3104),
.B(n_2803),
.C(n_2889),
.Y(n_3707)
);

NOR2x2_ASAP7_75t_L g3708 ( 
.A(n_3352),
.B(n_2408),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3458),
.B(n_3075),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3555),
.B(n_3091),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_L g3711 ( 
.A1(n_3340),
.A2(n_3335),
.B1(n_3369),
.B2(n_3481),
.Y(n_3711)
);

NAND3xp33_ASAP7_75t_L g3712 ( 
.A(n_3477),
.B(n_2406),
.C(n_2257),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3448),
.B(n_3457),
.Y(n_3713)
);

NOR2xp67_ASAP7_75t_L g3714 ( 
.A(n_3427),
.B(n_2249),
.Y(n_3714)
);

AOI22xp33_ASAP7_75t_L g3715 ( 
.A1(n_3481),
.A2(n_2857),
.B1(n_2837),
.B2(n_3096),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3384),
.Y(n_3716)
);

INVx2_ASAP7_75t_SL g3717 ( 
.A(n_3443),
.Y(n_3717)
);

AOI22xp33_ASAP7_75t_L g3718 ( 
.A1(n_3569),
.A2(n_3098),
.B1(n_3175),
.B2(n_725),
.Y(n_3718)
);

AOI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3477),
.A2(n_2549),
.B1(n_2541),
.B2(n_2752),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3347),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_SL g3721 ( 
.A(n_3473),
.B(n_3140),
.Y(n_3721)
);

INVxp67_ASAP7_75t_SL g3722 ( 
.A(n_3376),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_SL g3723 ( 
.A(n_3473),
.B(n_2241),
.Y(n_3723)
);

AOI22xp5_ASAP7_75t_L g3724 ( 
.A1(n_3499),
.A2(n_2549),
.B1(n_2762),
.B2(n_2752),
.Y(n_3724)
);

OAI22xp5_ASAP7_75t_L g3725 ( 
.A1(n_3409),
.A2(n_3059),
.B1(n_2904),
.B2(n_2829),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_SL g3726 ( 
.A(n_3377),
.B(n_2266),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3383),
.B(n_3435),
.Y(n_3727)
);

NOR2xp33_ASAP7_75t_L g3728 ( 
.A(n_3383),
.B(n_3435),
.Y(n_3728)
);

INVx2_ASAP7_75t_SL g3729 ( 
.A(n_3358),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3429),
.B(n_3207),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3349),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3499),
.A2(n_2762),
.B1(n_2269),
.B2(n_2268),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3351),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_SL g3734 ( 
.A(n_3544),
.B(n_2205),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3429),
.B(n_3216),
.Y(n_3735)
);

HB1xp67_ASAP7_75t_L g3736 ( 
.A(n_3288),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3353),
.Y(n_3737)
);

INVx4_ASAP7_75t_L g3738 ( 
.A(n_3394),
.Y(n_3738)
);

INVx4_ASAP7_75t_L g3739 ( 
.A(n_3394),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3380),
.B(n_3219),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3357),
.Y(n_3741)
);

NOR2xp67_ASAP7_75t_L g3742 ( 
.A(n_3455),
.B(n_2206),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3320),
.B(n_2334),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3360),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3431),
.B(n_3159),
.Y(n_3745)
);

AND2x4_ASAP7_75t_L g3746 ( 
.A(n_3471),
.B(n_2870),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3388),
.Y(n_3747)
);

AOI22xp33_ASAP7_75t_L g3748 ( 
.A1(n_3598),
.A2(n_3175),
.B1(n_725),
.B2(n_830),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3431),
.B(n_2858),
.Y(n_3749)
);

NOR2xp33_ASAP7_75t_L g3750 ( 
.A(n_3449),
.B(n_2183),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_SL g3751 ( 
.A(n_3544),
.B(n_3498),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_SL g3752 ( 
.A(n_3498),
.B(n_2497),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3361),
.Y(n_3753)
);

AOI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3522),
.A2(n_2533),
.B1(n_2518),
.B2(n_2474),
.Y(n_3754)
);

AOI22xp33_ASAP7_75t_L g3755 ( 
.A1(n_3356),
.A2(n_3175),
.B1(n_830),
.B2(n_861),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3590),
.B(n_2866),
.Y(n_3756)
);

AOI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_3522),
.A2(n_2533),
.B1(n_2518),
.B2(n_2474),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3587),
.B(n_2866),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3587),
.B(n_2785),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3365),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3589),
.B(n_3204),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3366),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_SL g3763 ( 
.A(n_3517),
.B(n_2608),
.Y(n_3763)
);

OR2x6_ASAP7_75t_L g3764 ( 
.A(n_3471),
.B(n_2797),
.Y(n_3764)
);

BUFx3_ASAP7_75t_L g3765 ( 
.A(n_3275),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3368),
.Y(n_3766)
);

INVx3_ASAP7_75t_L g3767 ( 
.A(n_3490),
.Y(n_3767)
);

OAI22xp5_ASAP7_75t_L g3768 ( 
.A1(n_3493),
.A2(n_2923),
.B1(n_2957),
.B2(n_2974),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3449),
.B(n_3488),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3589),
.B(n_2870),
.Y(n_3770)
);

OR2x2_ASAP7_75t_L g3771 ( 
.A(n_3325),
.B(n_2290),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3464),
.B(n_2295),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3389),
.B(n_3071),
.Y(n_3773)
);

OAI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_3493),
.A2(n_3175),
.B1(n_3050),
.B2(n_2946),
.Y(n_3774)
);

NOR2xp33_ASAP7_75t_L g3775 ( 
.A(n_3488),
.B(n_2183),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3389),
.B(n_3074),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3576),
.B(n_3074),
.Y(n_3777)
);

NOR2xp67_ASAP7_75t_L g3778 ( 
.A(n_3312),
.B(n_2573),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3578),
.B(n_3077),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3403),
.Y(n_3780)
);

AOI22xp33_ASAP7_75t_L g3781 ( 
.A1(n_3399),
.A2(n_830),
.B1(n_861),
.B2(n_777),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_SL g3782 ( 
.A(n_3517),
.B(n_2353),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3370),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3413),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3608),
.B(n_3609),
.Y(n_3785)
);

INVx2_ASAP7_75t_SL g3786 ( 
.A(n_3397),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_SL g3787 ( 
.A(n_3430),
.B(n_3022),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3609),
.B(n_3077),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_SL g3789 ( 
.A(n_3547),
.B(n_2353),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_SL g3790 ( 
.A(n_3547),
.B(n_2295),
.Y(n_3790)
);

NOR2xp33_ASAP7_75t_SL g3791 ( 
.A(n_3236),
.B(n_2495),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3291),
.Y(n_3792)
);

NOR2xp33_ASAP7_75t_L g3793 ( 
.A(n_3503),
.B(n_2192),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3297),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3298),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3601),
.B(n_3612),
.Y(n_3796)
);

BUFx6f_ASAP7_75t_L g3797 ( 
.A(n_3254),
.Y(n_3797)
);

NOR2xp33_ASAP7_75t_L g3798 ( 
.A(n_3503),
.B(n_2192),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3559),
.B(n_3081),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3299),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3497),
.B(n_3081),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_L g3802 ( 
.A(n_3548),
.B(n_2196),
.Y(n_3802)
);

INVx5_ASAP7_75t_L g3803 ( 
.A(n_3254),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3300),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3497),
.B(n_3083),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3467),
.B(n_2303),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3603),
.B(n_3083),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_3581),
.B(n_2303),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3416),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3422),
.Y(n_3810)
);

OR2x6_ASAP7_75t_L g3811 ( 
.A(n_3490),
.B(n_2797),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3302),
.B(n_3084),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3541),
.B(n_3045),
.Y(n_3813)
);

INVxp67_ASAP7_75t_L g3814 ( 
.A(n_3577),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_SL g3815 ( 
.A(n_3309),
.B(n_3076),
.Y(n_3815)
);

NOR2xp67_ASAP7_75t_L g3816 ( 
.A(n_3456),
.B(n_2573),
.Y(n_3816)
);

NOR2xp33_ASAP7_75t_L g3817 ( 
.A(n_3344),
.B(n_2196),
.Y(n_3817)
);

INVx3_ASAP7_75t_L g3818 ( 
.A(n_3491),
.Y(n_3818)
);

INVx1_ASAP7_75t_SL g3819 ( 
.A(n_3344),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3306),
.B(n_3089),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_SL g3821 ( 
.A(n_3273),
.B(n_2946),
.Y(n_3821)
);

BUFx6f_ASAP7_75t_L g3822 ( 
.A(n_3307),
.Y(n_3822)
);

AND2x4_ASAP7_75t_L g3823 ( 
.A(n_3469),
.B(n_3018),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3273),
.B(n_2946),
.Y(n_3824)
);

INVx8_ASAP7_75t_L g3825 ( 
.A(n_3557),
.Y(n_3825)
);

NOR2xp33_ASAP7_75t_L g3826 ( 
.A(n_3595),
.B(n_2197),
.Y(n_3826)
);

AND2x4_ASAP7_75t_L g3827 ( 
.A(n_3469),
.B(n_3018),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3399),
.A2(n_861),
.B1(n_1041),
.B2(n_1032),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_SL g3829 ( 
.A(n_3289),
.B(n_3050),
.Y(n_3829)
);

BUFx5_ASAP7_75t_L g3830 ( 
.A(n_3552),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3485),
.Y(n_3831)
);

INVx3_ASAP7_75t_L g3832 ( 
.A(n_3491),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3313),
.B(n_3093),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_SL g3834 ( 
.A(n_3539),
.B(n_3050),
.Y(n_3834)
);

INVx8_ASAP7_75t_L g3835 ( 
.A(n_3557),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3315),
.B(n_3097),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3487),
.Y(n_3837)
);

HB1xp67_ASAP7_75t_L g3838 ( 
.A(n_3288),
.Y(n_3838)
);

INVxp67_ASAP7_75t_L g3839 ( 
.A(n_3577),
.Y(n_3839)
);

INVx2_ASAP7_75t_SL g3840 ( 
.A(n_3562),
.Y(n_3840)
);

BUFx12f_ASAP7_75t_L g3841 ( 
.A(n_3483),
.Y(n_3841)
);

NOR2xp33_ASAP7_75t_L g3842 ( 
.A(n_3595),
.B(n_2197),
.Y(n_3842)
);

AOI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3399),
.A2(n_1003),
.B1(n_887),
.B2(n_969),
.Y(n_3843)
);

INVx8_ASAP7_75t_L g3844 ( 
.A(n_3557),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3317),
.B(n_3097),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3318),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3319),
.B(n_3099),
.Y(n_3847)
);

OAI22xp5_ASAP7_75t_L g3848 ( 
.A1(n_3546),
.A2(n_3050),
.B1(n_2946),
.B2(n_2991),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3323),
.B(n_3099),
.Y(n_3849)
);

NOR2xp33_ASAP7_75t_L g3850 ( 
.A(n_3410),
.B(n_2199),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3310),
.B(n_2946),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3581),
.B(n_2325),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3463),
.B(n_2199),
.Y(n_3853)
);

AOI22xp33_ASAP7_75t_L g3854 ( 
.A1(n_3399),
.A2(n_1003),
.B1(n_887),
.B2(n_969),
.Y(n_3854)
);

BUFx3_ASAP7_75t_L g3855 ( 
.A(n_3373),
.Y(n_3855)
);

BUFx12f_ASAP7_75t_L g3856 ( 
.A(n_3419),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3512),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3283),
.B(n_2946),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_L g3859 ( 
.A(n_3501),
.B(n_2207),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3324),
.B(n_3024),
.Y(n_3860)
);

NOR2xp33_ASAP7_75t_L g3861 ( 
.A(n_3507),
.B(n_2325),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3328),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3329),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3605),
.B(n_3034),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3428),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_3285),
.B(n_3050),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3286),
.B(n_2556),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3520),
.Y(n_3868)
);

INVx2_ASAP7_75t_SL g3869 ( 
.A(n_3301),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3432),
.Y(n_3870)
);

OAI22xp5_ASAP7_75t_L g3871 ( 
.A1(n_3507),
.A2(n_2991),
.B1(n_3086),
.B2(n_2969),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3529),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3613),
.B(n_3060),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3594),
.B(n_3060),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3260),
.B(n_2333),
.Y(n_3875)
);

INVx3_ASAP7_75t_L g3876 ( 
.A(n_3570),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3532),
.B(n_3078),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_3532),
.B(n_2333),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3434),
.Y(n_3879)
);

NOR2xp33_ASAP7_75t_L g3880 ( 
.A(n_3535),
.B(n_3540),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3260),
.B(n_2333),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3535),
.B(n_3170),
.Y(n_3882)
);

NOR3xp33_ASAP7_75t_L g3883 ( 
.A(n_3354),
.B(n_1994),
.C(n_2301),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3267),
.A2(n_3230),
.B(n_3227),
.Y(n_3884)
);

AND2x4_ASAP7_75t_SL g3885 ( 
.A(n_3321),
.B(n_3046),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_SL g3886 ( 
.A(n_3287),
.B(n_3115),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3400),
.B(n_3115),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_SL g3888 ( 
.A(n_3400),
.B(n_3115),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3436),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3440),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3441),
.Y(n_3891)
);

NOR2xp33_ASAP7_75t_SL g3892 ( 
.A(n_3263),
.B(n_2502),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3406),
.B(n_3506),
.Y(n_3893)
);

INVx4_ASAP7_75t_L g3894 ( 
.A(n_3307),
.Y(n_3894)
);

AOI22xp5_ASAP7_75t_L g3895 ( 
.A1(n_3508),
.A2(n_2512),
.B1(n_2301),
.B2(n_2502),
.Y(n_3895)
);

OAI221xp5_ASAP7_75t_L g3896 ( 
.A1(n_3276),
.A2(n_2186),
.B1(n_2200),
.B2(n_2187),
.C(n_2177),
.Y(n_3896)
);

BUFx3_ASAP7_75t_L g3897 ( 
.A(n_3600),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_SL g3898 ( 
.A(n_3406),
.B(n_3414),
.Y(n_3898)
);

AOI22xp5_ASAP7_75t_L g3899 ( 
.A1(n_3508),
.A2(n_3551),
.B1(n_3249),
.B2(n_3305),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3414),
.B(n_3210),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_3234),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_3418),
.B(n_3115),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3418),
.B(n_3210),
.Y(n_3903)
);

AND2x4_ASAP7_75t_L g3904 ( 
.A(n_3563),
.B(n_3573),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3573),
.B(n_3046),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3454),
.B(n_3218),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_SL g3907 ( 
.A(n_3474),
.B(n_3115),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3474),
.B(n_2992),
.Y(n_3908)
);

NOR2xp33_ASAP7_75t_L g3909 ( 
.A(n_3235),
.B(n_2512),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3506),
.B(n_3238),
.Y(n_3910)
);

BUFx6f_ASAP7_75t_SL g3911 ( 
.A(n_3592),
.Y(n_3911)
);

INVx2_ASAP7_75t_L g3912 ( 
.A(n_3237),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3239),
.B(n_2992),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3599),
.B(n_1946),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3241),
.B(n_2994),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_SL g3916 ( 
.A(n_3533),
.B(n_3267),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3243),
.B(n_2994),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_SL g3918 ( 
.A(n_3326),
.B(n_3343),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3244),
.B(n_2996),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3245),
.B(n_2996),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3250),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3445),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3252),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3447),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3255),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3256),
.B(n_2999),
.Y(n_3926)
);

NOR2xp33_ASAP7_75t_L g3927 ( 
.A(n_3258),
.B(n_2498),
.Y(n_3927)
);

INVx2_ASAP7_75t_SL g3928 ( 
.A(n_3364),
.Y(n_3928)
);

INVx3_ASAP7_75t_L g3929 ( 
.A(n_3307),
.Y(n_3929)
);

AOI22xp5_ASAP7_75t_L g3930 ( 
.A1(n_3551),
.A2(n_2505),
.B1(n_1875),
.B2(n_1874),
.Y(n_3930)
);

OAI22xp33_ASAP7_75t_L g3931 ( 
.A1(n_3305),
.A2(n_2408),
.B1(n_1086),
.B2(n_1082),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3266),
.B(n_2999),
.Y(n_3932)
);

NAND3xp33_ASAP7_75t_L g3933 ( 
.A(n_3582),
.B(n_2097),
.C(n_2505),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3269),
.B(n_3015),
.Y(n_3934)
);

INVxp33_ASAP7_75t_L g3935 ( 
.A(n_3314),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3270),
.B(n_3015),
.Y(n_3936)
);

INVx3_ASAP7_75t_L g3937 ( 
.A(n_3307),
.Y(n_3937)
);

NOR3xp33_ASAP7_75t_L g3938 ( 
.A(n_3462),
.B(n_2104),
.C(n_2038),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3450),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3451),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3271),
.B(n_3020),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3277),
.B(n_2561),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3399),
.A2(n_1003),
.B1(n_887),
.B2(n_969),
.Y(n_3943)
);

CKINVDCx5p33_ASAP7_75t_R g3944 ( 
.A(n_3511),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3278),
.B(n_2561),
.Y(n_3945)
);

OR2x2_ASAP7_75t_L g3946 ( 
.A(n_3339),
.B(n_2109),
.Y(n_3946)
);

NOR2xp33_ASAP7_75t_L g3947 ( 
.A(n_3279),
.B(n_3280),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3617),
.Y(n_3948)
);

A2O1A1Ixp33_ASAP7_75t_L g3949 ( 
.A1(n_3682),
.A2(n_3446),
.B(n_3282),
.C(n_3281),
.Y(n_3949)
);

AOI22xp5_ASAP7_75t_L g3950 ( 
.A1(n_3655),
.A2(n_2364),
.B1(n_2368),
.B2(n_2355),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3655),
.B(n_2578),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3697),
.B(n_3523),
.Y(n_3952)
);

BUFx6f_ASAP7_75t_L g3953 ( 
.A(n_3633),
.Y(n_3953)
);

NOR2x1p5_ASAP7_75t_L g3954 ( 
.A(n_3933),
.B(n_2418),
.Y(n_3954)
);

HB1xp67_ASAP7_75t_L g3955 ( 
.A(n_3638),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3697),
.B(n_3523),
.Y(n_3956)
);

BUFx6f_ASAP7_75t_L g3957 ( 
.A(n_3633),
.Y(n_3957)
);

HB1xp67_ASAP7_75t_L g3958 ( 
.A(n_3736),
.Y(n_3958)
);

NOR2xp67_ASAP7_75t_L g3959 ( 
.A(n_3796),
.B(n_3712),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3695),
.B(n_3785),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3711),
.A2(n_3248),
.B1(n_3233),
.B2(n_2564),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3626),
.Y(n_3962)
);

BUFx3_ASAP7_75t_L g3963 ( 
.A(n_3637),
.Y(n_3963)
);

AND2x4_ASAP7_75t_L g3964 ( 
.A(n_3904),
.B(n_3504),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3893),
.B(n_3552),
.Y(n_3965)
);

AOI22xp33_ASAP7_75t_L g3966 ( 
.A1(n_3711),
.A2(n_2564),
.B1(n_3552),
.B2(n_3565),
.Y(n_3966)
);

AOI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3645),
.A2(n_2368),
.B1(n_2370),
.B2(n_2364),
.Y(n_3967)
);

INVx4_ASAP7_75t_L g3968 ( 
.A(n_3633),
.Y(n_3968)
);

AOI22xp5_ASAP7_75t_L g3969 ( 
.A1(n_3645),
.A2(n_2372),
.B1(n_2388),
.B2(n_2370),
.Y(n_3969)
);

HB1xp67_ASAP7_75t_L g3970 ( 
.A(n_3736),
.Y(n_3970)
);

AND2x6_ASAP7_75t_SL g3971 ( 
.A(n_3859),
.B(n_3261),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3627),
.B(n_3552),
.Y(n_3972)
);

CKINVDCx20_ASAP7_75t_R g3973 ( 
.A(n_3855),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3901),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3634),
.Y(n_3975)
);

NOR2xp33_ASAP7_75t_R g3976 ( 
.A(n_3791),
.B(n_2372),
.Y(n_3976)
);

BUFx6f_ASAP7_75t_L g3977 ( 
.A(n_3633),
.Y(n_3977)
);

BUFx6f_ASAP7_75t_L g3978 ( 
.A(n_3803),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_3912),
.Y(n_3979)
);

O2A1O1Ixp33_ASAP7_75t_L g3980 ( 
.A1(n_3721),
.A2(n_2142),
.B(n_2143),
.C(n_2128),
.Y(n_3980)
);

OAI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3895),
.A2(n_3521),
.B1(n_3614),
.B2(n_3511),
.Y(n_3981)
);

NOR2xp33_ASAP7_75t_L g3982 ( 
.A(n_3946),
.B(n_2394),
.Y(n_3982)
);

BUFx3_ASAP7_75t_L g3983 ( 
.A(n_3765),
.Y(n_3983)
);

NOR2xp33_ASAP7_75t_L g3984 ( 
.A(n_3819),
.B(n_2464),
.Y(n_3984)
);

AND2x4_ASAP7_75t_L g3985 ( 
.A(n_3904),
.B(n_3505),
.Y(n_3985)
);

AND3x1_ASAP7_75t_SL g3986 ( 
.A(n_3896),
.B(n_789),
.C(n_764),
.Y(n_3986)
);

INVx3_ASAP7_75t_L g3987 ( 
.A(n_3702),
.Y(n_3987)
);

AOI22xp5_ASAP7_75t_L g3988 ( 
.A1(n_3853),
.A2(n_2470),
.B1(n_2464),
.B2(n_3350),
.Y(n_3988)
);

NOR2x1p5_ASAP7_75t_L g3989 ( 
.A(n_3856),
.B(n_2460),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3701),
.Y(n_3990)
);

BUFx6f_ASAP7_75t_L g3991 ( 
.A(n_3803),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3643),
.B(n_3452),
.Y(n_3992)
);

OAI22xp5_ASAP7_75t_SL g3993 ( 
.A1(n_3700),
.A2(n_2595),
.B1(n_2602),
.B2(n_2606),
.Y(n_3993)
);

INVx4_ASAP7_75t_L g3994 ( 
.A(n_3803),
.Y(n_3994)
);

BUFx6f_ASAP7_75t_L g3995 ( 
.A(n_3803),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3628),
.B(n_3624),
.Y(n_3996)
);

OAI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_3658),
.A2(n_3446),
.B(n_3232),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3644),
.B(n_3552),
.Y(n_3998)
);

OAI21xp33_ASAP7_75t_L g3999 ( 
.A1(n_3640),
.A2(n_2465),
.B(n_2461),
.Y(n_3999)
);

AOI22xp5_ASAP7_75t_L g4000 ( 
.A1(n_3853),
.A2(n_2470),
.B1(n_3385),
.B2(n_3521),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3650),
.B(n_3453),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3720),
.Y(n_4002)
);

NOR2xp33_ASAP7_75t_SL g4003 ( 
.A(n_3931),
.B(n_3614),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3652),
.B(n_3459),
.Y(n_4004)
);

HB1xp67_ASAP7_75t_L g4005 ( 
.A(n_3838),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3921),
.Y(n_4006)
);

BUFx6f_ASAP7_75t_L g4007 ( 
.A(n_3705),
.Y(n_4007)
);

INVx2_ASAP7_75t_SL g4008 ( 
.A(n_3647),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3731),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3667),
.B(n_2343),
.Y(n_4010)
);

AND3x2_ASAP7_75t_SL g4011 ( 
.A(n_3708),
.B(n_3054),
.C(n_2954),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3923),
.Y(n_4012)
);

AOI22xp33_ASAP7_75t_L g4013 ( 
.A1(n_3698),
.A2(n_2564),
.B1(n_3054),
.B2(n_2954),
.Y(n_4013)
);

INVx2_ASAP7_75t_L g4014 ( 
.A(n_3925),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3641),
.B(n_3460),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3733),
.Y(n_4016)
);

BUFx6f_ASAP7_75t_L g4017 ( 
.A(n_3705),
.Y(n_4017)
);

INVx2_ASAP7_75t_SL g4018 ( 
.A(n_3885),
.Y(n_4018)
);

INVx5_ASAP7_75t_L g4019 ( 
.A(n_3705),
.Y(n_4019)
);

INVx2_ASAP7_75t_SL g4020 ( 
.A(n_3623),
.Y(n_4020)
);

HB1xp67_ASAP7_75t_L g4021 ( 
.A(n_3678),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3641),
.B(n_3465),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3737),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_SL g4024 ( 
.A(n_3620),
.B(n_2461),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3741),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_3722),
.B(n_3468),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_SL g4027 ( 
.A(n_3732),
.B(n_2465),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3744),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3753),
.Y(n_4029)
);

BUFx2_ASAP7_75t_L g4030 ( 
.A(n_3772),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3722),
.B(n_3470),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3880),
.B(n_3476),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3880),
.B(n_3479),
.Y(n_4033)
);

BUFx6f_ASAP7_75t_L g4034 ( 
.A(n_3705),
.Y(n_4034)
);

AND2x4_ASAP7_75t_L g4035 ( 
.A(n_3746),
.B(n_3905),
.Y(n_4035)
);

BUFx6f_ASAP7_75t_L g4036 ( 
.A(n_3797),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_3911),
.Y(n_4037)
);

INVx2_ASAP7_75t_SL g4038 ( 
.A(n_3629),
.Y(n_4038)
);

NAND2x1p5_ASAP7_75t_L g4039 ( 
.A(n_3621),
.B(n_3579),
.Y(n_4039)
);

AND2x2_ASAP7_75t_SL g4040 ( 
.A(n_3673),
.B(n_3899),
.Y(n_4040)
);

INVx6_ASAP7_75t_L g4041 ( 
.A(n_3841),
.Y(n_4041)
);

AND2x6_ASAP7_75t_SL g4042 ( 
.A(n_3909),
.B(n_2612),
.Y(n_4042)
);

AOI22xp33_ASAP7_75t_SL g4043 ( 
.A1(n_3661),
.A2(n_2648),
.B1(n_2674),
.B2(n_2619),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_3850),
.B(n_2479),
.Y(n_4044)
);

NOR2x1p5_ASAP7_75t_L g4045 ( 
.A(n_3761),
.B(n_2479),
.Y(n_4045)
);

OR2x6_ASAP7_75t_L g4046 ( 
.A(n_3825),
.B(n_2797),
.Y(n_4046)
);

INVx3_ASAP7_75t_L g4047 ( 
.A(n_3702),
.Y(n_4047)
);

INVx5_ASAP7_75t_L g4048 ( 
.A(n_3797),
.Y(n_4048)
);

CKINVDCx5p33_ASAP7_75t_R g4049 ( 
.A(n_3944),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3760),
.Y(n_4050)
);

AND2x6_ASAP7_75t_L g4051 ( 
.A(n_3621),
.B(n_3480),
.Y(n_4051)
);

AOI22xp5_ASAP7_75t_L g4052 ( 
.A1(n_3914),
.A2(n_2539),
.B1(n_2562),
.B2(n_2532),
.Y(n_4052)
);

AND2x6_ASAP7_75t_SL g4053 ( 
.A(n_3909),
.B(n_2619),
.Y(n_4053)
);

OAI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3755),
.A2(n_3486),
.B1(n_3489),
.B2(n_3482),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3762),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3692),
.B(n_3492),
.Y(n_4056)
);

INVx4_ASAP7_75t_L g4057 ( 
.A(n_3797),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3766),
.Y(n_4058)
);

INVx1_ASAP7_75t_SL g4059 ( 
.A(n_3743),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_SL g4060 ( 
.A(n_3931),
.B(n_2585),
.Y(n_4060)
);

INVx1_ASAP7_75t_SL g4061 ( 
.A(n_3806),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_SL g4062 ( 
.A(n_3672),
.B(n_2586),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3783),
.Y(n_4063)
);

INVxp67_ASAP7_75t_L g4064 ( 
.A(n_3817),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3713),
.B(n_3494),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_L g4066 ( 
.A(n_3653),
.B(n_2344),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3792),
.Y(n_4067)
);

AND2x6_ASAP7_75t_SL g4068 ( 
.A(n_3631),
.B(n_2674),
.Y(n_4068)
);

NAND2x1p5_ASAP7_75t_L g4069 ( 
.A(n_3669),
.B(n_3579),
.Y(n_4069)
);

BUFx2_ASAP7_75t_L g4070 ( 
.A(n_3875),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3794),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3795),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3800),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_3694),
.B(n_3699),
.Y(n_4074)
);

AOI21xp5_ASAP7_75t_L g4075 ( 
.A1(n_3916),
.A2(n_3502),
.B(n_3484),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3684),
.B(n_3495),
.Y(n_4076)
);

INVx4_ASAP7_75t_L g4077 ( 
.A(n_3797),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3804),
.Y(n_4078)
);

INVx5_ASAP7_75t_L g4079 ( 
.A(n_3822),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3846),
.Y(n_4080)
);

INVxp67_ASAP7_75t_L g4081 ( 
.A(n_3631),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_3862),
.Y(n_4082)
);

NAND2xp33_ASAP7_75t_L g4083 ( 
.A(n_3938),
.B(n_2797),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3863),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3685),
.B(n_3496),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3898),
.B(n_3500),
.Y(n_4086)
);

NOR3xp33_ASAP7_75t_SL g4087 ( 
.A(n_3660),
.B(n_2586),
.C(n_2361),
.Y(n_4087)
);

AND2x4_ASAP7_75t_L g4088 ( 
.A(n_3738),
.B(n_3510),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_3898),
.B(n_3591),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_SL g4090 ( 
.A(n_3672),
.B(n_3662),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3910),
.B(n_3593),
.Y(n_4091)
);

INVx2_ASAP7_75t_SL g4092 ( 
.A(n_3717),
.Y(n_4092)
);

BUFx3_ASAP7_75t_L g4093 ( 
.A(n_3786),
.Y(n_4093)
);

OAI21xp5_ASAP7_75t_L g4094 ( 
.A1(n_3658),
.A2(n_3327),
.B(n_3574),
.Y(n_4094)
);

CKINVDCx5p33_ASAP7_75t_R g4095 ( 
.A(n_3897),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3808),
.B(n_3513),
.Y(n_4096)
);

AND2x4_ASAP7_75t_L g4097 ( 
.A(n_3738),
.B(n_3514),
.Y(n_4097)
);

AOI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3861),
.A2(n_2682),
.B1(n_3054),
.B2(n_2346),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_SL g4099 ( 
.A(n_3826),
.B(n_3515),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_3865),
.Y(n_4100)
);

BUFx6f_ASAP7_75t_L g4101 ( 
.A(n_3822),
.Y(n_4101)
);

HB1xp67_ASAP7_75t_L g4102 ( 
.A(n_3771),
.Y(n_4102)
);

OAI22xp5_ASAP7_75t_SL g4103 ( 
.A1(n_3755),
.A2(n_2682),
.B1(n_3412),
.B2(n_3322),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_3870),
.Y(n_4104)
);

BUFx6f_ASAP7_75t_L g4105 ( 
.A(n_3822),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3879),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3618),
.B(n_3615),
.Y(n_4107)
);

BUFx3_ASAP7_75t_L g4108 ( 
.A(n_3840),
.Y(n_4108)
);

BUFx12f_ASAP7_75t_L g4109 ( 
.A(n_3928),
.Y(n_4109)
);

INVxp67_ASAP7_75t_SL g4110 ( 
.A(n_3740),
.Y(n_4110)
);

BUFx6f_ASAP7_75t_L g4111 ( 
.A(n_3822),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3889),
.Y(n_4112)
);

AOI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_3916),
.A2(n_3502),
.B(n_3484),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_3618),
.B(n_3580),
.Y(n_4114)
);

INVx3_ASAP7_75t_L g4115 ( 
.A(n_3702),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3890),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3891),
.Y(n_4117)
);

AOI21xp33_ASAP7_75t_L g4118 ( 
.A1(n_3625),
.A2(n_3327),
.B(n_3574),
.Y(n_4118)
);

NAND2x1p5_ASAP7_75t_L g4119 ( 
.A(n_3669),
.B(n_3579),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3826),
.B(n_3518),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3654),
.B(n_3588),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3657),
.B(n_3596),
.Y(n_4122)
);

INVx4_ASAP7_75t_L g4123 ( 
.A(n_3825),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3842),
.B(n_3519),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3659),
.B(n_3602),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3922),
.Y(n_4126)
);

BUFx8_ASAP7_75t_L g4127 ( 
.A(n_3942),
.Y(n_4127)
);

INVx2_ASAP7_75t_SL g4128 ( 
.A(n_3639),
.Y(n_4128)
);

BUFx12f_ASAP7_75t_L g4129 ( 
.A(n_3649),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3924),
.Y(n_4130)
);

INVx2_ASAP7_75t_SL g4131 ( 
.A(n_3729),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3939),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3630),
.B(n_3606),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_3869),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_3940),
.Y(n_4135)
);

NOR2xp67_ASAP7_75t_L g4136 ( 
.A(n_3814),
.B(n_2363),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3635),
.B(n_3538),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3947),
.Y(n_4138)
);

OR2x6_ASAP7_75t_L g4139 ( 
.A(n_3835),
.B(n_3844),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3908),
.B(n_3543),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_SL g4141 ( 
.A(n_3759),
.B(n_3524),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_3852),
.B(n_3526),
.Y(n_4142)
);

NOR2xp33_ASAP7_75t_L g4143 ( 
.A(n_3935),
.B(n_2373),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3947),
.Y(n_4144)
);

AND2x4_ASAP7_75t_L g4145 ( 
.A(n_3739),
.B(n_3527),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3651),
.Y(n_4146)
);

BUFx6f_ASAP7_75t_L g4147 ( 
.A(n_3835),
.Y(n_4147)
);

BUFx6f_ASAP7_75t_L g4148 ( 
.A(n_3835),
.Y(n_4148)
);

AOI22xp33_ASAP7_75t_L g4149 ( 
.A1(n_3625),
.A2(n_2564),
.B1(n_3412),
.B2(n_2875),
.Y(n_4149)
);

BUFx4f_ASAP7_75t_L g4150 ( 
.A(n_3844),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_3656),
.Y(n_4151)
);

INVx2_ASAP7_75t_SL g4152 ( 
.A(n_3881),
.Y(n_4152)
);

NOR2xp33_ASAP7_75t_L g4153 ( 
.A(n_3719),
.B(n_2373),
.Y(n_4153)
);

HB1xp67_ASAP7_75t_L g4154 ( 
.A(n_3727),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_SL g4155 ( 
.A(n_3660),
.B(n_2374),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3663),
.Y(n_4156)
);

CKINVDCx5p33_ASAP7_75t_R g4157 ( 
.A(n_3636),
.Y(n_4157)
);

INVx2_ASAP7_75t_SL g4158 ( 
.A(n_3945),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3675),
.Y(n_4159)
);

AOI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_3878),
.A2(n_2374),
.B1(n_2391),
.B2(n_2377),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3677),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3679),
.Y(n_4162)
);

AOI22xp33_ASAP7_75t_L g4163 ( 
.A1(n_3748),
.A2(n_2564),
.B1(n_2875),
.B2(n_2807),
.Y(n_4163)
);

NAND3xp33_ASAP7_75t_SL g4164 ( 
.A(n_3883),
.B(n_2391),
.C(n_2377),
.Y(n_4164)
);

NOR2x1p5_ASAP7_75t_L g4165 ( 
.A(n_3671),
.B(n_3371),
.Y(n_4165)
);

AND2x4_ASAP7_75t_L g4166 ( 
.A(n_3739),
.B(n_3823),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3773),
.B(n_3604),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_3776),
.B(n_3607),
.Y(n_4168)
);

INVx2_ASAP7_75t_SL g4169 ( 
.A(n_3844),
.Y(n_4169)
);

INVx5_ASAP7_75t_L g4170 ( 
.A(n_3764),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3788),
.B(n_3710),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_3930),
.B(n_3374),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3665),
.B(n_3545),
.Y(n_4173)
);

INVx2_ASAP7_75t_SL g4174 ( 
.A(n_3823),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_SL g4175 ( 
.A(n_3688),
.B(n_2807),
.Y(n_4175)
);

BUFx3_ASAP7_75t_L g4176 ( 
.A(n_3728),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3687),
.Y(n_4177)
);

AOI22xp33_ASAP7_75t_L g4178 ( 
.A1(n_3748),
.A2(n_2875),
.B1(n_2807),
.B2(n_2117),
.Y(n_4178)
);

OAI21xp33_ASAP7_75t_L g4179 ( 
.A1(n_3802),
.A2(n_1037),
.B(n_1012),
.Y(n_4179)
);

INVx2_ASAP7_75t_SL g4180 ( 
.A(n_3827),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_3668),
.B(n_3567),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3703),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_3673),
.B(n_3568),
.Y(n_4183)
);

INVx2_ASAP7_75t_SL g4184 ( 
.A(n_3827),
.Y(n_4184)
);

BUFx4f_ASAP7_75t_L g4185 ( 
.A(n_3764),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3706),
.Y(n_4186)
);

AND2x4_ASAP7_75t_L g4187 ( 
.A(n_3751),
.B(n_3375),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_3696),
.B(n_3378),
.Y(n_4188)
);

AND3x1_ASAP7_75t_L g4189 ( 
.A(n_3883),
.B(n_1032),
.C(n_777),
.Y(n_4189)
);

OAI21xp5_ASAP7_75t_L g4190 ( 
.A1(n_3616),
.A2(n_3466),
.B(n_3142),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_3927),
.B(n_3381),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3716),
.Y(n_4192)
);

NOR2xp33_ASAP7_75t_L g4193 ( 
.A(n_3723),
.B(n_3724),
.Y(n_4193)
);

INVx3_ASAP7_75t_L g4194 ( 
.A(n_3894),
.Y(n_4194)
);

OAI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_3781),
.A2(n_3553),
.B1(n_3556),
.B2(n_3549),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3696),
.B(n_3387),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_3747),
.Y(n_4197)
);

AND2x6_ASAP7_75t_SL g4198 ( 
.A(n_3769),
.B(n_761),
.Y(n_4198)
);

BUFx2_ASAP7_75t_L g4199 ( 
.A(n_3839),
.Y(n_4199)
);

AOI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3790),
.A2(n_3938),
.B1(n_3789),
.B2(n_3782),
.Y(n_4200)
);

AOI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_3693),
.A2(n_2823),
.B1(n_3132),
.B2(n_3118),
.Y(n_4201)
);

AOI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_3734),
.A2(n_3132),
.B1(n_3118),
.B2(n_2969),
.Y(n_4202)
);

AOI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_3754),
.A2(n_3132),
.B1(n_2969),
.B2(n_3086),
.Y(n_4203)
);

INVx2_ASAP7_75t_SL g4204 ( 
.A(n_3769),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_3900),
.B(n_3564),
.Y(n_4205)
);

INVx3_ASAP7_75t_L g4206 ( 
.A(n_3894),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_3780),
.Y(n_4207)
);

INVx2_ASAP7_75t_L g4208 ( 
.A(n_3784),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_3809),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3903),
.B(n_3566),
.Y(n_4210)
);

INVx5_ASAP7_75t_L g4211 ( 
.A(n_3764),
.Y(n_4211)
);

CKINVDCx5p33_ASAP7_75t_R g4212 ( 
.A(n_3757),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3810),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_3906),
.B(n_3571),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3664),
.B(n_3572),
.Y(n_4215)
);

OR2x6_ASAP7_75t_L g4216 ( 
.A(n_3690),
.B(n_2921),
.Y(n_4216)
);

BUFx6f_ASAP7_75t_L g4217 ( 
.A(n_3929),
.Y(n_4217)
);

AND2x4_ASAP7_75t_L g4218 ( 
.A(n_3767),
.B(n_3390),
.Y(n_4218)
);

OAI22xp5_ASAP7_75t_SL g4219 ( 
.A1(n_3718),
.A2(n_734),
.B1(n_756),
.B2(n_683),
.Y(n_4219)
);

AOI22xp33_ASAP7_75t_L g4220 ( 
.A1(n_3718),
.A2(n_3648),
.B1(n_3666),
.B2(n_3632),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_SL g4221 ( 
.A(n_3674),
.B(n_3391),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3831),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_3683),
.B(n_3392),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_SL g4224 ( 
.A(n_3770),
.B(n_3393),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3837),
.Y(n_4225)
);

INVx2_ASAP7_75t_SL g4226 ( 
.A(n_3752),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_SL g4227 ( 
.A(n_3704),
.B(n_3396),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3857),
.Y(n_4228)
);

INVx1_ASAP7_75t_SL g4229 ( 
.A(n_3726),
.Y(n_4229)
);

HB1xp67_ASAP7_75t_L g4230 ( 
.A(n_3749),
.Y(n_4230)
);

O2A1O1Ixp33_ASAP7_75t_L g4231 ( 
.A1(n_3689),
.A2(n_934),
.B(n_963),
.C(n_921),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_3670),
.B(n_3401),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3868),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3872),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_3758),
.B(n_3560),
.Y(n_4235)
);

NOR2xp33_ASAP7_75t_L g4236 ( 
.A(n_3892),
.B(n_2991),
.Y(n_4236)
);

AOI21xp5_ASAP7_75t_L g4237 ( 
.A1(n_3884),
.A2(n_3768),
.B(n_3646),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3619),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_3622),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_3812),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3860),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_3750),
.B(n_3402),
.Y(n_4242)
);

AND2x4_ASAP7_75t_L g4243 ( 
.A(n_3811),
.B(n_3404),
.Y(n_4243)
);

INVx3_ASAP7_75t_L g4244 ( 
.A(n_3818),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3820),
.Y(n_4245)
);

NOR3xp33_ASAP7_75t_L g4246 ( 
.A(n_3763),
.B(n_934),
.C(n_921),
.Y(n_4246)
);

NAND2xp33_ASAP7_75t_SL g4247 ( 
.A(n_3691),
.B(n_3579),
.Y(n_4247)
);

INVxp67_ASAP7_75t_L g4248 ( 
.A(n_3775),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_3715),
.B(n_3561),
.Y(n_4249)
);

CKINVDCx5p33_ASAP7_75t_R g4250 ( 
.A(n_3775),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_3715),
.B(n_3575),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_3799),
.B(n_3405),
.Y(n_4252)
);

AOI22xp33_ASAP7_75t_L g4253 ( 
.A1(n_3680),
.A2(n_2117),
.B1(n_2031),
.B2(n_3132),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_3833),
.Y(n_4254)
);

AND2x4_ASAP7_75t_L g4255 ( 
.A(n_3811),
.B(n_3408),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_3836),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_3845),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_3730),
.B(n_3610),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_3847),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_3849),
.Y(n_4260)
);

BUFx4f_ASAP7_75t_L g4261 ( 
.A(n_3937),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_3793),
.B(n_3415),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_3735),
.B(n_3583),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3913),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_3787),
.B(n_3584),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_3915),
.Y(n_4266)
);

AOI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_3829),
.A2(n_3597),
.B(n_3585),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_3917),
.Y(n_4268)
);

AND2x6_ASAP7_75t_L g4269 ( 
.A(n_3818),
.B(n_3417),
.Y(n_4269)
);

AOI22xp5_ASAP7_75t_L g4270 ( 
.A1(n_3742),
.A2(n_3132),
.B1(n_3149),
.B2(n_2921),
.Y(n_4270)
);

INVxp67_ASAP7_75t_SL g4271 ( 
.A(n_3801),
.Y(n_4271)
);

NOR2xp33_ASAP7_75t_L g4272 ( 
.A(n_3793),
.B(n_3149),
.Y(n_4272)
);

BUFx6f_ASAP7_75t_L g4273 ( 
.A(n_3937),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3919),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_3920),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_3709),
.B(n_3420),
.Y(n_4276)
);

OAI21xp5_ASAP7_75t_L g4277 ( 
.A1(n_3616),
.A2(n_3142),
.B(n_3333),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3948),
.Y(n_4278)
);

AOI22xp33_ASAP7_75t_L g4279 ( 
.A1(n_4219),
.A2(n_4040),
.B1(n_4003),
.B2(n_4193),
.Y(n_4279)
);

INVx3_ASAP7_75t_SL g4280 ( 
.A(n_4049),
.Y(n_4280)
);

INVx3_ASAP7_75t_L g4281 ( 
.A(n_4217),
.Y(n_4281)
);

OR2x4_ASAP7_75t_L g4282 ( 
.A(n_4164),
.B(n_3798),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3962),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_3952),
.B(n_3676),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_3974),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_3979),
.Y(n_4286)
);

OAI22xp5_ASAP7_75t_L g4287 ( 
.A1(n_3961),
.A2(n_3781),
.B1(n_3843),
.B2(n_3828),
.Y(n_4287)
);

NOR2xp33_ASAP7_75t_L g4288 ( 
.A(n_4010),
.B(n_3864),
.Y(n_4288)
);

BUFx6f_ASAP7_75t_L g4289 ( 
.A(n_4129),
.Y(n_4289)
);

AND2x4_ASAP7_75t_L g4290 ( 
.A(n_4139),
.B(n_4243),
.Y(n_4290)
);

BUFx3_ASAP7_75t_L g4291 ( 
.A(n_3983),
.Y(n_4291)
);

AND2x2_ASAP7_75t_SL g4292 ( 
.A(n_4185),
.B(n_3828),
.Y(n_4292)
);

OAI221xp5_ASAP7_75t_L g4293 ( 
.A1(n_4003),
.A2(n_3943),
.B1(n_3854),
.B2(n_3843),
.C(n_3707),
.Y(n_4293)
);

INVxp67_ASAP7_75t_SL g4294 ( 
.A(n_4015),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3975),
.Y(n_4295)
);

BUFx3_ASAP7_75t_L g4296 ( 
.A(n_3973),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4006),
.Y(n_4297)
);

OAI221xp5_ASAP7_75t_L g4298 ( 
.A1(n_4179),
.A2(n_3943),
.B1(n_3854),
.B2(n_3681),
.C(n_3686),
.Y(n_4298)
);

INVx3_ASAP7_75t_L g4299 ( 
.A(n_4217),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4012),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3952),
.B(n_3787),
.Y(n_4301)
);

NOR2xp33_ASAP7_75t_R g4302 ( 
.A(n_4157),
.B(n_3830),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_3956),
.B(n_3830),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_3956),
.B(n_3830),
.Y(n_4304)
);

HB1xp67_ASAP7_75t_L g4305 ( 
.A(n_3958),
.Y(n_4305)
);

INVx4_ASAP7_75t_L g4306 ( 
.A(n_3953),
.Y(n_4306)
);

INVxp67_ASAP7_75t_L g4307 ( 
.A(n_3970),
.Y(n_4307)
);

INVxp67_ASAP7_75t_SL g4308 ( 
.A(n_4015),
.Y(n_4308)
);

NOR2xp33_ASAP7_75t_L g4309 ( 
.A(n_4176),
.B(n_3873),
.Y(n_4309)
);

OR2x6_ASAP7_75t_L g4310 ( 
.A(n_4216),
.B(n_3725),
.Y(n_4310)
);

CKINVDCx5p33_ASAP7_75t_R g4311 ( 
.A(n_4037),
.Y(n_4311)
);

BUFx10_ASAP7_75t_L g4312 ( 
.A(n_4041),
.Y(n_4312)
);

NOR2xp33_ASAP7_75t_L g4313 ( 
.A(n_4250),
.B(n_3874),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4074),
.B(n_3830),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4014),
.Y(n_4315)
);

CKINVDCx5p33_ASAP7_75t_R g4316 ( 
.A(n_4134),
.Y(n_4316)
);

INVxp67_ASAP7_75t_SL g4317 ( 
.A(n_4022),
.Y(n_4317)
);

NAND3xp33_ASAP7_75t_SL g4318 ( 
.A(n_3966),
.B(n_3686),
.C(n_3745),
.Y(n_4318)
);

AOI21xp5_ASAP7_75t_L g4319 ( 
.A1(n_3997),
.A2(n_3829),
.B(n_3834),
.Y(n_4319)
);

INVx3_ASAP7_75t_L g4320 ( 
.A(n_4217),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4058),
.Y(n_4321)
);

AND2x4_ASAP7_75t_L g4322 ( 
.A(n_4139),
.B(n_3886),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4204),
.B(n_4061),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4061),
.B(n_3830),
.Y(n_4324)
);

BUFx6f_ASAP7_75t_L g4325 ( 
.A(n_4147),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_4171),
.B(n_3926),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4171),
.B(n_3932),
.Y(n_4327)
);

NOR2xp33_ASAP7_75t_L g4328 ( 
.A(n_3982),
.B(n_3778),
.Y(n_4328)
);

OR2x6_ASAP7_75t_L g4329 ( 
.A(n_4216),
.B(n_4237),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_3960),
.B(n_3934),
.Y(n_4330)
);

INVx2_ASAP7_75t_SL g4331 ( 
.A(n_4108),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_3990),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4002),
.Y(n_4333)
);

INVx4_ASAP7_75t_L g4334 ( 
.A(n_3953),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3960),
.B(n_3936),
.Y(n_4335)
);

BUFx6f_ASAP7_75t_L g4336 ( 
.A(n_4147),
.Y(n_4336)
);

BUFx12f_ASAP7_75t_L g4337 ( 
.A(n_4041),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4032),
.B(n_3941),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_4032),
.B(n_3887),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4009),
.Y(n_4340)
);

BUFx6f_ASAP7_75t_L g4341 ( 
.A(n_4147),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4016),
.Y(n_4342)
);

AOI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4200),
.A2(n_3816),
.B1(n_3714),
.B2(n_3642),
.Y(n_4343)
);

INVx3_ASAP7_75t_L g4344 ( 
.A(n_4273),
.Y(n_4344)
);

INVxp67_ASAP7_75t_SL g4345 ( 
.A(n_4022),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4023),
.Y(n_4346)
);

AO21x2_ASAP7_75t_L g4347 ( 
.A1(n_4075),
.A2(n_3851),
.B(n_3815),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4067),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4072),
.Y(n_4349)
);

HB1xp67_ASAP7_75t_L g4350 ( 
.A(n_4005),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_SL g4351 ( 
.A(n_3959),
.B(n_3756),
.Y(n_4351)
);

BUFx2_ASAP7_75t_L g4352 ( 
.A(n_3955),
.Y(n_4352)
);

CKINVDCx20_ASAP7_75t_R g4353 ( 
.A(n_3976),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4033),
.B(n_3887),
.Y(n_4354)
);

NOR2xp33_ASAP7_75t_L g4355 ( 
.A(n_3984),
.B(n_734),
.Y(n_4355)
);

NOR3xp33_ASAP7_75t_SL g4356 ( 
.A(n_3999),
.B(n_845),
.C(n_844),
.Y(n_4356)
);

BUFx6f_ASAP7_75t_L g4357 ( 
.A(n_4148),
.Y(n_4357)
);

AND2x4_ASAP7_75t_L g4358 ( 
.A(n_4139),
.B(n_3886),
.Y(n_4358)
);

AND2x4_ASAP7_75t_L g4359 ( 
.A(n_4243),
.B(n_3821),
.Y(n_4359)
);

INVx2_ASAP7_75t_SL g4360 ( 
.A(n_4093),
.Y(n_4360)
);

INVx1_ASAP7_75t_SL g4361 ( 
.A(n_4199),
.Y(n_4361)
);

AOI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_4212),
.A2(n_3813),
.B1(n_3815),
.B2(n_3774),
.Y(n_4362)
);

INVx5_ASAP7_75t_L g4363 ( 
.A(n_4051),
.Y(n_4363)
);

INVxp67_ASAP7_75t_L g4364 ( 
.A(n_4138),
.Y(n_4364)
);

NOR3xp33_ASAP7_75t_SL g4365 ( 
.A(n_4060),
.B(n_849),
.C(n_847),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4080),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4025),
.Y(n_4367)
);

AND2x4_ASAP7_75t_L g4368 ( 
.A(n_4255),
.B(n_3821),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4028),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4082),
.Y(n_4370)
);

NOR2xp33_ASAP7_75t_L g4371 ( 
.A(n_3950),
.B(n_756),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_4033),
.B(n_3888),
.Y(n_4372)
);

OAI21xp5_ASAP7_75t_L g4373 ( 
.A1(n_3949),
.A2(n_3813),
.B(n_3867),
.Y(n_4373)
);

OR2x6_ASAP7_75t_L g4374 ( 
.A(n_4216),
.B(n_3824),
.Y(n_4374)
);

OR2x6_ASAP7_75t_L g4375 ( 
.A(n_4046),
.B(n_3824),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_3996),
.B(n_3888),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4100),
.Y(n_4377)
);

INVx3_ASAP7_75t_L g4378 ( 
.A(n_4273),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4029),
.Y(n_4379)
);

OR2x2_ASAP7_75t_L g4380 ( 
.A(n_4154),
.B(n_3877),
.Y(n_4380)
);

OAI221xp5_ASAP7_75t_L g4381 ( 
.A1(n_4027),
.A2(n_1031),
.B1(n_1045),
.B2(n_1002),
.C(n_963),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4104),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4106),
.Y(n_4383)
);

NOR2x1p5_ASAP7_75t_L g4384 ( 
.A(n_3987),
.B(n_3882),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4050),
.Y(n_4385)
);

NAND2x1p5_ASAP7_75t_L g4386 ( 
.A(n_4170),
.B(n_3902),
.Y(n_4386)
);

NAND2x1p5_ASAP7_75t_L g4387 ( 
.A(n_4170),
.B(n_3902),
.Y(n_4387)
);

INVxp67_ASAP7_75t_SL g4388 ( 
.A(n_4026),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4116),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_3996),
.B(n_3907),
.Y(n_4390)
);

BUFx6f_ASAP7_75t_L g4391 ( 
.A(n_4148),
.Y(n_4391)
);

AOI22xp33_ASAP7_75t_L g4392 ( 
.A1(n_4103),
.A2(n_1032),
.B1(n_1050),
.B2(n_1041),
.Y(n_4392)
);

BUFx6f_ASAP7_75t_L g4393 ( 
.A(n_4148),
.Y(n_4393)
);

NOR2xp33_ASAP7_75t_R g4394 ( 
.A(n_4095),
.B(n_3832),
.Y(n_4394)
);

AND3x1_ASAP7_75t_SL g4395 ( 
.A(n_3954),
.B(n_764),
.C(n_761),
.Y(n_4395)
);

BUFx3_ASAP7_75t_L g4396 ( 
.A(n_4109),
.Y(n_4396)
);

BUFx6f_ASAP7_75t_L g4397 ( 
.A(n_4150),
.Y(n_4397)
);

AND2x4_ASAP7_75t_L g4398 ( 
.A(n_4255),
.B(n_3858),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4096),
.B(n_4142),
.Y(n_4399)
);

INVx5_ASAP7_75t_L g4400 ( 
.A(n_4051),
.Y(n_4400)
);

AOI22xp5_ASAP7_75t_L g4401 ( 
.A1(n_4024),
.A2(n_853),
.B1(n_854),
.B2(n_851),
.Y(n_4401)
);

INVx5_ASAP7_75t_L g4402 ( 
.A(n_4051),
.Y(n_4402)
);

OR2x6_ASAP7_75t_L g4403 ( 
.A(n_4046),
.B(n_3965),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4055),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4271),
.B(n_3907),
.Y(n_4405)
);

OR2x6_ASAP7_75t_L g4406 ( 
.A(n_4046),
.B(n_3851),
.Y(n_4406)
);

INVx2_ASAP7_75t_SL g4407 ( 
.A(n_4020),
.Y(n_4407)
);

NOR3xp33_ASAP7_75t_SL g4408 ( 
.A(n_3981),
.B(n_856),
.C(n_855),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_4126),
.Y(n_4409)
);

INVxp67_ASAP7_75t_SL g4410 ( 
.A(n_4026),
.Y(n_4410)
);

AOI22xp5_ASAP7_75t_L g4411 ( 
.A1(n_3951),
.A2(n_859),
.B1(n_860),
.B2(n_858),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_SL g4412 ( 
.A(n_4081),
.B(n_3876),
.Y(n_4412)
);

BUFx6f_ASAP7_75t_L g4413 ( 
.A(n_4150),
.Y(n_4413)
);

INVx2_ASAP7_75t_L g4414 ( 
.A(n_4130),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4110),
.B(n_3805),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4135),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4264),
.B(n_3807),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4063),
.Y(n_4418)
);

NAND3xp33_ASAP7_75t_SL g4419 ( 
.A(n_3980),
.B(n_780),
.C(n_826),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4071),
.Y(n_4420)
);

NAND3xp33_ASAP7_75t_SL g4421 ( 
.A(n_3967),
.B(n_780),
.C(n_826),
.Y(n_4421)
);

BUFx2_ASAP7_75t_L g4422 ( 
.A(n_4035),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4073),
.Y(n_4423)
);

NOR2xp33_ASAP7_75t_L g4424 ( 
.A(n_3969),
.B(n_838),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4078),
.Y(n_4425)
);

INVx2_ASAP7_75t_L g4426 ( 
.A(n_4146),
.Y(n_4426)
);

BUFx6f_ASAP7_75t_L g4427 ( 
.A(n_3953),
.Y(n_4427)
);

INVx4_ASAP7_75t_L g4428 ( 
.A(n_3957),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_4151),
.Y(n_4429)
);

BUFx3_ASAP7_75t_L g4430 ( 
.A(n_4008),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4084),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4192),
.Y(n_4432)
);

AND2x2_ASAP7_75t_L g4433 ( 
.A(n_4030),
.B(n_3777),
.Y(n_4433)
);

AND2x2_ASAP7_75t_SL g4434 ( 
.A(n_4185),
.B(n_891),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_SL g4435 ( 
.A(n_4044),
.B(n_3876),
.Y(n_4435)
);

AND2x4_ASAP7_75t_L g4436 ( 
.A(n_3987),
.B(n_3858),
.Y(n_4436)
);

CKINVDCx5p33_ASAP7_75t_R g4437 ( 
.A(n_4127),
.Y(n_4437)
);

BUFx6f_ASAP7_75t_L g4438 ( 
.A(n_3957),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_4197),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4207),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4208),
.Y(n_4441)
);

BUFx2_ASAP7_75t_L g4442 ( 
.A(n_4166),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4209),
.Y(n_4443)
);

HB1xp67_ASAP7_75t_L g4444 ( 
.A(n_4102),
.Y(n_4444)
);

BUFx3_ASAP7_75t_L g4445 ( 
.A(n_4127),
.Y(n_4445)
);

HB1xp67_ASAP7_75t_L g4446 ( 
.A(n_4059),
.Y(n_4446)
);

BUFx6f_ASAP7_75t_L g4447 ( 
.A(n_3957),
.Y(n_4447)
);

BUFx3_ASAP7_75t_L g4448 ( 
.A(n_3963),
.Y(n_4448)
);

NOR3xp33_ASAP7_75t_SL g4449 ( 
.A(n_4062),
.B(n_4155),
.C(n_3993),
.Y(n_4449)
);

AND2x4_ASAP7_75t_L g4450 ( 
.A(n_4047),
.B(n_3866),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4112),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4266),
.B(n_3779),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4117),
.Y(n_4453)
);

INVx3_ASAP7_75t_L g4454 ( 
.A(n_4273),
.Y(n_4454)
);

NOR3xp33_ASAP7_75t_SL g4455 ( 
.A(n_4153),
.B(n_4066),
.C(n_4090),
.Y(n_4455)
);

INVx4_ASAP7_75t_L g4456 ( 
.A(n_3977),
.Y(n_4456)
);

BUFx3_ASAP7_75t_L g4457 ( 
.A(n_4018),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4268),
.B(n_3421),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4274),
.B(n_3423),
.Y(n_4459)
);

AOI22x1_ASAP7_75t_L g4460 ( 
.A1(n_4165),
.A2(n_890),
.B1(n_923),
.B2(n_874),
.Y(n_4460)
);

BUFx10_ASAP7_75t_L g4461 ( 
.A(n_3989),
.Y(n_4461)
);

AND2x4_ASAP7_75t_L g4462 ( 
.A(n_4047),
.B(n_3866),
.Y(n_4462)
);

BUFx6f_ASAP7_75t_L g4463 ( 
.A(n_3977),
.Y(n_4463)
);

BUFx6f_ASAP7_75t_L g4464 ( 
.A(n_3977),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4132),
.Y(n_4465)
);

NAND2x1p5_ASAP7_75t_L g4466 ( 
.A(n_4170),
.B(n_3834),
.Y(n_4466)
);

INVx5_ASAP7_75t_L g4467 ( 
.A(n_4051),
.Y(n_4467)
);

BUFx6f_ASAP7_75t_L g4468 ( 
.A(n_3978),
.Y(n_4468)
);

INVx1_ASAP7_75t_SL g4469 ( 
.A(n_4242),
.Y(n_4469)
);

BUFx2_ASAP7_75t_L g4470 ( 
.A(n_4070),
.Y(n_4470)
);

BUFx4f_ASAP7_75t_L g4471 ( 
.A(n_3978),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4275),
.B(n_3424),
.Y(n_4472)
);

NAND3xp33_ASAP7_75t_SL g4473 ( 
.A(n_4229),
.B(n_972),
.C(n_960),
.Y(n_4473)
);

AND2x4_ASAP7_75t_L g4474 ( 
.A(n_4115),
.B(n_3425),
.Y(n_4474)
);

INVx3_ASAP7_75t_L g4475 ( 
.A(n_4057),
.Y(n_4475)
);

BUFx4f_ASAP7_75t_L g4476 ( 
.A(n_3978),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_3965),
.B(n_3426),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4031),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4086),
.Y(n_4479)
);

AND2x4_ASAP7_75t_L g4480 ( 
.A(n_4115),
.B(n_3918),
.Y(n_4480)
);

INVx5_ASAP7_75t_L g4481 ( 
.A(n_4269),
.Y(n_4481)
);

INVx2_ASAP7_75t_SL g4482 ( 
.A(n_4038),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4001),
.B(n_3528),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_4001),
.B(n_3530),
.Y(n_4484)
);

AND2x4_ASAP7_75t_L g4485 ( 
.A(n_4123),
.B(n_3918),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_L g4486 ( 
.A(n_4004),
.B(n_3531),
.Y(n_4486)
);

OR2x6_ASAP7_75t_L g4487 ( 
.A(n_4113),
.B(n_3871),
.Y(n_4487)
);

INVx3_ASAP7_75t_L g4488 ( 
.A(n_4057),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4089),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4004),
.B(n_3105),
.Y(n_4490)
);

NOR2xp33_ASAP7_75t_R g4491 ( 
.A(n_4158),
.B(n_2921),
.Y(n_4491)
);

NOR2xp33_ASAP7_75t_R g4492 ( 
.A(n_4152),
.B(n_2921),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_L g4493 ( 
.A(n_3988),
.B(n_960),
.Y(n_4493)
);

BUFx6f_ASAP7_75t_L g4494 ( 
.A(n_3991),
.Y(n_4494)
);

BUFx12f_ASAP7_75t_L g4495 ( 
.A(n_4045),
.Y(n_4495)
);

INVx5_ASAP7_75t_L g4496 ( 
.A(n_4269),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4089),
.Y(n_4497)
);

NAND2x1p5_ASAP7_75t_L g4498 ( 
.A(n_4211),
.B(n_2780),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4056),
.B(n_3105),
.Y(n_4499)
);

BUFx3_ASAP7_75t_L g4500 ( 
.A(n_4092),
.Y(n_4500)
);

INVx5_ASAP7_75t_L g4501 ( 
.A(n_4269),
.Y(n_4501)
);

NOR3xp33_ASAP7_75t_SL g4502 ( 
.A(n_4143),
.B(n_875),
.C(n_873),
.Y(n_4502)
);

NOR2xp33_ASAP7_75t_L g4503 ( 
.A(n_4064),
.B(n_972),
.Y(n_4503)
);

OR2x6_ASAP7_75t_SL g4504 ( 
.A(n_4011),
.B(n_3972),
.Y(n_4504)
);

AND2x4_ASAP7_75t_L g4505 ( 
.A(n_4123),
.B(n_3294),
.Y(n_4505)
);

HB1xp67_ASAP7_75t_L g4506 ( 
.A(n_4230),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_4056),
.B(n_2896),
.Y(n_4507)
);

CKINVDCx8_ASAP7_75t_R g4508 ( 
.A(n_4068),
.Y(n_4508)
);

AND2x4_ASAP7_75t_L g4509 ( 
.A(n_4211),
.B(n_3294),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_4156),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4076),
.B(n_2896),
.Y(n_4511)
);

INVx1_ASAP7_75t_SL g4512 ( 
.A(n_4262),
.Y(n_4512)
);

INVx3_ASAP7_75t_L g4513 ( 
.A(n_4077),
.Y(n_4513)
);

INVx4_ASAP7_75t_L g4514 ( 
.A(n_3991),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_4076),
.B(n_2903),
.Y(n_4515)
);

INVx1_ASAP7_75t_SL g4516 ( 
.A(n_4188),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4159),
.Y(n_4517)
);

OR2x2_ASAP7_75t_SL g4518 ( 
.A(n_4021),
.B(n_4198),
.Y(n_4518)
);

NOR3xp33_ASAP7_75t_SL g4519 ( 
.A(n_4172),
.B(n_880),
.C(n_878),
.Y(n_4519)
);

BUFx10_ASAP7_75t_L g4520 ( 
.A(n_4236),
.Y(n_4520)
);

AOI22xp5_ASAP7_75t_L g4521 ( 
.A1(n_4098),
.A2(n_883),
.B1(n_884),
.B2(n_881),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_4161),
.Y(n_4522)
);

INVx4_ASAP7_75t_L g4523 ( 
.A(n_3991),
.Y(n_4523)
);

INVx3_ASAP7_75t_L g4524 ( 
.A(n_4077),
.Y(n_4524)
);

OR2x6_ASAP7_75t_L g4525 ( 
.A(n_3997),
.B(n_4249),
.Y(n_4525)
);

OR2x2_ASAP7_75t_SL g4526 ( 
.A(n_4241),
.B(n_891),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4162),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4085),
.B(n_2903),
.Y(n_4528)
);

BUFx2_ASAP7_75t_L g4529 ( 
.A(n_4007),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_4177),
.Y(n_4530)
);

INVx3_ASAP7_75t_L g4531 ( 
.A(n_3995),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_4182),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4186),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_4229),
.B(n_3848),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4213),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4222),
.Y(n_4536)
);

BUFx6f_ASAP7_75t_L g4537 ( 
.A(n_3995),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4225),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4085),
.B(n_2912),
.Y(n_4539)
);

INVx3_ASAP7_75t_L g4540 ( 
.A(n_3995),
.Y(n_4540)
);

BUFx10_ASAP7_75t_L g4541 ( 
.A(n_4131),
.Y(n_4541)
);

NOR2xp33_ASAP7_75t_R g4542 ( 
.A(n_4174),
.B(n_3132),
.Y(n_4542)
);

AND2x4_ASAP7_75t_L g4543 ( 
.A(n_4211),
.B(n_3294),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4121),
.B(n_4122),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_4121),
.B(n_2912),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4228),
.Y(n_4546)
);

INVxp67_ASAP7_75t_L g4547 ( 
.A(n_4144),
.Y(n_4547)
);

BUFx6f_ASAP7_75t_L g4548 ( 
.A(n_4007),
.Y(n_4548)
);

AND2x4_ASAP7_75t_L g4549 ( 
.A(n_3964),
.B(n_3395),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4122),
.B(n_2914),
.Y(n_4550)
);

INVx2_ASAP7_75t_SL g4551 ( 
.A(n_4128),
.Y(n_4551)
);

BUFx6f_ASAP7_75t_L g4552 ( 
.A(n_4007),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4233),
.Y(n_4553)
);

OAI21xp5_ASAP7_75t_L g4554 ( 
.A1(n_4220),
.A2(n_2897),
.B(n_3585),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4234),
.Y(n_4555)
);

AND2x6_ASAP7_75t_SL g4556 ( 
.A(n_4272),
.B(n_768),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_L g4557 ( 
.A(n_4125),
.B(n_2914),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4238),
.Y(n_4558)
);

INVx5_ASAP7_75t_L g4559 ( 
.A(n_3968),
.Y(n_4559)
);

BUFx6f_ASAP7_75t_L g4560 ( 
.A(n_4017),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4125),
.B(n_2915),
.Y(n_4561)
);

OAI22xp5_ASAP7_75t_L g4562 ( 
.A1(n_4189),
.A2(n_1012),
.B1(n_1037),
.B2(n_979),
.Y(n_4562)
);

AOI22xp33_ASAP7_75t_L g4563 ( 
.A1(n_4149),
.A2(n_1041),
.B1(n_1050),
.B2(n_949),
.Y(n_4563)
);

O2A1O1Ixp33_ASAP7_75t_L g4564 ( 
.A1(n_4191),
.A2(n_1002),
.B(n_1045),
.C(n_1031),
.Y(n_4564)
);

BUFx4f_ASAP7_75t_SL g4565 ( 
.A(n_4169),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4239),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4235),
.B(n_2915),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4265),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4265),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4249),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_3972),
.B(n_2917),
.Y(n_4571)
);

OR2x6_ASAP7_75t_L g4572 ( 
.A(n_4251),
.B(n_4267),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4251),
.Y(n_4573)
);

NAND2x1p5_ASAP7_75t_L g4574 ( 
.A(n_3968),
.B(n_2780),
.Y(n_4574)
);

BUFx3_ASAP7_75t_L g4575 ( 
.A(n_4261),
.Y(n_4575)
);

OAI22xp5_ASAP7_75t_L g4576 ( 
.A1(n_4189),
.A2(n_1071),
.B1(n_1082),
.B2(n_979),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4183),
.B(n_2924),
.Y(n_4577)
);

BUFx2_ASAP7_75t_L g4578 ( 
.A(n_4017),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_3964),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4183),
.Y(n_4580)
);

BUFx6f_ASAP7_75t_L g4581 ( 
.A(n_4017),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_3985),
.Y(n_4582)
);

HB1xp67_ASAP7_75t_L g4583 ( 
.A(n_4196),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_3985),
.Y(n_4584)
);

NOR2xp33_ASAP7_75t_L g4585 ( 
.A(n_4248),
.B(n_1071),
.Y(n_4585)
);

INVxp67_ASAP7_75t_L g4586 ( 
.A(n_4099),
.Y(n_4586)
);

NOR2xp33_ASAP7_75t_R g4587 ( 
.A(n_4180),
.B(n_2898),
.Y(n_4587)
);

INVx1_ASAP7_75t_SL g4588 ( 
.A(n_4120),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4218),
.Y(n_4589)
);

NOR2xp67_ASAP7_75t_L g4590 ( 
.A(n_4226),
.B(n_2787),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4173),
.B(n_2924),
.Y(n_4591)
);

INVx3_ASAP7_75t_L g4592 ( 
.A(n_4034),
.Y(n_4592)
);

CKINVDCx16_ASAP7_75t_R g4593 ( 
.A(n_4052),
.Y(n_4593)
);

BUFx6f_ASAP7_75t_L g4594 ( 
.A(n_4034),
.Y(n_4594)
);

INVx2_ASAP7_75t_SL g4595 ( 
.A(n_4034),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_4259),
.Y(n_4596)
);

NAND2xp5_ASAP7_75t_L g4597 ( 
.A(n_4173),
.B(n_4181),
.Y(n_4597)
);

NAND3xp33_ASAP7_75t_SL g4598 ( 
.A(n_4231),
.B(n_1084),
.C(n_1086),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4276),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4221),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4065),
.B(n_1511),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4223),
.Y(n_4602)
);

BUFx10_ASAP7_75t_L g4603 ( 
.A(n_4042),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4227),
.Y(n_4604)
);

NOR2xp33_ASAP7_75t_L g4605 ( 
.A(n_4000),
.B(n_3971),
.Y(n_4605)
);

AO22x1_ASAP7_75t_L g4606 ( 
.A1(n_4088),
.A2(n_4097),
.B1(n_4145),
.B2(n_4246),
.Y(n_4606)
);

INVx4_ASAP7_75t_L g4607 ( 
.A(n_4019),
.Y(n_4607)
);

INVx2_ASAP7_75t_L g4608 ( 
.A(n_4260),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4184),
.B(n_1514),
.Y(n_4609)
);

CKINVDCx5p33_ASAP7_75t_R g4610 ( 
.A(n_4087),
.Y(n_4610)
);

INVx1_ASAP7_75t_SL g4611 ( 
.A(n_4124),
.Y(n_4611)
);

INVx2_ASAP7_75t_L g4612 ( 
.A(n_4187),
.Y(n_4612)
);

AOI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4175),
.A2(n_901),
.B1(n_902),
.B2(n_899),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4181),
.B(n_2929),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4232),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4240),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4258),
.B(n_2929),
.Y(n_4617)
);

INVx4_ASAP7_75t_L g4618 ( 
.A(n_4019),
.Y(n_4618)
);

NAND2x1p5_ASAP7_75t_L g4619 ( 
.A(n_3994),
.B(n_2787),
.Y(n_4619)
);

BUFx4f_ASAP7_75t_L g4620 ( 
.A(n_4036),
.Y(n_4620)
);

BUFx6f_ASAP7_75t_L g4621 ( 
.A(n_4036),
.Y(n_4621)
);

INVx2_ASAP7_75t_SL g4622 ( 
.A(n_4101),
.Y(n_4622)
);

BUFx6f_ASAP7_75t_L g4623 ( 
.A(n_4101),
.Y(n_4623)
);

OR2x6_ASAP7_75t_L g4624 ( 
.A(n_3998),
.B(n_4277),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4263),
.B(n_2871),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4187),
.Y(n_4626)
);

INVx3_ASAP7_75t_L g4627 ( 
.A(n_4101),
.Y(n_4627)
);

OR2x2_ASAP7_75t_L g4628 ( 
.A(n_4303),
.B(n_3998),
.Y(n_4628)
);

AOI22xp33_ASAP7_75t_L g4629 ( 
.A1(n_4279),
.A2(n_4043),
.B1(n_4163),
.B2(n_4083),
.Y(n_4629)
);

O2A1O1Ixp33_ASAP7_75t_L g4630 ( 
.A1(n_4421),
.A2(n_4419),
.B(n_4598),
.C(n_4576),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_SL g4631 ( 
.A(n_4455),
.B(n_4136),
.Y(n_4631)
);

BUFx6f_ASAP7_75t_L g4632 ( 
.A(n_4291),
.Y(n_4632)
);

NOR2xp33_ASAP7_75t_L g4633 ( 
.A(n_4288),
.B(n_4160),
.Y(n_4633)
);

AOI21xp5_ASAP7_75t_L g4634 ( 
.A1(n_4293),
.A2(n_4094),
.B(n_4118),
.Y(n_4634)
);

INVx4_ASAP7_75t_L g4635 ( 
.A(n_4397),
.Y(n_4635)
);

AOI21xp5_ASAP7_75t_L g4636 ( 
.A1(n_4293),
.A2(n_4419),
.B(n_4319),
.Y(n_4636)
);

AOI221xp5_ASAP7_75t_L g4637 ( 
.A1(n_4421),
.A2(n_4576),
.B1(n_4562),
.B2(n_4424),
.C(n_4371),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4544),
.B(n_4224),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4278),
.Y(n_4639)
);

OAI22xp5_ASAP7_75t_L g4640 ( 
.A1(n_4593),
.A2(n_4408),
.B1(n_4434),
.B2(n_4449),
.Y(n_4640)
);

AOI21xp5_ASAP7_75t_L g4641 ( 
.A1(n_4319),
.A2(n_4094),
.B(n_4118),
.Y(n_4641)
);

OR2x2_ASAP7_75t_L g4642 ( 
.A(n_4303),
.B(n_4304),
.Y(n_4642)
);

OAI21x1_ASAP7_75t_L g4643 ( 
.A1(n_4554),
.A2(n_4277),
.B(n_4190),
.Y(n_4643)
);

BUFx6f_ASAP7_75t_L g4644 ( 
.A(n_4397),
.Y(n_4644)
);

AND2x2_ASAP7_75t_SL g4645 ( 
.A(n_4292),
.B(n_4013),
.Y(n_4645)
);

INVx2_ASAP7_75t_L g4646 ( 
.A(n_4321),
.Y(n_4646)
);

AOI21xp5_ASAP7_75t_L g4647 ( 
.A1(n_4572),
.A2(n_4091),
.B(n_4247),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4597),
.B(n_4141),
.Y(n_4648)
);

INVx2_ASAP7_75t_SL g4649 ( 
.A(n_4541),
.Y(n_4649)
);

BUFx2_ASAP7_75t_L g4650 ( 
.A(n_4394),
.Y(n_4650)
);

OAI21xp33_ASAP7_75t_L g4651 ( 
.A1(n_4493),
.A2(n_1084),
.B(n_4215),
.Y(n_4651)
);

AOI22xp5_ASAP7_75t_L g4652 ( 
.A1(n_4287),
.A2(n_3986),
.B1(n_4054),
.B2(n_4178),
.Y(n_4652)
);

AOI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4572),
.A2(n_4091),
.B(n_4140),
.Y(n_4653)
);

HB1xp67_ASAP7_75t_L g4654 ( 
.A(n_4446),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_4506),
.B(n_4245),
.Y(n_4655)
);

OR2x6_ASAP7_75t_L g4656 ( 
.A(n_4329),
.B(n_4190),
.Y(n_4656)
);

O2A1O1Ixp33_ASAP7_75t_L g4657 ( 
.A1(n_4562),
.A2(n_4381),
.B(n_4473),
.C(n_4298),
.Y(n_4657)
);

AOI21xp5_ASAP7_75t_L g4658 ( 
.A1(n_4572),
.A2(n_4140),
.B(n_3992),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_SL g4659 ( 
.A(n_4343),
.B(n_4263),
.Y(n_4659)
);

NOR2xp33_ASAP7_75t_L g4660 ( 
.A(n_4313),
.B(n_4053),
.Y(n_4660)
);

OAI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_4392),
.A2(n_4114),
.B1(n_4107),
.B2(n_4203),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_SL g4662 ( 
.A(n_4520),
.B(n_4252),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4516),
.B(n_4254),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4516),
.B(n_4256),
.Y(n_4664)
);

A2O1A1Ixp33_ASAP7_75t_L g4665 ( 
.A1(n_4519),
.A2(n_4270),
.B(n_4114),
.C(n_4107),
.Y(n_4665)
);

A2O1A1Ixp33_ASAP7_75t_SL g4666 ( 
.A1(n_4605),
.A2(n_4194),
.B(n_4206),
.C(n_4244),
.Y(n_4666)
);

AOI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_4287),
.A2(n_770),
.B1(n_775),
.B2(n_768),
.Y(n_4667)
);

NOR2xp33_ASAP7_75t_SL g4668 ( 
.A(n_4316),
.B(n_3994),
.Y(n_4668)
);

BUFx3_ASAP7_75t_L g4669 ( 
.A(n_4296),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4580),
.B(n_4257),
.Y(n_4670)
);

OAI21xp33_ASAP7_75t_L g4671 ( 
.A1(n_4355),
.A2(n_904),
.B(n_903),
.Y(n_4671)
);

NOR3xp33_ASAP7_75t_SL g4672 ( 
.A(n_4610),
.B(n_909),
.C(n_907),
.Y(n_4672)
);

O2A1O1Ixp33_ASAP7_75t_L g4673 ( 
.A1(n_4473),
.A2(n_775),
.B(n_778),
.C(n_770),
.Y(n_4673)
);

NOR2x1_ASAP7_75t_L g4674 ( 
.A(n_4351),
.B(n_4133),
.Y(n_4674)
);

AOI21xp5_ASAP7_75t_L g4675 ( 
.A1(n_4329),
.A2(n_4168),
.B(n_4167),
.Y(n_4675)
);

NAND3xp33_ASAP7_75t_L g4676 ( 
.A(n_4613),
.B(n_789),
.C(n_786),
.Y(n_4676)
);

NOR2xp33_ASAP7_75t_L g4677 ( 
.A(n_4309),
.B(n_912),
.Y(n_4677)
);

AND2x4_ASAP7_75t_L g4678 ( 
.A(n_4290),
.B(n_4019),
.Y(n_4678)
);

INVx4_ASAP7_75t_L g4679 ( 
.A(n_4397),
.Y(n_4679)
);

AOI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4329),
.A2(n_4168),
.B(n_4167),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4323),
.B(n_4105),
.Y(n_4681)
);

OAI22xp5_ASAP7_75t_L g4682 ( 
.A1(n_4526),
.A2(n_4201),
.B1(n_4202),
.B2(n_4253),
.Y(n_4682)
);

AND2x4_ASAP7_75t_L g4683 ( 
.A(n_4290),
.B(n_4048),
.Y(n_4683)
);

NOR2xp67_ASAP7_75t_L g4684 ( 
.A(n_4363),
.B(n_4205),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_SL g4685 ( 
.A(n_4363),
.B(n_4210),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4283),
.Y(n_4686)
);

AND2x4_ASAP7_75t_L g4687 ( 
.A(n_4612),
.B(n_4048),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4295),
.Y(n_4688)
);

INVx5_ASAP7_75t_L g4689 ( 
.A(n_4607),
.Y(n_4689)
);

CKINVDCx16_ASAP7_75t_R g4690 ( 
.A(n_4353),
.Y(n_4690)
);

OAI21x1_ASAP7_75t_L g4691 ( 
.A1(n_4554),
.A2(n_4373),
.B(n_3550),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_SL g4692 ( 
.A(n_4363),
.B(n_4210),
.Y(n_4692)
);

NAND3xp33_ASAP7_75t_L g4693 ( 
.A(n_4460),
.B(n_810),
.C(n_809),
.Y(n_4693)
);

AOI21xp5_ASAP7_75t_L g4694 ( 
.A1(n_4373),
.A2(n_4214),
.B(n_3597),
.Y(n_4694)
);

NAND3xp33_ASAP7_75t_SL g4695 ( 
.A(n_4521),
.B(n_4564),
.C(n_4508),
.Y(n_4695)
);

AOI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4415),
.A2(n_4214),
.B(n_4137),
.Y(n_4696)
);

NAND3xp33_ASAP7_75t_SL g4697 ( 
.A(n_4564),
.B(n_915),
.C(n_913),
.Y(n_4697)
);

OA22x2_ASAP7_75t_L g4698 ( 
.A1(n_4588),
.A2(n_863),
.B1(n_889),
.B2(n_828),
.Y(n_4698)
);

AND2x4_ASAP7_75t_L g4699 ( 
.A(n_4626),
.B(n_4048),
.Y(n_4699)
);

NAND2x1p5_ASAP7_75t_L g4700 ( 
.A(n_4363),
.B(n_4079),
.Y(n_4700)
);

OAI22xp5_ASAP7_75t_L g4701 ( 
.A1(n_4518),
.A2(n_4195),
.B1(n_4069),
.B2(n_4119),
.Y(n_4701)
);

OAI22xp5_ASAP7_75t_L g4702 ( 
.A1(n_4282),
.A2(n_4195),
.B1(n_4069),
.B2(n_4119),
.Y(n_4702)
);

BUFx6f_ASAP7_75t_L g4703 ( 
.A(n_4413),
.Y(n_4703)
);

BUFx6f_ASAP7_75t_L g4704 ( 
.A(n_4413),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_SL g4705 ( 
.A(n_4400),
.B(n_4039),
.Y(n_4705)
);

AOI21xp5_ASAP7_75t_L g4706 ( 
.A1(n_4347),
.A2(n_3525),
.B(n_3259),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4469),
.B(n_4105),
.Y(n_4707)
);

CKINVDCx5p33_ASAP7_75t_R g4708 ( 
.A(n_4280),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4512),
.B(n_4105),
.Y(n_4709)
);

HB1xp67_ASAP7_75t_L g4710 ( 
.A(n_4444),
.Y(n_4710)
);

A2O1A1Ixp33_ASAP7_75t_L g4711 ( 
.A1(n_4356),
.A2(n_820),
.B(n_827),
.C(n_819),
.Y(n_4711)
);

INVx2_ASAP7_75t_L g4712 ( 
.A(n_4348),
.Y(n_4712)
);

NOR2xp33_ASAP7_75t_L g4713 ( 
.A(n_4556),
.B(n_917),
.Y(n_4713)
);

AOI22xp33_ASAP7_75t_L g4714 ( 
.A1(n_4318),
.A2(n_916),
.B1(n_918),
.B2(n_908),
.Y(n_4714)
);

NAND3xp33_ASAP7_75t_SL g4715 ( 
.A(n_4365),
.B(n_922),
.C(n_920),
.Y(n_4715)
);

INVxp67_ASAP7_75t_SL g4716 ( 
.A(n_4305),
.Y(n_4716)
);

AND2x2_ASAP7_75t_L g4717 ( 
.A(n_4512),
.B(n_4111),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4380),
.B(n_4111),
.Y(n_4718)
);

OAI22xp5_ASAP7_75t_L g4719 ( 
.A1(n_4282),
.A2(n_4039),
.B1(n_4079),
.B2(n_835),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_L g4720 ( 
.A(n_4583),
.B(n_4111),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4399),
.B(n_4079),
.Y(n_4721)
);

O2A1O1Ixp33_ASAP7_75t_L g4722 ( 
.A1(n_4534),
.A2(n_835),
.B(n_846),
.C(n_833),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4349),
.Y(n_4723)
);

OR2x2_ASAP7_75t_L g4724 ( 
.A(n_4304),
.B(n_1521),
.Y(n_4724)
);

AOI21xp5_ASAP7_75t_L g4725 ( 
.A1(n_4347),
.A2(n_3525),
.B(n_3259),
.Y(n_4725)
);

AND2x4_ASAP7_75t_L g4726 ( 
.A(n_4359),
.B(n_4368),
.Y(n_4726)
);

A2O1A1Ixp33_ASAP7_75t_SL g4727 ( 
.A1(n_4503),
.A2(n_1523),
.B(n_1524),
.C(n_1522),
.Y(n_4727)
);

BUFx12f_ASAP7_75t_L g4728 ( 
.A(n_4312),
.Y(n_4728)
);

AND2x4_ASAP7_75t_L g4729 ( 
.A(n_4359),
.B(n_3395),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_SL g4730 ( 
.A(n_4400),
.B(n_2062),
.Y(n_4730)
);

INVx2_ASAP7_75t_L g4731 ( 
.A(n_4366),
.Y(n_4731)
);

AOI21xp5_ASAP7_75t_L g4732 ( 
.A1(n_4326),
.A2(n_2789),
.B(n_2787),
.Y(n_4732)
);

NOR4xp25_ASAP7_75t_SL g4733 ( 
.A(n_4437),
.B(n_930),
.C(n_938),
.D(n_926),
.Y(n_4733)
);

BUFx6f_ASAP7_75t_L g4734 ( 
.A(n_4413),
.Y(n_4734)
);

AOI21xp5_ASAP7_75t_L g4735 ( 
.A1(n_4326),
.A2(n_2798),
.B(n_2789),
.Y(n_4735)
);

AOI21xp5_ASAP7_75t_L g4736 ( 
.A1(n_4327),
.A2(n_2798),
.B(n_2789),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4324),
.B(n_848),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4350),
.B(n_1311),
.Y(n_4738)
);

NOR2xp33_ASAP7_75t_L g4739 ( 
.A(n_4328),
.B(n_928),
.Y(n_4739)
);

CKINVDCx5p33_ASAP7_75t_R g4740 ( 
.A(n_4311),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4611),
.B(n_1311),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4611),
.B(n_1311),
.Y(n_4742)
);

CKINVDCx5p33_ASAP7_75t_R g4743 ( 
.A(n_4337),
.Y(n_4743)
);

NAND2x1p5_ASAP7_75t_L g4744 ( 
.A(n_4400),
.B(n_2798),
.Y(n_4744)
);

OR2x6_ASAP7_75t_L g4745 ( 
.A(n_4606),
.B(n_2808),
.Y(n_4745)
);

CKINVDCx20_ASAP7_75t_R g4746 ( 
.A(n_4565),
.Y(n_4746)
);

INVxp67_ASAP7_75t_SL g4747 ( 
.A(n_4405),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_SL g4748 ( 
.A(n_4402),
.B(n_2070),
.Y(n_4748)
);

OAI22xp5_ASAP7_75t_L g4749 ( 
.A1(n_4504),
.A2(n_4362),
.B1(n_4361),
.B2(n_4563),
.Y(n_4749)
);

NOR2xp33_ASAP7_75t_L g4750 ( 
.A(n_4331),
.B(n_4422),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4332),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_SL g4752 ( 
.A(n_4402),
.B(n_2070),
.Y(n_4752)
);

INVx4_ASAP7_75t_L g4753 ( 
.A(n_4607),
.Y(n_4753)
);

NOR3xp33_ASAP7_75t_L g4754 ( 
.A(n_4435),
.B(n_863),
.C(n_862),
.Y(n_4754)
);

INVx3_ASAP7_75t_SL g4755 ( 
.A(n_4312),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4333),
.Y(n_4756)
);

O2A1O1Ixp5_ASAP7_75t_SL g4757 ( 
.A1(n_4586),
.A2(n_866),
.B(n_867),
.C(n_865),
.Y(n_4757)
);

BUFx6f_ASAP7_75t_L g4758 ( 
.A(n_4575),
.Y(n_4758)
);

AOI21xp5_ASAP7_75t_L g4759 ( 
.A1(n_4294),
.A2(n_4317),
.B(n_4308),
.Y(n_4759)
);

A2O1A1Ixp33_ASAP7_75t_L g4760 ( 
.A1(n_4502),
.A2(n_866),
.B(n_867),
.C(n_865),
.Y(n_4760)
);

NOR3xp33_ASAP7_75t_L g4761 ( 
.A(n_4585),
.B(n_4284),
.C(n_4601),
.Y(n_4761)
);

NOR2xp33_ASAP7_75t_L g4762 ( 
.A(n_4360),
.B(n_931),
.Y(n_4762)
);

BUFx6f_ASAP7_75t_L g4763 ( 
.A(n_4500),
.Y(n_4763)
);

BUFx12f_ASAP7_75t_L g4764 ( 
.A(n_4461),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4470),
.B(n_868),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4433),
.B(n_868),
.Y(n_4766)
);

AOI21xp5_ASAP7_75t_L g4767 ( 
.A1(n_4317),
.A2(n_4388),
.B(n_4345),
.Y(n_4767)
);

AOI22xp5_ASAP7_75t_L g4768 ( 
.A1(n_4395),
.A2(n_877),
.B1(n_888),
.B2(n_871),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4314),
.B(n_1326),
.Y(n_4769)
);

OAI21x1_ASAP7_75t_L g4770 ( 
.A1(n_4466),
.A2(n_2897),
.B(n_2972),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4314),
.B(n_1326),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_SL g4772 ( 
.A(n_4402),
.B(n_2071),
.Y(n_4772)
);

AOI22xp33_ASAP7_75t_L g4773 ( 
.A1(n_4310),
.A2(n_4403),
.B1(n_4603),
.B2(n_4368),
.Y(n_4773)
);

A2O1A1Ixp33_ASAP7_75t_L g4774 ( 
.A1(n_4411),
.A2(n_896),
.B(n_897),
.C(n_894),
.Y(n_4774)
);

OAI22x1_ASAP7_75t_L g4775 ( 
.A1(n_4361),
.A2(n_896),
.B1(n_897),
.B2(n_894),
.Y(n_4775)
);

OAI22xp5_ASAP7_75t_L g4776 ( 
.A1(n_4310),
.A2(n_4384),
.B1(n_4547),
.B2(n_4364),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_SL g4777 ( 
.A(n_4467),
.B(n_4481),
.Y(n_4777)
);

A2O1A1Ixp33_ASAP7_75t_SL g4778 ( 
.A1(n_4475),
.A2(n_1526),
.B(n_1528),
.C(n_1525),
.Y(n_4778)
);

AOI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4345),
.A2(n_2839),
.B(n_2808),
.Y(n_4779)
);

A2O1A1Ixp33_ASAP7_75t_L g4780 ( 
.A1(n_4401),
.A2(n_906),
.B(n_911),
.C(n_905),
.Y(n_4780)
);

BUFx6f_ASAP7_75t_L g4781 ( 
.A(n_4548),
.Y(n_4781)
);

INVxp67_ASAP7_75t_L g4782 ( 
.A(n_4352),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4307),
.B(n_4376),
.Y(n_4783)
);

O2A1O1Ixp33_ASAP7_75t_L g4784 ( 
.A1(n_4412),
.A2(n_906),
.B(n_911),
.C(n_905),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4370),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4307),
.B(n_1326),
.Y(n_4786)
);

INVxp67_ASAP7_75t_L g4787 ( 
.A(n_4551),
.Y(n_4787)
);

BUFx6f_ASAP7_75t_L g4788 ( 
.A(n_4548),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4377),
.Y(n_4789)
);

AOI21xp5_ASAP7_75t_L g4790 ( 
.A1(n_4388),
.A2(n_2839),
.B(n_2808),
.Y(n_4790)
);

OR2x6_ASAP7_75t_L g4791 ( 
.A(n_4374),
.B(n_2839),
.Y(n_4791)
);

BUFx6f_ASAP7_75t_L g4792 ( 
.A(n_4548),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4376),
.B(n_932),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4390),
.B(n_933),
.Y(n_4794)
);

NOR3xp33_ASAP7_75t_SL g4795 ( 
.A(n_4599),
.B(n_936),
.C(n_935),
.Y(n_4795)
);

OR2x6_ASAP7_75t_SL g4796 ( 
.A(n_4301),
.B(n_4579),
.Y(n_4796)
);

INVx3_ASAP7_75t_L g4797 ( 
.A(n_4325),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4340),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4410),
.A2(n_2879),
.B(n_2861),
.Y(n_4799)
);

HB1xp67_ASAP7_75t_L g4800 ( 
.A(n_4600),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4342),
.Y(n_4801)
);

OAI21x1_ASAP7_75t_L g4802 ( 
.A1(n_4466),
.A2(n_2879),
.B(n_2861),
.Y(n_4802)
);

INVxp67_ASAP7_75t_L g4803 ( 
.A(n_4407),
.Y(n_4803)
);

NAND2x1p5_ASAP7_75t_L g4804 ( 
.A(n_4481),
.B(n_2861),
.Y(n_4804)
);

AND2x4_ASAP7_75t_L g4805 ( 
.A(n_4403),
.B(n_3395),
.Y(n_4805)
);

AOI22xp33_ASAP7_75t_SL g4806 ( 
.A1(n_4302),
.A2(n_1060),
.B1(n_1072),
.B2(n_949),
.Y(n_4806)
);

INVx8_ASAP7_75t_L g4807 ( 
.A(n_4509),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4346),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4390),
.B(n_939),
.Y(n_4809)
);

OAI21x1_ASAP7_75t_L g4810 ( 
.A1(n_4386),
.A2(n_3229),
.B(n_3194),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4367),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4602),
.B(n_940),
.Y(n_4812)
);

AND2x4_ASAP7_75t_SL g4813 ( 
.A(n_4289),
.B(n_2898),
.Y(n_4813)
);

AND2x4_ASAP7_75t_L g4814 ( 
.A(n_4403),
.B(n_3611),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_4604),
.B(n_941),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4615),
.B(n_4479),
.Y(n_4816)
);

OR2x6_ASAP7_75t_L g4817 ( 
.A(n_4374),
.B(n_2876),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4489),
.B(n_4497),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4478),
.B(n_942),
.Y(n_4819)
);

AO21x1_ASAP7_75t_L g4820 ( 
.A1(n_4616),
.A2(n_945),
.B(n_944),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4369),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4379),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4382),
.Y(n_4823)
);

OR2x6_ASAP7_75t_L g4824 ( 
.A(n_4374),
.B(n_2876),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_4383),
.Y(n_4825)
);

BUFx3_ASAP7_75t_L g4826 ( 
.A(n_4430),
.Y(n_4826)
);

AOI22xp5_ASAP7_75t_L g4827 ( 
.A1(n_4301),
.A2(n_951),
.B1(n_952),
.B2(n_948),
.Y(n_4827)
);

O2A1O1Ixp33_ASAP7_75t_L g4828 ( 
.A1(n_4330),
.A2(n_4335),
.B(n_951),
.C(n_952),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4385),
.Y(n_4829)
);

BUFx6f_ASAP7_75t_L g4830 ( 
.A(n_4552),
.Y(n_4830)
);

BUFx12f_ASAP7_75t_L g4831 ( 
.A(n_4461),
.Y(n_4831)
);

BUFx12f_ASAP7_75t_L g4832 ( 
.A(n_4289),
.Y(n_4832)
);

BUFx6f_ASAP7_75t_SL g4833 ( 
.A(n_4445),
.Y(n_4833)
);

A2O1A1Ixp33_ASAP7_75t_L g4834 ( 
.A1(n_4496),
.A2(n_4501),
.B(n_4476),
.C(n_4471),
.Y(n_4834)
);

INVx5_ASAP7_75t_L g4835 ( 
.A(n_4618),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4404),
.Y(n_4836)
);

BUFx3_ASAP7_75t_L g4837 ( 
.A(n_4457),
.Y(n_4837)
);

AOI21xp5_ASAP7_75t_L g4838 ( 
.A1(n_4338),
.A2(n_3144),
.B(n_3138),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_SL g4839 ( 
.A(n_4496),
.B(n_2092),
.Y(n_4839)
);

OAI22xp5_ASAP7_75t_L g4840 ( 
.A1(n_4338),
.A2(n_966),
.B1(n_968),
.B2(n_964),
.Y(n_4840)
);

AOI21xp5_ASAP7_75t_L g4841 ( 
.A1(n_4487),
.A2(n_3144),
.B(n_3138),
.Y(n_4841)
);

AOI21xp5_ASAP7_75t_L g4842 ( 
.A1(n_4487),
.A2(n_4501),
.B(n_4496),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4418),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4420),
.Y(n_4844)
);

A2O1A1Ixp33_ASAP7_75t_SL g4845 ( 
.A1(n_4475),
.A2(n_1533),
.B(n_916),
.C(n_918),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_L g4846 ( 
.A(n_4568),
.B(n_943),
.Y(n_4846)
);

AOI21xp5_ASAP7_75t_L g4847 ( 
.A1(n_4487),
.A2(n_3144),
.B(n_3138),
.Y(n_4847)
);

OAI22xp5_ASAP7_75t_L g4848 ( 
.A1(n_4482),
.A2(n_4375),
.B1(n_4501),
.B2(n_4496),
.Y(n_4848)
);

A2O1A1Ixp33_ASAP7_75t_L g4849 ( 
.A1(n_4501),
.A2(n_973),
.B(n_974),
.C(n_971),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4423),
.Y(n_4850)
);

OAI22xp5_ASAP7_75t_L g4851 ( 
.A1(n_4375),
.A2(n_974),
.B1(n_976),
.B2(n_973),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4425),
.Y(n_4852)
);

INVx5_ASAP7_75t_L g4853 ( 
.A(n_4618),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4569),
.B(n_947),
.Y(n_4854)
);

BUFx2_ASAP7_75t_L g4855 ( 
.A(n_4442),
.Y(n_4855)
);

AND2x4_ASAP7_75t_L g4856 ( 
.A(n_4375),
.B(n_3611),
.Y(n_4856)
);

OAI21x1_ASAP7_75t_L g4857 ( 
.A1(n_4386),
.A2(n_3221),
.B(n_3214),
.Y(n_4857)
);

AOI21xp5_ASAP7_75t_L g4858 ( 
.A1(n_4417),
.A2(n_3144),
.B(n_3138),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4417),
.A2(n_2993),
.B(n_2961),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4596),
.B(n_4608),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4570),
.B(n_4573),
.Y(n_4861)
);

OAI22x1_ASAP7_75t_L g4862 ( 
.A1(n_4431),
.A2(n_982),
.B1(n_984),
.B2(n_978),
.Y(n_4862)
);

O2A1O1Ixp33_ASAP7_75t_L g4863 ( 
.A1(n_4452),
.A2(n_984),
.B(n_986),
.C(n_981),
.Y(n_4863)
);

INVx4_ASAP7_75t_L g4864 ( 
.A(n_4427),
.Y(n_4864)
);

BUFx2_ASAP7_75t_L g4865 ( 
.A(n_4529),
.Y(n_4865)
);

BUFx3_ASAP7_75t_L g4866 ( 
.A(n_4396),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4339),
.B(n_953),
.Y(n_4867)
);

BUFx6f_ASAP7_75t_L g4868 ( 
.A(n_4552),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4339),
.B(n_958),
.Y(n_4869)
);

NOR2xp33_ASAP7_75t_L g4870 ( 
.A(n_4582),
.B(n_959),
.Y(n_4870)
);

O2A1O1Ixp33_ASAP7_75t_L g4871 ( 
.A1(n_4477),
.A2(n_991),
.B(n_992),
.C(n_987),
.Y(n_4871)
);

OAI22xp5_ASAP7_75t_L g4872 ( 
.A1(n_4398),
.A2(n_4372),
.B1(n_4354),
.B2(n_4584),
.Y(n_4872)
);

HB1xp67_ASAP7_75t_L g4873 ( 
.A(n_4624),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4389),
.Y(n_4874)
);

NOR2xp67_ASAP7_75t_SL g4875 ( 
.A(n_4495),
.B(n_2793),
.Y(n_4875)
);

OAI22xp5_ASAP7_75t_SL g4876 ( 
.A1(n_4448),
.A2(n_993),
.B1(n_996),
.B2(n_990),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_4354),
.B(n_961),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4372),
.B(n_962),
.Y(n_4878)
);

AOI21xp5_ASAP7_75t_L g4879 ( 
.A1(n_4525),
.A2(n_4406),
.B(n_4617),
.Y(n_4879)
);

O2A1O1Ixp33_ASAP7_75t_L g4880 ( 
.A1(n_4477),
.A2(n_997),
.B(n_1004),
.C(n_993),
.Y(n_4880)
);

BUFx6f_ASAP7_75t_L g4881 ( 
.A(n_4552),
.Y(n_4881)
);

AND2x2_ASAP7_75t_SL g4882 ( 
.A(n_4322),
.B(n_908),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4409),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4451),
.Y(n_4884)
);

BUFx2_ASAP7_75t_L g4885 ( 
.A(n_4578),
.Y(n_4885)
);

INVx2_ASAP7_75t_L g4886 ( 
.A(n_4414),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4453),
.Y(n_4887)
);

NOR2xp67_ASAP7_75t_L g4888 ( 
.A(n_4559),
.B(n_4517),
.Y(n_4888)
);

BUFx6f_ASAP7_75t_L g4889 ( 
.A(n_4560),
.Y(n_4889)
);

INVx2_ASAP7_75t_L g4890 ( 
.A(n_4416),
.Y(n_4890)
);

NOR2xp33_ASAP7_75t_L g4891 ( 
.A(n_4589),
.B(n_970),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4465),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4522),
.Y(n_4893)
);

INVx3_ASAP7_75t_L g4894 ( 
.A(n_4325),
.Y(n_4894)
);

NOR2xp33_ASAP7_75t_L g4895 ( 
.A(n_4609),
.B(n_4281),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_SL g4896 ( 
.A(n_4358),
.B(n_2093),
.Y(n_4896)
);

INVx4_ASAP7_75t_L g4897 ( 
.A(n_4427),
.Y(n_4897)
);

A2O1A1Ixp33_ASAP7_75t_L g4898 ( 
.A1(n_4476),
.A2(n_1009),
.B(n_1011),
.C(n_1005),
.Y(n_4898)
);

NOR2xp33_ASAP7_75t_L g4899 ( 
.A(n_4299),
.B(n_977),
.Y(n_4899)
);

AND2x4_ASAP7_75t_L g4900 ( 
.A(n_4480),
.B(n_3611),
.Y(n_4900)
);

CKINVDCx6p67_ASAP7_75t_R g4901 ( 
.A(n_4325),
.Y(n_4901)
);

O2A1O1Ixp33_ASAP7_75t_L g4902 ( 
.A1(n_4458),
.A2(n_1009),
.B(n_1011),
.C(n_1005),
.Y(n_4902)
);

INVx1_ASAP7_75t_SL g4903 ( 
.A(n_4299),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4535),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4510),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4527),
.B(n_980),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_4530),
.Y(n_4907)
);

AOI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4591),
.A2(n_2958),
.B(n_2947),
.Y(n_4908)
);

BUFx6f_ASAP7_75t_L g4909 ( 
.A(n_4560),
.Y(n_4909)
);

INVx2_ASAP7_75t_SL g4910 ( 
.A(n_4560),
.Y(n_4910)
);

O2A1O1Ixp33_ASAP7_75t_L g4911 ( 
.A1(n_4458),
.A2(n_1019),
.B(n_1022),
.C(n_1016),
.Y(n_4911)
);

AOI21xp5_ASAP7_75t_L g4912 ( 
.A1(n_4591),
.A2(n_2979),
.B(n_2947),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4536),
.Y(n_4913)
);

INVx3_ASAP7_75t_L g4914 ( 
.A(n_4336),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_4532),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4546),
.Y(n_4916)
);

INVx2_ASAP7_75t_L g4917 ( 
.A(n_4533),
.Y(n_4917)
);

HB1xp67_ASAP7_75t_L g4918 ( 
.A(n_4553),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_SL g4919 ( 
.A(n_4491),
.B(n_3326),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_L g4920 ( 
.A1(n_4614),
.A2(n_2981),
.B(n_2979),
.Y(n_4920)
);

AOI21xp5_ASAP7_75t_L g4921 ( 
.A1(n_4614),
.A2(n_2981),
.B(n_2979),
.Y(n_4921)
);

A2O1A1Ixp33_ASAP7_75t_SL g4922 ( 
.A1(n_4488),
.A2(n_954),
.B(n_967),
.C(n_929),
.Y(n_4922)
);

HB1xp67_ASAP7_75t_L g4923 ( 
.A(n_4558),
.Y(n_4923)
);

AND2x2_ASAP7_75t_L g4924 ( 
.A(n_4538),
.B(n_1016),
.Y(n_4924)
);

BUFx6f_ASAP7_75t_L g4925 ( 
.A(n_4581),
.Y(n_4925)
);

BUFx6f_ASAP7_75t_L g4926 ( 
.A(n_4581),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4639),
.Y(n_4927)
);

BUFx3_ASAP7_75t_L g4928 ( 
.A(n_4746),
.Y(n_4928)
);

AOI211x1_ASAP7_75t_L g4929 ( 
.A1(n_4695),
.A2(n_1038),
.B(n_1043),
.C(n_1033),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4747),
.B(n_4566),
.Y(n_4930)
);

AOI21xp5_ASAP7_75t_L g4931 ( 
.A1(n_4636),
.A2(n_4511),
.B(n_4507),
.Y(n_4931)
);

OAI21xp5_ASAP7_75t_L g4932 ( 
.A1(n_4630),
.A2(n_4590),
.B(n_4387),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4654),
.B(n_4555),
.Y(n_4933)
);

OAI21xp5_ASAP7_75t_L g4934 ( 
.A1(n_4657),
.A2(n_4485),
.B(n_4472),
.Y(n_4934)
);

AOI21xp5_ASAP7_75t_L g4935 ( 
.A1(n_4658),
.A2(n_4511),
.B(n_4507),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4918),
.Y(n_4936)
);

O2A1O1Ixp33_ASAP7_75t_L g4937 ( 
.A1(n_4637),
.A2(n_1043),
.B(n_1046),
.C(n_1038),
.Y(n_4937)
);

HB1xp67_ASAP7_75t_L g4938 ( 
.A(n_4710),
.Y(n_4938)
);

INVx2_ASAP7_75t_SL g4939 ( 
.A(n_4632),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4783),
.B(n_4696),
.Y(n_4940)
);

AO31x2_ASAP7_75t_L g4941 ( 
.A1(n_4842),
.A2(n_4571),
.A3(n_4577),
.B(n_4528),
.Y(n_4941)
);

AOI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_4640),
.A2(n_4485),
.B1(n_4450),
.B2(n_4462),
.Y(n_4942)
);

NOR2xp33_ASAP7_75t_L g4943 ( 
.A(n_4633),
.B(n_4336),
.Y(n_4943)
);

AOI21x1_ASAP7_75t_L g4944 ( 
.A1(n_4631),
.A2(n_4472),
.B(n_4459),
.Y(n_4944)
);

AOI21x1_ASAP7_75t_SL g4945 ( 
.A1(n_4867),
.A2(n_4877),
.B(n_4869),
.Y(n_4945)
);

AOI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_4759),
.A2(n_4528),
.B(n_4515),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4923),
.Y(n_4947)
);

AOI21xp5_ASAP7_75t_L g4948 ( 
.A1(n_4767),
.A2(n_4653),
.B(n_4675),
.Y(n_4948)
);

AO31x2_ASAP7_75t_L g4949 ( 
.A1(n_4641),
.A2(n_4571),
.A3(n_4577),
.B(n_4539),
.Y(n_4949)
);

A2O1A1Ixp33_ASAP7_75t_L g4950 ( 
.A1(n_4651),
.A2(n_1048),
.B(n_1049),
.C(n_1046),
.Y(n_4950)
);

OAI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4667),
.A2(n_4459),
.B(n_4450),
.Y(n_4951)
);

OA21x2_ASAP7_75t_L g4952 ( 
.A1(n_4879),
.A2(n_4484),
.B(n_4483),
.Y(n_4952)
);

OAI21x1_ASAP7_75t_L g4953 ( 
.A1(n_4841),
.A2(n_4539),
.B(n_4515),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4716),
.B(n_4436),
.Y(n_4954)
);

AOI21xp5_ASAP7_75t_L g4955 ( 
.A1(n_4680),
.A2(n_4550),
.B(n_4545),
.Y(n_4955)
);

A2O1A1Ixp33_ASAP7_75t_L g4956 ( 
.A1(n_4828),
.A2(n_1049),
.B(n_1052),
.C(n_1048),
.Y(n_4956)
);

OAI21x1_ASAP7_75t_L g4957 ( 
.A1(n_4847),
.A2(n_4486),
.B(n_4484),
.Y(n_4957)
);

BUFx2_ASAP7_75t_L g4958 ( 
.A(n_4865),
.Y(n_4958)
);

INVx8_ASAP7_75t_L g4959 ( 
.A(n_4728),
.Y(n_4959)
);

AOI22xp5_ASAP7_75t_L g4960 ( 
.A1(n_4761),
.A2(n_4462),
.B1(n_4436),
.B2(n_4549),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4642),
.B(n_4285),
.Y(n_4961)
);

BUFx12f_ASAP7_75t_L g4962 ( 
.A(n_4743),
.Y(n_4962)
);

NOR2xp33_ASAP7_75t_SL g4963 ( 
.A(n_4708),
.B(n_4882),
.Y(n_4963)
);

AO31x2_ASAP7_75t_L g4964 ( 
.A1(n_4848),
.A2(n_4550),
.A3(n_4557),
.B(n_4545),
.Y(n_4964)
);

BUFx6f_ASAP7_75t_L g4965 ( 
.A(n_4632),
.Y(n_4965)
);

AOI21xp5_ASAP7_75t_L g4966 ( 
.A1(n_4694),
.A2(n_4561),
.B(n_4557),
.Y(n_4966)
);

OAI21x1_ASAP7_75t_L g4967 ( 
.A1(n_4691),
.A2(n_4838),
.B(n_4858),
.Y(n_4967)
);

AOI21x1_ASAP7_75t_L g4968 ( 
.A1(n_4888),
.A2(n_4297),
.B(n_4286),
.Y(n_4968)
);

OR2x6_ASAP7_75t_L g4969 ( 
.A(n_4745),
.B(n_4509),
.Y(n_4969)
);

AOI21x1_ASAP7_75t_L g4970 ( 
.A1(n_4888),
.A2(n_4315),
.B(n_4300),
.Y(n_4970)
);

AOI21xp5_ASAP7_75t_L g4971 ( 
.A1(n_4634),
.A2(n_4567),
.B(n_4561),
.Y(n_4971)
);

OAI22xp5_ASAP7_75t_L g4972 ( 
.A1(n_4629),
.A2(n_4652),
.B1(n_4806),
.B2(n_4645),
.Y(n_4972)
);

OAI21xp5_ASAP7_75t_L g4973 ( 
.A1(n_4676),
.A2(n_4474),
.B(n_1065),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4686),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_SL g4975 ( 
.A(n_4674),
.B(n_4341),
.Y(n_4975)
);

BUFx2_ASAP7_75t_L g4976 ( 
.A(n_4885),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_SL g4977 ( 
.A(n_4668),
.B(n_4341),
.Y(n_4977)
);

HB1xp67_ASAP7_75t_L g4978 ( 
.A(n_4800),
.Y(n_4978)
);

OAI21x1_ASAP7_75t_L g4979 ( 
.A1(n_4706),
.A2(n_4625),
.B(n_4499),
.Y(n_4979)
);

NOR2xp67_ASAP7_75t_L g4980 ( 
.A(n_4649),
.B(n_4559),
.Y(n_4980)
);

NOR2xp33_ASAP7_75t_SL g4981 ( 
.A(n_4690),
.B(n_4306),
.Y(n_4981)
);

AO31x2_ASAP7_75t_L g4982 ( 
.A1(n_4725),
.A2(n_4820),
.A3(n_4647),
.B(n_4776),
.Y(n_4982)
);

INVx2_ASAP7_75t_L g4983 ( 
.A(n_4688),
.Y(n_4983)
);

AOI21xp5_ASAP7_75t_L g4984 ( 
.A1(n_4777),
.A2(n_4543),
.B(n_4490),
.Y(n_4984)
);

AOI21xp5_ASAP7_75t_L g4985 ( 
.A1(n_4684),
.A2(n_4498),
.B(n_4559),
.Y(n_4985)
);

AOI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4684),
.A2(n_4559),
.B(n_4620),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4726),
.B(n_4357),
.Y(n_4987)
);

OAI21x1_ASAP7_75t_L g4988 ( 
.A1(n_4643),
.A2(n_4619),
.B(n_4574),
.Y(n_4988)
);

OAI21x1_ASAP7_75t_L g4989 ( 
.A1(n_4770),
.A2(n_4619),
.B(n_4574),
.Y(n_4989)
);

BUFx6f_ASAP7_75t_L g4990 ( 
.A(n_4632),
.Y(n_4990)
);

OAI21x1_ASAP7_75t_L g4991 ( 
.A1(n_4779),
.A2(n_4799),
.B(n_4790),
.Y(n_4991)
);

OAI21x1_ASAP7_75t_L g4992 ( 
.A1(n_4802),
.A2(n_4513),
.B(n_4488),
.Y(n_4992)
);

OAI21x1_ASAP7_75t_L g4993 ( 
.A1(n_4810),
.A2(n_4524),
.B(n_4513),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_4628),
.B(n_4655),
.Y(n_4994)
);

O2A1O1Ixp5_ASAP7_75t_SL g4995 ( 
.A1(n_4662),
.A2(n_1074),
.B(n_1077),
.C(n_1067),
.Y(n_4995)
);

BUFx2_ASAP7_75t_L g4996 ( 
.A(n_4855),
.Y(n_4996)
);

AO31x2_ASAP7_75t_L g4997 ( 
.A1(n_4702),
.A2(n_4428),
.A3(n_4456),
.B(n_4334),
.Y(n_4997)
);

OAI21x1_ASAP7_75t_L g4998 ( 
.A1(n_4857),
.A2(n_4524),
.B(n_4426),
.Y(n_4998)
);

AOI21x1_ASAP7_75t_SL g4999 ( 
.A1(n_4878),
.A2(n_4505),
.B(n_4549),
.Y(n_4999)
);

INVxp67_ASAP7_75t_L g5000 ( 
.A(n_4766),
.Y(n_5000)
);

OAI21x1_ASAP7_75t_L g5001 ( 
.A1(n_4732),
.A2(n_4432),
.B(n_4429),
.Y(n_5001)
);

OAI21x1_ASAP7_75t_L g5002 ( 
.A1(n_4735),
.A2(n_4440),
.B(n_4439),
.Y(n_5002)
);

OAI21x1_ASAP7_75t_L g5003 ( 
.A1(n_4736),
.A2(n_4443),
.B(n_4441),
.Y(n_5003)
);

BUFx6f_ASAP7_75t_L g5004 ( 
.A(n_4763),
.Y(n_5004)
);

AOI21xp5_ASAP7_75t_L g5005 ( 
.A1(n_4834),
.A2(n_4692),
.B(n_4685),
.Y(n_5005)
);

BUFx3_ASAP7_75t_L g5006 ( 
.A(n_4832),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4751),
.Y(n_5007)
);

CKINVDCx5p33_ASAP7_75t_R g5008 ( 
.A(n_4740),
.Y(n_5008)
);

BUFx2_ASAP7_75t_SL g5009 ( 
.A(n_4833),
.Y(n_5009)
);

INVx2_ASAP7_75t_SL g5010 ( 
.A(n_4763),
.Y(n_5010)
);

BUFx6f_ASAP7_75t_L g5011 ( 
.A(n_4763),
.Y(n_5011)
);

OAI21xp5_ASAP7_75t_SL g5012 ( 
.A1(n_4697),
.A2(n_1081),
.B(n_1079),
.Y(n_5012)
);

AO31x2_ASAP7_75t_L g5013 ( 
.A1(n_4872),
.A2(n_4514),
.A3(n_4523),
.B(n_4456),
.Y(n_5013)
);

OAI22xp5_ASAP7_75t_L g5014 ( 
.A1(n_4714),
.A2(n_4540),
.B1(n_4531),
.B2(n_4620),
.Y(n_5014)
);

OAI21xp5_ASAP7_75t_L g5015 ( 
.A1(n_4693),
.A2(n_1083),
.B(n_1081),
.Y(n_5015)
);

O2A1O1Ixp5_ASAP7_75t_SL g5016 ( 
.A1(n_4659),
.A2(n_1085),
.B(n_1083),
.C(n_4592),
.Y(n_5016)
);

AOI21xp5_ASAP7_75t_L g5017 ( 
.A1(n_4666),
.A2(n_4505),
.B(n_4514),
.Y(n_5017)
);

INVx3_ASAP7_75t_L g5018 ( 
.A(n_4753),
.Y(n_5018)
);

INVx2_ASAP7_75t_L g5019 ( 
.A(n_4756),
.Y(n_5019)
);

INVx3_ASAP7_75t_L g5020 ( 
.A(n_4753),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4816),
.B(n_4320),
.Y(n_5021)
);

OR2x2_ASAP7_75t_L g5022 ( 
.A(n_4873),
.B(n_4320),
.Y(n_5022)
);

AOI21xp5_ASAP7_75t_L g5023 ( 
.A1(n_4730),
.A2(n_4523),
.B(n_4540),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4798),
.Y(n_5024)
);

AO22x2_ASAP7_75t_L g5025 ( 
.A1(n_4801),
.A2(n_4622),
.B1(n_4595),
.B2(n_4378),
.Y(n_5025)
);

CKINVDCx9p33_ASAP7_75t_R g5026 ( 
.A(n_4650),
.Y(n_5026)
);

OAI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4863),
.A2(n_954),
.B(n_929),
.Y(n_5027)
);

AOI21xp5_ASAP7_75t_L g5028 ( 
.A1(n_4748),
.A2(n_2982),
.B(n_2981),
.Y(n_5028)
);

INVx2_ASAP7_75t_SL g5029 ( 
.A(n_4826),
.Y(n_5029)
);

A2O1A1Ixp33_ASAP7_75t_L g5030 ( 
.A1(n_4660),
.A2(n_4880),
.B(n_4871),
.C(n_4711),
.Y(n_5030)
);

OAI21x1_ASAP7_75t_L g5031 ( 
.A1(n_4908),
.A2(n_4627),
.B(n_4592),
.Y(n_5031)
);

OAI21x1_ASAP7_75t_L g5032 ( 
.A1(n_4912),
.A2(n_4627),
.B(n_4378),
.Y(n_5032)
);

AO31x2_ASAP7_75t_L g5033 ( 
.A1(n_4701),
.A2(n_1014),
.A3(n_1042),
.B(n_967),
.Y(n_5033)
);

OAI21xp5_ASAP7_75t_L g5034 ( 
.A1(n_4739),
.A2(n_1042),
.B(n_1014),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_L g5035 ( 
.A(n_4782),
.B(n_4344),
.Y(n_5035)
);

AOI21xp5_ASAP7_75t_L g5036 ( 
.A1(n_4752),
.A2(n_3003),
.B(n_2982),
.Y(n_5036)
);

INVx3_ASAP7_75t_L g5037 ( 
.A(n_4905),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_4663),
.B(n_4454),
.Y(n_5038)
);

NAND3x1_ASAP7_75t_L g5039 ( 
.A(n_4750),
.B(n_4454),
.C(n_4393),
.Y(n_5039)
);

OAI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4902),
.A2(n_1073),
.B(n_1042),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4664),
.B(n_4391),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4737),
.B(n_4391),
.Y(n_5042)
);

AOI21xp5_ASAP7_75t_L g5043 ( 
.A1(n_4772),
.A2(n_3003),
.B(n_2982),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4808),
.Y(n_5044)
);

NOR2xp67_ASAP7_75t_L g5045 ( 
.A(n_4787),
.B(n_4391),
.Y(n_5045)
);

AOI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4839),
.A2(n_3012),
.B(n_3003),
.Y(n_5046)
);

CKINVDCx20_ASAP7_75t_R g5047 ( 
.A(n_4669),
.Y(n_5047)
);

INVx5_ASAP7_75t_L g5048 ( 
.A(n_4745),
.Y(n_5048)
);

OAI21xp5_ASAP7_75t_L g5049 ( 
.A1(n_4911),
.A2(n_1073),
.B(n_1070),
.Y(n_5049)
);

AND2x6_ASAP7_75t_L g5050 ( 
.A(n_4856),
.B(n_4427),
.Y(n_5050)
);

AOI21xp33_ASAP7_75t_L g5051 ( 
.A1(n_4719),
.A2(n_4447),
.B(n_4438),
.Y(n_5051)
);

OA21x2_ASAP7_75t_L g5052 ( 
.A1(n_4773),
.A2(n_995),
.B(n_988),
.Y(n_5052)
);

OAI21x1_ASAP7_75t_L g5053 ( 
.A1(n_4920),
.A2(n_4921),
.B(n_4705),
.Y(n_5053)
);

OAI21xp5_ASAP7_75t_L g5054 ( 
.A1(n_4677),
.A2(n_999),
.B(n_998),
.Y(n_5054)
);

BUFx3_ASAP7_75t_L g5055 ( 
.A(n_4837),
.Y(n_5055)
);

INVx3_ASAP7_75t_L g5056 ( 
.A(n_4907),
.Y(n_5056)
);

AOI21xp5_ASAP7_75t_L g5057 ( 
.A1(n_4656),
.A2(n_3014),
.B(n_3012),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_L g5058 ( 
.A(n_4861),
.B(n_4594),
.Y(n_5058)
);

OAI21x1_ASAP7_75t_L g5059 ( 
.A1(n_4700),
.A2(n_3194),
.B(n_3184),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_4915),
.B(n_4594),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_4917),
.B(n_4621),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_4648),
.B(n_4621),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4764),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4811),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4821),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_4822),
.Y(n_5066)
);

BUFx2_ASAP7_75t_L g5067 ( 
.A(n_4717),
.Y(n_5067)
);

OAI21x1_ASAP7_75t_L g5068 ( 
.A1(n_4757),
.A2(n_4771),
.B(n_4769),
.Y(n_5068)
);

BUFx6f_ASAP7_75t_L g5069 ( 
.A(n_4755),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4818),
.B(n_4621),
.Y(n_5070)
);

INVxp67_ASAP7_75t_L g5071 ( 
.A(n_4765),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4638),
.B(n_4623),
.Y(n_5072)
);

OAI22xp5_ASAP7_75t_L g5073 ( 
.A1(n_4749),
.A2(n_4447),
.B1(n_4464),
.B2(n_4438),
.Y(n_5073)
);

INVx5_ASAP7_75t_L g5074 ( 
.A(n_4831),
.Y(n_5074)
);

BUFx6f_ASAP7_75t_L g5075 ( 
.A(n_4758),
.Y(n_5075)
);

AOI21x1_ASAP7_75t_L g5076 ( 
.A1(n_4793),
.A2(n_2928),
.B(n_2899),
.Y(n_5076)
);

AOI21xp5_ASAP7_75t_L g5077 ( 
.A1(n_4656),
.A2(n_3014),
.B(n_3012),
.Y(n_5077)
);

INVx8_ASAP7_75t_L g5078 ( 
.A(n_4833),
.Y(n_5078)
);

OAI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_4774),
.A2(n_4780),
.B(n_4760),
.Y(n_5079)
);

AO31x2_ASAP7_75t_L g5080 ( 
.A1(n_4665),
.A2(n_4661),
.A3(n_4682),
.B(n_4893),
.Y(n_5080)
);

AND2x2_ASAP7_75t_L g5081 ( 
.A(n_4681),
.B(n_4438),
.Y(n_5081)
);

AOI21xp5_ASAP7_75t_L g5082 ( 
.A1(n_4656),
.A2(n_3014),
.B(n_3029),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_4904),
.B(n_4623),
.Y(n_5083)
);

AO31x2_ASAP7_75t_L g5084 ( 
.A1(n_4913),
.A2(n_2928),
.A3(n_2899),
.B(n_3184),
.Y(n_5084)
);

OAI21xp5_ASAP7_75t_L g5085 ( 
.A1(n_4827),
.A2(n_1007),
.B(n_1006),
.Y(n_5085)
);

AND2x6_ASAP7_75t_L g5086 ( 
.A(n_4856),
.B(n_4447),
.Y(n_5086)
);

NAND3xp33_ASAP7_75t_SL g5087 ( 
.A(n_4713),
.B(n_4587),
.C(n_4542),
.Y(n_5087)
);

AOI21x1_ASAP7_75t_L g5088 ( 
.A1(n_4794),
.A2(n_3200),
.B(n_3197),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4916),
.B(n_4463),
.Y(n_5089)
);

A2O1A1Ixp33_ASAP7_75t_L g5090 ( 
.A1(n_4827),
.A2(n_1036),
.B(n_1055),
.C(n_1023),
.Y(n_5090)
);

AO31x2_ASAP7_75t_L g5091 ( 
.A1(n_4851),
.A2(n_3221),
.A3(n_3229),
.B(n_3214),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4829),
.B(n_4463),
.Y(n_5092)
);

NAND3xp33_ASAP7_75t_L g5093 ( 
.A(n_4754),
.B(n_4468),
.C(n_4464),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_4836),
.B(n_4464),
.Y(n_5094)
);

OAI21x1_ASAP7_75t_SL g5095 ( 
.A1(n_4670),
.A2(n_5),
.B(n_6),
.Y(n_5095)
);

INVx3_ASAP7_75t_L g5096 ( 
.A(n_4646),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4843),
.Y(n_5097)
);

AO21x1_ASAP7_75t_L g5098 ( 
.A1(n_4809),
.A2(n_6),
.B(n_7),
.Y(n_5098)
);

NAND2xp5_ASAP7_75t_L g5099 ( 
.A(n_4844),
.B(n_4850),
.Y(n_5099)
);

OAI21xp5_ASAP7_75t_L g5100 ( 
.A1(n_4840),
.A2(n_1018),
.B(n_1008),
.Y(n_5100)
);

BUFx2_ASAP7_75t_L g5101 ( 
.A(n_4796),
.Y(n_5101)
);

INVx4_ASAP7_75t_L g5102 ( 
.A(n_4781),
.Y(n_5102)
);

AO32x2_ASAP7_75t_L g5103 ( 
.A1(n_4876),
.A2(n_1072),
.A3(n_1060),
.B1(n_949),
.B2(n_2792),
.Y(n_5103)
);

AOI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4859),
.A2(n_4494),
.B(n_4468),
.Y(n_5104)
);

AND2x4_ASAP7_75t_L g5105 ( 
.A(n_4852),
.B(n_4468),
.Y(n_5105)
);

BUFx6f_ASAP7_75t_L g5106 ( 
.A(n_4758),
.Y(n_5106)
);

INVx5_ASAP7_75t_L g5107 ( 
.A(n_4689),
.Y(n_5107)
);

BUFx2_ASAP7_75t_L g5108 ( 
.A(n_4720),
.Y(n_5108)
);

AOI21x1_ASAP7_75t_L g5109 ( 
.A1(n_4786),
.A2(n_3211),
.B(n_3201),
.Y(n_5109)
);

INVxp67_ASAP7_75t_SL g5110 ( 
.A(n_4707),
.Y(n_5110)
);

BUFx6f_ASAP7_75t_L g5111 ( 
.A(n_4758),
.Y(n_5111)
);

AO21x2_ASAP7_75t_L g5112 ( 
.A1(n_4738),
.A2(n_4492),
.B(n_3109),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_SL g5113 ( 
.A(n_4724),
.B(n_4494),
.Y(n_5113)
);

NOR2xp67_ASAP7_75t_L g5114 ( 
.A(n_4803),
.B(n_4537),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4884),
.Y(n_5115)
);

NOR2xp33_ASAP7_75t_L g5116 ( 
.A(n_4866),
.B(n_4537),
.Y(n_5116)
);

AND2x2_ASAP7_75t_L g5117 ( 
.A(n_4721),
.B(n_4887),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4892),
.Y(n_5118)
);

OAI21x1_ASAP7_75t_L g5119 ( 
.A1(n_4744),
.A2(n_4804),
.B(n_4919),
.Y(n_5119)
);

AOI21x1_ASAP7_75t_L g5120 ( 
.A1(n_4741),
.A2(n_2129),
.B(n_2124),
.Y(n_5120)
);

OAI21x1_ASAP7_75t_L g5121 ( 
.A1(n_4896),
.A2(n_3123),
.B(n_3108),
.Y(n_5121)
);

AND2x4_ASAP7_75t_L g5122 ( 
.A(n_4817),
.B(n_4824),
.Y(n_5122)
);

AO21x2_ASAP7_75t_L g5123 ( 
.A1(n_4742),
.A2(n_3125),
.B(n_3123),
.Y(n_5123)
);

OAI21x1_ASAP7_75t_SL g5124 ( 
.A1(n_4860),
.A2(n_4709),
.B(n_4718),
.Y(n_5124)
);

INVx3_ASAP7_75t_L g5125 ( 
.A(n_4712),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4723),
.Y(n_5126)
);

OAI21x1_ASAP7_75t_L g5127 ( 
.A1(n_4731),
.A2(n_3129),
.B(n_3125),
.Y(n_5127)
);

HB1xp67_ASAP7_75t_L g5128 ( 
.A(n_4785),
.Y(n_5128)
);

AOI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_4778),
.A2(n_3023),
.B(n_3020),
.Y(n_5129)
);

OAI21x1_ASAP7_75t_L g5130 ( 
.A1(n_4789),
.A2(n_4825),
.B(n_4823),
.Y(n_5130)
);

BUFx10_ASAP7_75t_L g5131 ( 
.A(n_4762),
.Y(n_5131)
);

OA21x2_ASAP7_75t_L g5132 ( 
.A1(n_4874),
.A2(n_1035),
.B(n_1028),
.Y(n_5132)
);

BUFx4f_ASAP7_75t_L g5133 ( 
.A(n_4644),
.Y(n_5133)
);

AOI21xp5_ASAP7_75t_L g5134 ( 
.A1(n_4727),
.A2(n_4845),
.B(n_4824),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_4883),
.B(n_1039),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_L g5136 ( 
.A(n_4886),
.B(n_1044),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_L g5137 ( 
.A(n_4890),
.B(n_4924),
.Y(n_5137)
);

AOI21x1_ASAP7_75t_L g5138 ( 
.A1(n_4819),
.A2(n_2129),
.B(n_2124),
.Y(n_5138)
);

AO31x2_ASAP7_75t_L g5139 ( 
.A1(n_4849),
.A2(n_3136),
.A3(n_3137),
.B(n_3129),
.Y(n_5139)
);

OAI21x1_ASAP7_75t_L g5140 ( 
.A1(n_4797),
.A2(n_4914),
.B(n_4894),
.Y(n_5140)
);

NAND2xp5_ASAP7_75t_L g5141 ( 
.A(n_4895),
.B(n_1053),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4903),
.B(n_1057),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_SL g5143 ( 
.A(n_4689),
.B(n_1060),
.Y(n_5143)
);

AOI21xp5_ASAP7_75t_L g5144 ( 
.A1(n_4817),
.A2(n_3026),
.B(n_3023),
.Y(n_5144)
);

AOI21xp5_ASAP7_75t_L g5145 ( 
.A1(n_4817),
.A2(n_3027),
.B(n_3026),
.Y(n_5145)
);

AOI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4824),
.A2(n_3030),
.B(n_3027),
.Y(n_5146)
);

INVx3_ASAP7_75t_L g5147 ( 
.A(n_4864),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_4791),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_4791),
.Y(n_5149)
);

INVx2_ASAP7_75t_L g5150 ( 
.A(n_4791),
.Y(n_5150)
);

AO31x2_ASAP7_75t_L g5151 ( 
.A1(n_4862),
.A2(n_3137),
.A3(n_3139),
.B(n_3136),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4922),
.A2(n_4854),
.B(n_4846),
.Y(n_5152)
);

OAI21xp33_ASAP7_75t_L g5153 ( 
.A1(n_4671),
.A2(n_1062),
.B(n_1061),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_4812),
.B(n_1063),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_L g5155 ( 
.A(n_4815),
.B(n_1066),
.Y(n_5155)
);

AOI21xp5_ASAP7_75t_L g5156 ( 
.A1(n_4805),
.A2(n_4814),
.B(n_4715),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_4698),
.Y(n_5157)
);

INVx6_ASAP7_75t_SL g5158 ( 
.A(n_4678),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_4678),
.B(n_4683),
.Y(n_5159)
);

OAI22x1_ASAP7_75t_L g5160 ( 
.A1(n_4814),
.A2(n_1076),
.B1(n_1078),
.B2(n_1075),
.Y(n_5160)
);

AND2x2_ASAP7_75t_L g5161 ( 
.A(n_4683),
.B(n_1072),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4687),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4687),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4699),
.Y(n_5164)
);

NOR2xp67_ASAP7_75t_L g5165 ( 
.A(n_4689),
.B(n_7),
.Y(n_5165)
);

BUFx6f_ASAP7_75t_L g5166 ( 
.A(n_4644),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_4699),
.Y(n_5167)
);

AOI21x1_ASAP7_75t_SL g5168 ( 
.A1(n_4906),
.A2(n_10),
.B(n_9),
.Y(n_5168)
);

INVx1_ASAP7_75t_SL g5169 ( 
.A(n_4644),
.Y(n_5169)
);

INVx3_ASAP7_75t_L g5170 ( 
.A(n_4864),
.Y(n_5170)
);

AND2x2_ASAP7_75t_L g5171 ( 
.A(n_4729),
.B(n_34),
.Y(n_5171)
);

AOI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_4835),
.A2(n_3033),
.B(n_2901),
.Y(n_5172)
);

NAND2x1p5_ASAP7_75t_L g5173 ( 
.A(n_4835),
.B(n_3130),
.Y(n_5173)
);

INVx4_ASAP7_75t_L g5174 ( 
.A(n_4781),
.Y(n_5174)
);

NAND2x1_ASAP7_75t_L g5175 ( 
.A(n_4897),
.B(n_2841),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_4775),
.B(n_34),
.Y(n_5176)
);

AND2x4_ASAP7_75t_L g5177 ( 
.A(n_4897),
.B(n_3053),
.Y(n_5177)
);

AND2x4_ASAP7_75t_L g5178 ( 
.A(n_4900),
.B(n_3053),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_4722),
.Y(n_5179)
);

OA21x2_ASAP7_75t_L g5180 ( 
.A1(n_4898),
.A2(n_3143),
.B(n_3141),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_4784),
.Y(n_5181)
);

AOI21xp5_ASAP7_75t_L g5182 ( 
.A1(n_4853),
.A2(n_2901),
.B(n_2900),
.Y(n_5182)
);

OA21x2_ASAP7_75t_L g5183 ( 
.A1(n_4768),
.A2(n_3145),
.B(n_3143),
.Y(n_5183)
);

OAI22xp33_ASAP7_75t_L g5184 ( 
.A1(n_4972),
.A2(n_4853),
.B1(n_4807),
.B2(n_4679),
.Y(n_5184)
);

INVx4_ASAP7_75t_L g5185 ( 
.A(n_5078),
.Y(n_5185)
);

BUFx6f_ASAP7_75t_L g5186 ( 
.A(n_5069),
.Y(n_5186)
);

INVx5_ASAP7_75t_L g5187 ( 
.A(n_5078),
.Y(n_5187)
);

AOI21xp5_ASAP7_75t_L g5188 ( 
.A1(n_4948),
.A2(n_4807),
.B(n_4673),
.Y(n_5188)
);

AND2x4_ASAP7_75t_L g5189 ( 
.A(n_5159),
.B(n_4910),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_5067),
.B(n_4635),
.Y(n_5190)
);

AND2x2_ASAP7_75t_L g5191 ( 
.A(n_5108),
.B(n_4635),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4927),
.Y(n_5192)
);

OAI22xp5_ASAP7_75t_L g5193 ( 
.A1(n_5030),
.A2(n_4795),
.B1(n_4679),
.B2(n_4768),
.Y(n_5193)
);

AOI21xp33_ASAP7_75t_SL g5194 ( 
.A1(n_4959),
.A2(n_4899),
.B(n_4891),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_4927),
.Y(n_5195)
);

AND2x4_ASAP7_75t_L g5196 ( 
.A(n_5162),
.B(n_4894),
.Y(n_5196)
);

OR2x2_ASAP7_75t_L g5197 ( 
.A(n_4938),
.B(n_4914),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_4940),
.B(n_4870),
.Y(n_5198)
);

NOR2xp33_ASAP7_75t_L g5199 ( 
.A(n_5069),
.B(n_4703),
.Y(n_5199)
);

AND2x2_ASAP7_75t_L g5200 ( 
.A(n_4958),
.B(n_4901),
.Y(n_5200)
);

NAND2xp5_ASAP7_75t_L g5201 ( 
.A(n_5110),
.B(n_4788),
.Y(n_5201)
);

AOI21xp5_ASAP7_75t_L g5202 ( 
.A1(n_5034),
.A2(n_4733),
.B(n_4813),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_4994),
.B(n_4788),
.Y(n_5203)
);

AOI21xp5_ASAP7_75t_L g5204 ( 
.A1(n_4966),
.A2(n_4704),
.B(n_4703),
.Y(n_5204)
);

AOI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_5152),
.A2(n_4704),
.B(n_4703),
.Y(n_5205)
);

AND2x4_ASAP7_75t_L g5206 ( 
.A(n_5163),
.B(n_4788),
.Y(n_5206)
);

O2A1O1Ixp5_ASAP7_75t_SL g5207 ( 
.A1(n_4975),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_5207)
);

AOI21xp5_ASAP7_75t_L g5208 ( 
.A1(n_4955),
.A2(n_4931),
.B(n_4935),
.Y(n_5208)
);

INVx3_ASAP7_75t_L g5209 ( 
.A(n_5140),
.Y(n_5209)
);

OA21x2_ASAP7_75t_L g5210 ( 
.A1(n_5005),
.A2(n_4672),
.B(n_3146),
.Y(n_5210)
);

OA21x2_ASAP7_75t_L g5211 ( 
.A1(n_5053),
.A2(n_3146),
.B(n_3145),
.Y(n_5211)
);

AOI21xp5_ASAP7_75t_L g5212 ( 
.A1(n_4971),
.A2(n_4734),
.B(n_4792),
.Y(n_5212)
);

AOI21xp5_ASAP7_75t_L g5213 ( 
.A1(n_4946),
.A2(n_4830),
.B(n_4792),
.Y(n_5213)
);

AND2x4_ASAP7_75t_L g5214 ( 
.A(n_5164),
.B(n_4792),
.Y(n_5214)
);

INVxp67_ASAP7_75t_L g5215 ( 
.A(n_4978),
.Y(n_5215)
);

NAND2x1p5_ASAP7_75t_L g5216 ( 
.A(n_5048),
.B(n_4875),
.Y(n_5216)
);

CKINVDCx5p33_ASAP7_75t_R g5217 ( 
.A(n_5008),
.Y(n_5217)
);

AOI22xp33_ASAP7_75t_L g5218 ( 
.A1(n_5101),
.A2(n_4868),
.B1(n_4881),
.B2(n_4830),
.Y(n_5218)
);

A2O1A1Ixp33_ASAP7_75t_L g5219 ( 
.A1(n_5012),
.A2(n_4868),
.B(n_4881),
.C(n_4830),
.Y(n_5219)
);

NAND2xp5_ASAP7_75t_L g5220 ( 
.A(n_4961),
.B(n_4868),
.Y(n_5220)
);

BUFx4f_ASAP7_75t_L g5221 ( 
.A(n_4959),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_5124),
.Y(n_5222)
);

INVx2_ASAP7_75t_L g5223 ( 
.A(n_5025),
.Y(n_5223)
);

OAI22xp5_ASAP7_75t_L g5224 ( 
.A1(n_5093),
.A2(n_4889),
.B1(n_4909),
.B2(n_4881),
.Y(n_5224)
);

A2O1A1Ixp33_ASAP7_75t_SL g5225 ( 
.A1(n_4932),
.A2(n_2134),
.B(n_2133),
.C(n_2025),
.Y(n_5225)
);

OR2x2_ASAP7_75t_L g5226 ( 
.A(n_4936),
.B(n_4889),
.Y(n_5226)
);

AOI22xp33_ASAP7_75t_L g5227 ( 
.A1(n_5052),
.A2(n_4925),
.B1(n_4926),
.B2(n_4909),
.Y(n_5227)
);

AOI22xp33_ASAP7_75t_L g5228 ( 
.A1(n_5052),
.A2(n_4925),
.B1(n_4926),
.B2(n_4909),
.Y(n_5228)
);

OAI22xp5_ASAP7_75t_L g5229 ( 
.A1(n_4929),
.A2(n_4926),
.B1(n_4925),
.B2(n_3156),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_L g5230 ( 
.A(n_5038),
.B(n_35),
.Y(n_5230)
);

AOI21xp5_ASAP7_75t_L g5231 ( 
.A1(n_5079),
.A2(n_3156),
.B(n_3151),
.Y(n_5231)
);

BUFx2_ASAP7_75t_L g5232 ( 
.A(n_5158),
.Y(n_5232)
);

AND2x2_ASAP7_75t_L g5233 ( 
.A(n_4976),
.B(n_9),
.Y(n_5233)
);

BUFx4f_ASAP7_75t_SL g5234 ( 
.A(n_4962),
.Y(n_5234)
);

BUFx3_ASAP7_75t_L g5235 ( 
.A(n_5047),
.Y(n_5235)
);

AOI22xp33_ASAP7_75t_L g5236 ( 
.A1(n_5098),
.A2(n_2134),
.B1(n_2133),
.B2(n_3053),
.Y(n_5236)
);

AND2x2_ASAP7_75t_L g5237 ( 
.A(n_4996),
.B(n_11),
.Y(n_5237)
);

OR2x2_ASAP7_75t_L g5238 ( 
.A(n_4947),
.B(n_11),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_5025),
.Y(n_5239)
);

AOI21xp5_ASAP7_75t_L g5240 ( 
.A1(n_5134),
.A2(n_3161),
.B(n_3151),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_L g5241 ( 
.A(n_5021),
.B(n_36),
.Y(n_5241)
);

INVx4_ASAP7_75t_L g5242 ( 
.A(n_5074),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_4930),
.B(n_36),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_5037),
.Y(n_5244)
);

BUFx2_ASAP7_75t_L g5245 ( 
.A(n_5158),
.Y(n_5245)
);

BUFx3_ASAP7_75t_L g5246 ( 
.A(n_4928),
.Y(n_5246)
);

AOI22xp5_ASAP7_75t_L g5247 ( 
.A1(n_4963),
.A2(n_4942),
.B1(n_5179),
.B2(n_4960),
.Y(n_5247)
);

BUFx2_ASAP7_75t_L g5248 ( 
.A(n_5026),
.Y(n_5248)
);

AO32x2_ASAP7_75t_L g5249 ( 
.A1(n_5073),
.A2(n_2966),
.A3(n_2984),
.B1(n_2891),
.B2(n_2862),
.Y(n_5249)
);

NAND2xp33_ASAP7_75t_L g5250 ( 
.A(n_5074),
.B(n_5063),
.Y(n_5250)
);

NOR2x1_ASAP7_75t_L g5251 ( 
.A(n_5009),
.B(n_2862),
.Y(n_5251)
);

OR2x2_ASAP7_75t_L g5252 ( 
.A(n_4933),
.B(n_11),
.Y(n_5252)
);

INVx5_ASAP7_75t_L g5253 ( 
.A(n_5107),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5007),
.Y(n_5254)
);

BUFx2_ASAP7_75t_L g5255 ( 
.A(n_5147),
.Y(n_5255)
);

OAI22xp5_ASAP7_75t_L g5256 ( 
.A1(n_5179),
.A2(n_3165),
.B1(n_2966),
.B2(n_2984),
.Y(n_5256)
);

AND2x2_ASAP7_75t_SL g5257 ( 
.A(n_4981),
.B(n_4952),
.Y(n_5257)
);

CKINVDCx16_ASAP7_75t_R g5258 ( 
.A(n_5006),
.Y(n_5258)
);

BUFx6f_ASAP7_75t_L g5259 ( 
.A(n_5075),
.Y(n_5259)
);

NOR2xp33_ASAP7_75t_L g5260 ( 
.A(n_5131),
.B(n_38),
.Y(n_5260)
);

AOI22xp5_ASAP7_75t_L g5261 ( 
.A1(n_5087),
.A2(n_3343),
.B1(n_3326),
.B2(n_2020),
.Y(n_5261)
);

BUFx4f_ASAP7_75t_L g5262 ( 
.A(n_5075),
.Y(n_5262)
);

AND2x2_ASAP7_75t_L g5263 ( 
.A(n_5117),
.B(n_12),
.Y(n_5263)
);

NAND2x1p5_ASAP7_75t_L g5264 ( 
.A(n_5048),
.B(n_2841),
.Y(n_5264)
);

AND2x4_ASAP7_75t_L g5265 ( 
.A(n_5167),
.B(n_12),
.Y(n_5265)
);

OR2x2_ASAP7_75t_L g5266 ( 
.A(n_5128),
.B(n_13),
.Y(n_5266)
);

INVx3_ASAP7_75t_SL g5267 ( 
.A(n_5074),
.Y(n_5267)
);

AND2x4_ASAP7_75t_L g5268 ( 
.A(n_5148),
.B(n_13),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_5024),
.Y(n_5269)
);

OAI22xp5_ASAP7_75t_L g5270 ( 
.A1(n_5157),
.A2(n_2966),
.B1(n_2984),
.B2(n_2891),
.Y(n_5270)
);

BUFx6f_ASAP7_75t_L g5271 ( 
.A(n_5075),
.Y(n_5271)
);

OAI22xp5_ASAP7_75t_L g5272 ( 
.A1(n_5181),
.A2(n_3092),
.B1(n_3117),
.B2(n_2891),
.Y(n_5272)
);

NOR2xp33_ASAP7_75t_L g5273 ( 
.A(n_5131),
.B(n_38),
.Y(n_5273)
);

AOI21xp5_ASAP7_75t_L g5274 ( 
.A1(n_4984),
.A2(n_3117),
.B(n_3092),
.Y(n_5274)
);

CKINVDCx5p33_ASAP7_75t_R g5275 ( 
.A(n_5055),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5044),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_5064),
.Y(n_5277)
);

BUFx6f_ASAP7_75t_L g5278 ( 
.A(n_5106),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5065),
.Y(n_5279)
);

AND2x4_ASAP7_75t_L g5280 ( 
.A(n_5149),
.B(n_13),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_5097),
.Y(n_5281)
);

BUFx6f_ASAP7_75t_L g5282 ( 
.A(n_5106),
.Y(n_5282)
);

NAND2x1p5_ASAP7_75t_L g5283 ( 
.A(n_5048),
.B(n_2841),
.Y(n_5283)
);

O2A1O1Ixp5_ASAP7_75t_SL g5284 ( 
.A1(n_5143),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_5284)
);

INVx3_ASAP7_75t_L g5285 ( 
.A(n_5018),
.Y(n_5285)
);

INVx3_ASAP7_75t_L g5286 ( 
.A(n_5018),
.Y(n_5286)
);

AND2x2_ASAP7_75t_L g5287 ( 
.A(n_4954),
.B(n_4987),
.Y(n_5287)
);

INVxp67_ASAP7_75t_SL g5288 ( 
.A(n_5130),
.Y(n_5288)
);

A2O1A1Ixp33_ASAP7_75t_L g5289 ( 
.A1(n_4937),
.A2(n_41),
.B(n_42),
.C(n_40),
.Y(n_5289)
);

AND2x4_ASAP7_75t_L g5290 ( 
.A(n_5150),
.B(n_14),
.Y(n_5290)
);

BUFx12f_ASAP7_75t_L g5291 ( 
.A(n_5161),
.Y(n_5291)
);

AND2x2_ASAP7_75t_L g5292 ( 
.A(n_5081),
.B(n_15),
.Y(n_5292)
);

NAND2xp5_ASAP7_75t_L g5293 ( 
.A(n_5096),
.B(n_41),
.Y(n_5293)
);

BUFx3_ASAP7_75t_L g5294 ( 
.A(n_4965),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5115),
.Y(n_5295)
);

BUFx6f_ASAP7_75t_L g5296 ( 
.A(n_5106),
.Y(n_5296)
);

AOI21xp5_ASAP7_75t_L g5297 ( 
.A1(n_5017),
.A2(n_3117),
.B(n_3092),
.Y(n_5297)
);

HB1xp67_ASAP7_75t_L g5298 ( 
.A(n_5096),
.Y(n_5298)
);

INVx2_ASAP7_75t_SL g5299 ( 
.A(n_4965),
.Y(n_5299)
);

AND2x4_ASAP7_75t_L g5300 ( 
.A(n_5122),
.B(n_17),
.Y(n_5300)
);

AOI21xp5_ASAP7_75t_L g5301 ( 
.A1(n_4985),
.A2(n_3128),
.B(n_2874),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_5056),
.Y(n_5302)
);

BUFx6f_ASAP7_75t_L g5303 ( 
.A(n_5111),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_5118),
.Y(n_5304)
);

INVx3_ASAP7_75t_L g5305 ( 
.A(n_5020),
.Y(n_5305)
);

BUFx2_ASAP7_75t_L g5306 ( 
.A(n_5170),
.Y(n_5306)
);

NAND2x1p5_ASAP7_75t_L g5307 ( 
.A(n_5107),
.B(n_2841),
.Y(n_5307)
);

INVx1_ASAP7_75t_SL g5308 ( 
.A(n_4990),
.Y(n_5308)
);

BUFx12f_ASAP7_75t_SL g5309 ( 
.A(n_5111),
.Y(n_5309)
);

INVx2_ASAP7_75t_L g5310 ( 
.A(n_5125),
.Y(n_5310)
);

AND2x2_ASAP7_75t_L g5311 ( 
.A(n_4939),
.B(n_19),
.Y(n_5311)
);

CKINVDCx11_ASAP7_75t_R g5312 ( 
.A(n_5111),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_4974),
.Y(n_5313)
);

NAND2xp5_ASAP7_75t_L g5314 ( 
.A(n_5126),
.B(n_42),
.Y(n_5314)
);

OAI22xp5_ASAP7_75t_L g5315 ( 
.A1(n_5156),
.A2(n_3128),
.B1(n_2874),
.B2(n_3000),
.Y(n_5315)
);

BUFx12f_ASAP7_75t_L g5316 ( 
.A(n_5029),
.Y(n_5316)
);

OAI21xp33_ASAP7_75t_L g5317 ( 
.A1(n_4934),
.A2(n_2083),
.B(n_19),
.Y(n_5317)
);

BUFx2_ASAP7_75t_L g5318 ( 
.A(n_5039),
.Y(n_5318)
);

AND2x4_ASAP7_75t_L g5319 ( 
.A(n_5122),
.B(n_5105),
.Y(n_5319)
);

AOI21xp5_ASAP7_75t_L g5320 ( 
.A1(n_4956),
.A2(n_3128),
.B(n_2874),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_4983),
.Y(n_5321)
);

AND2x2_ASAP7_75t_L g5322 ( 
.A(n_5022),
.B(n_20),
.Y(n_5322)
);

BUFx6f_ASAP7_75t_L g5323 ( 
.A(n_4990),
.Y(n_5323)
);

INVx5_ASAP7_75t_L g5324 ( 
.A(n_5107),
.Y(n_5324)
);

INVx1_ASAP7_75t_SL g5325 ( 
.A(n_5004),
.Y(n_5325)
);

INVx3_ASAP7_75t_L g5326 ( 
.A(n_5020),
.Y(n_5326)
);

AND2x4_ASAP7_75t_L g5327 ( 
.A(n_5105),
.B(n_20),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5019),
.Y(n_5328)
);

OR2x6_ASAP7_75t_L g5329 ( 
.A(n_4977),
.B(n_2841),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5066),
.Y(n_5330)
);

AOI21xp5_ASAP7_75t_L g5331 ( 
.A1(n_5104),
.A2(n_3000),
.B(n_2874),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_5058),
.B(n_43),
.Y(n_5332)
);

CKINVDCx20_ASAP7_75t_R g5333 ( 
.A(n_5042),
.Y(n_5333)
);

INVx1_ASAP7_75t_SL g5334 ( 
.A(n_5004),
.Y(n_5334)
);

INVx3_ASAP7_75t_L g5335 ( 
.A(n_5004),
.Y(n_5335)
);

AOI21xp5_ASAP7_75t_L g5336 ( 
.A1(n_4986),
.A2(n_3000),
.B(n_2874),
.Y(n_5336)
);

NOR2x1_ASAP7_75t_L g5337 ( 
.A(n_4980),
.B(n_3000),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_L g5338 ( 
.A(n_5070),
.B(n_45),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_5099),
.Y(n_5339)
);

AOI22xp33_ASAP7_75t_L g5340 ( 
.A1(n_5132),
.A2(n_2065),
.B1(n_2676),
.B2(n_2665),
.Y(n_5340)
);

INVx2_ASAP7_75t_SL g5341 ( 
.A(n_5011),
.Y(n_5341)
);

AND2x2_ASAP7_75t_L g5342 ( 
.A(n_5000),
.B(n_21),
.Y(n_5342)
);

BUFx3_ASAP7_75t_L g5343 ( 
.A(n_5011),
.Y(n_5343)
);

AOI21xp5_ASAP7_75t_L g5344 ( 
.A1(n_5090),
.A2(n_3130),
.B(n_3070),
.Y(n_5344)
);

AOI22xp33_ASAP7_75t_L g5345 ( 
.A1(n_5132),
.A2(n_2678),
.B1(n_2686),
.B2(n_2676),
.Y(n_5345)
);

BUFx6f_ASAP7_75t_L g5346 ( 
.A(n_5166),
.Y(n_5346)
);

OAI22xp5_ASAP7_75t_L g5347 ( 
.A1(n_4969),
.A2(n_3130),
.B1(n_3171),
.B2(n_3070),
.Y(n_5347)
);

AND2x4_ASAP7_75t_L g5348 ( 
.A(n_4997),
.B(n_21),
.Y(n_5348)
);

AOI222xp33_ASAP7_75t_L g5349 ( 
.A1(n_5085),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.C1(n_24),
.C2(n_26),
.Y(n_5349)
);

OAI22xp5_ASAP7_75t_L g5350 ( 
.A1(n_4969),
.A2(n_3130),
.B1(n_3171),
.B2(n_3070),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_5041),
.B(n_46),
.Y(n_5351)
);

AND2x2_ASAP7_75t_L g5352 ( 
.A(n_5010),
.B(n_5071),
.Y(n_5352)
);

AND2x4_ASAP7_75t_L g5353 ( 
.A(n_4997),
.B(n_23),
.Y(n_5353)
);

AND2x4_ASAP7_75t_L g5354 ( 
.A(n_4997),
.B(n_24),
.Y(n_5354)
);

AND2x2_ASAP7_75t_L g5355 ( 
.A(n_5035),
.B(n_27),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_5083),
.Y(n_5356)
);

AOI21xp5_ASAP7_75t_L g5357 ( 
.A1(n_5054),
.A2(n_3171),
.B(n_2906),
.Y(n_5357)
);

BUFx6f_ASAP7_75t_L g5358 ( 
.A(n_5166),
.Y(n_5358)
);

INVx3_ASAP7_75t_L g5359 ( 
.A(n_5102),
.Y(n_5359)
);

OR2x6_ASAP7_75t_L g5360 ( 
.A(n_5045),
.B(n_3171),
.Y(n_5360)
);

OR2x6_ASAP7_75t_L g5361 ( 
.A(n_5114),
.B(n_1140),
.Y(n_5361)
);

BUFx12f_ASAP7_75t_L g5362 ( 
.A(n_5171),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5089),
.Y(n_5363)
);

OAI21xp33_ASAP7_75t_L g5364 ( 
.A1(n_5176),
.A2(n_27),
.B(n_28),
.Y(n_5364)
);

INVx5_ASAP7_75t_SL g5365 ( 
.A(n_5177),
.Y(n_5365)
);

BUFx6f_ASAP7_75t_L g5366 ( 
.A(n_5133),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_5092),
.Y(n_5367)
);

INVx1_ASAP7_75t_SL g5368 ( 
.A(n_5169),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_5062),
.B(n_48),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_4968),
.Y(n_5370)
);

INVx3_ASAP7_75t_L g5371 ( 
.A(n_5102),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5072),
.B(n_49),
.Y(n_5372)
);

INVxp67_ASAP7_75t_SL g5373 ( 
.A(n_5137),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_L g5374 ( 
.A(n_4949),
.B(n_50),
.Y(n_5374)
);

OAI22xp5_ASAP7_75t_L g5375 ( 
.A1(n_4943),
.A2(n_2907),
.B1(n_2908),
.B2(n_2900),
.Y(n_5375)
);

INVx1_ASAP7_75t_L g5376 ( 
.A(n_5094),
.Y(n_5376)
);

BUFx3_ASAP7_75t_L g5377 ( 
.A(n_5116),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_4941),
.Y(n_5378)
);

AOI21xp5_ASAP7_75t_L g5379 ( 
.A1(n_5057),
.A2(n_2908),
.B(n_2907),
.Y(n_5379)
);

AND2x4_ASAP7_75t_L g5380 ( 
.A(n_5013),
.B(n_28),
.Y(n_5380)
);

AO21x2_ASAP7_75t_L g5381 ( 
.A1(n_4944),
.A2(n_29),
.B(n_30),
.Y(n_5381)
);

NAND2x1p5_ASAP7_75t_L g5382 ( 
.A(n_5119),
.B(n_2676),
.Y(n_5382)
);

AOI22xp33_ASAP7_75t_L g5383 ( 
.A1(n_5153),
.A2(n_2686),
.B1(n_2694),
.B2(n_2678),
.Y(n_5383)
);

INVx2_ASAP7_75t_L g5384 ( 
.A(n_4970),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5013),
.Y(n_5385)
);

CKINVDCx5p33_ASAP7_75t_R g5386 ( 
.A(n_5133),
.Y(n_5386)
);

BUFx3_ASAP7_75t_L g5387 ( 
.A(n_5050),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_4941),
.Y(n_5388)
);

OAI22xp5_ASAP7_75t_L g5389 ( 
.A1(n_4951),
.A2(n_5165),
.B1(n_5113),
.B2(n_5014),
.Y(n_5389)
);

AND2x2_ASAP7_75t_SL g5390 ( 
.A(n_5174),
.B(n_51),
.Y(n_5390)
);

BUFx6f_ASAP7_75t_L g5391 ( 
.A(n_5175),
.Y(n_5391)
);

HB1xp67_ASAP7_75t_L g5392 ( 
.A(n_5013),
.Y(n_5392)
);

OR2x2_ASAP7_75t_SL g5393 ( 
.A(n_5141),
.B(n_30),
.Y(n_5393)
);

AOI22xp33_ASAP7_75t_L g5394 ( 
.A1(n_5160),
.A2(n_2686),
.B1(n_2694),
.B2(n_2678),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_4941),
.Y(n_5395)
);

CKINVDCx5p33_ASAP7_75t_R g5396 ( 
.A(n_5060),
.Y(n_5396)
);

A2O1A1Ixp33_ASAP7_75t_L g5397 ( 
.A1(n_5027),
.A2(n_53),
.B(n_54),
.C(n_52),
.Y(n_5397)
);

NAND2xp5_ASAP7_75t_L g5398 ( 
.A(n_4949),
.B(n_53),
.Y(n_5398)
);

HB1xp67_ASAP7_75t_L g5399 ( 
.A(n_4964),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_5192),
.Y(n_5400)
);

AOI22xp33_ASAP7_75t_L g5401 ( 
.A1(n_5208),
.A2(n_5040),
.B1(n_5049),
.B2(n_5095),
.Y(n_5401)
);

BUFx10_ASAP7_75t_L g5402 ( 
.A(n_5260),
.Y(n_5402)
);

INVx6_ASAP7_75t_L g5403 ( 
.A(n_5187),
.Y(n_5403)
);

AOI22xp33_ASAP7_75t_L g5404 ( 
.A1(n_5349),
.A2(n_5068),
.B1(n_5100),
.B2(n_5178),
.Y(n_5404)
);

AOI22xp33_ASAP7_75t_SL g5405 ( 
.A1(n_5257),
.A2(n_5080),
.B1(n_4973),
.B2(n_5086),
.Y(n_5405)
);

OAI22xp33_ASAP7_75t_L g5406 ( 
.A1(n_5248),
.A2(n_5077),
.B1(n_5080),
.B2(n_5051),
.Y(n_5406)
);

CKINVDCx20_ASAP7_75t_R g5407 ( 
.A(n_5234),
.Y(n_5407)
);

INVx1_ASAP7_75t_SL g5408 ( 
.A(n_5312),
.Y(n_5408)
);

AOI22xp33_ASAP7_75t_L g5409 ( 
.A1(n_5317),
.A2(n_5112),
.B1(n_5155),
.B2(n_5154),
.Y(n_5409)
);

INVx6_ASAP7_75t_L g5410 ( 
.A(n_5187),
.Y(n_5410)
);

BUFx2_ASAP7_75t_L g5411 ( 
.A(n_5267),
.Y(n_5411)
);

CKINVDCx11_ASAP7_75t_R g5412 ( 
.A(n_5258),
.Y(n_5412)
);

AOI22xp33_ASAP7_75t_SL g5413 ( 
.A1(n_5390),
.A2(n_5086),
.B1(n_5015),
.B2(n_5103),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_5195),
.Y(n_5414)
);

NAND2xp5_ASAP7_75t_L g5415 ( 
.A(n_5373),
.B(n_4964),
.Y(n_5415)
);

INVx2_ASAP7_75t_L g5416 ( 
.A(n_5222),
.Y(n_5416)
);

AOI21xp5_ASAP7_75t_SL g5417 ( 
.A1(n_5210),
.A2(n_5183),
.B(n_5173),
.Y(n_5417)
);

OAI22xp33_ASAP7_75t_R g5418 ( 
.A1(n_5273),
.A2(n_4945),
.B1(n_5103),
.B2(n_5168),
.Y(n_5418)
);

BUFx3_ASAP7_75t_L g5419 ( 
.A(n_5316),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_5209),
.Y(n_5420)
);

INVxp67_ASAP7_75t_L g5421 ( 
.A(n_5198),
.Y(n_5421)
);

AOI22xp33_ASAP7_75t_L g5422 ( 
.A1(n_5364),
.A2(n_5184),
.B1(n_5210),
.B2(n_5193),
.Y(n_5422)
);

AOI22xp33_ASAP7_75t_L g5423 ( 
.A1(n_5188),
.A2(n_4979),
.B1(n_4957),
.B2(n_4967),
.Y(n_5423)
);

INVx6_ASAP7_75t_L g5424 ( 
.A(n_5187),
.Y(n_5424)
);

INVx5_ASAP7_75t_L g5425 ( 
.A(n_5242),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_5209),
.Y(n_5426)
);

AOI22xp33_ASAP7_75t_SL g5427 ( 
.A1(n_5389),
.A2(n_5103),
.B1(n_4999),
.B2(n_5135),
.Y(n_5427)
);

INVx8_ASAP7_75t_L g5428 ( 
.A(n_5186),
.Y(n_5428)
);

BUFx3_ASAP7_75t_L g5429 ( 
.A(n_5235),
.Y(n_5429)
);

INVx1_ASAP7_75t_SL g5430 ( 
.A(n_5191),
.Y(n_5430)
);

AOI22xp33_ASAP7_75t_L g5431 ( 
.A1(n_5380),
.A2(n_5353),
.B1(n_5354),
.B2(n_5348),
.Y(n_5431)
);

INVx2_ASAP7_75t_SL g5432 ( 
.A(n_5186),
.Y(n_5432)
);

AOI22xp33_ASAP7_75t_SL g5433 ( 
.A1(n_5318),
.A2(n_5136),
.B1(n_4988),
.B2(n_5142),
.Y(n_5433)
);

CKINVDCx5p33_ASAP7_75t_R g5434 ( 
.A(n_5217),
.Y(n_5434)
);

AOI22xp33_ASAP7_75t_L g5435 ( 
.A1(n_5380),
.A2(n_5177),
.B1(n_5180),
.B2(n_5183),
.Y(n_5435)
);

AND2x4_ASAP7_75t_L g5436 ( 
.A(n_5348),
.B(n_5032),
.Y(n_5436)
);

CKINVDCx11_ASAP7_75t_R g5437 ( 
.A(n_5291),
.Y(n_5437)
);

OAI22xp33_ASAP7_75t_L g5438 ( 
.A1(n_5247),
.A2(n_5023),
.B1(n_5061),
.B2(n_5138),
.Y(n_5438)
);

AOI22xp33_ASAP7_75t_L g5439 ( 
.A1(n_5353),
.A2(n_5180),
.B1(n_4953),
.B2(n_4991),
.Y(n_5439)
);

INVx6_ASAP7_75t_L g5440 ( 
.A(n_5185),
.Y(n_5440)
);

CKINVDCx11_ASAP7_75t_R g5441 ( 
.A(n_5246),
.Y(n_5441)
);

OAI22xp33_ASAP7_75t_L g5442 ( 
.A1(n_5374),
.A2(n_5145),
.B1(n_5146),
.B2(n_5144),
.Y(n_5442)
);

BUFx2_ASAP7_75t_L g5443 ( 
.A(n_5309),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5254),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_5223),
.Y(n_5445)
);

AOI22xp33_ASAP7_75t_SL g5446 ( 
.A1(n_5381),
.A2(n_5398),
.B1(n_5242),
.B2(n_5300),
.Y(n_5446)
);

AOI22xp33_ASAP7_75t_L g5447 ( 
.A1(n_5344),
.A2(n_5123),
.B1(n_5031),
.B2(n_5082),
.Y(n_5447)
);

INVx2_ASAP7_75t_L g5448 ( 
.A(n_5239),
.Y(n_5448)
);

CKINVDCx5p33_ASAP7_75t_R g5449 ( 
.A(n_5275),
.Y(n_5449)
);

AOI22xp33_ASAP7_75t_L g5450 ( 
.A1(n_5202),
.A2(n_5001),
.B1(n_5003),
.B2(n_5002),
.Y(n_5450)
);

BUFx6f_ASAP7_75t_L g5451 ( 
.A(n_5221),
.Y(n_5451)
);

AOI22xp33_ASAP7_75t_SL g5452 ( 
.A1(n_5300),
.A2(n_5033),
.B1(n_4982),
.B2(n_4989),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5269),
.Y(n_5453)
);

INVx3_ASAP7_75t_L g5454 ( 
.A(n_5391),
.Y(n_5454)
);

INVx2_ASAP7_75t_L g5455 ( 
.A(n_5370),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_5276),
.Y(n_5456)
);

OAI22xp33_ASAP7_75t_L g5457 ( 
.A1(n_5261),
.A2(n_5088),
.B1(n_5076),
.B2(n_5120),
.Y(n_5457)
);

AOI22xp33_ASAP7_75t_SL g5458 ( 
.A1(n_5327),
.A2(n_5033),
.B1(n_4982),
.B2(n_4992),
.Y(n_5458)
);

AOI22xp5_ASAP7_75t_L g5459 ( 
.A1(n_5397),
.A2(n_4950),
.B1(n_5172),
.B2(n_5182),
.Y(n_5459)
);

OAI22xp5_ASAP7_75t_L g5460 ( 
.A1(n_5227),
.A2(n_5109),
.B1(n_5036),
.B2(n_5043),
.Y(n_5460)
);

INVx3_ASAP7_75t_L g5461 ( 
.A(n_5391),
.Y(n_5461)
);

AOI22xp33_ASAP7_75t_SL g5462 ( 
.A1(n_5327),
.A2(n_5033),
.B1(n_4982),
.B2(n_4993),
.Y(n_5462)
);

AOI22xp33_ASAP7_75t_L g5463 ( 
.A1(n_5315),
.A2(n_5028),
.B1(n_5046),
.B2(n_4998),
.Y(n_5463)
);

INVx8_ASAP7_75t_L g5464 ( 
.A(n_5361),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_5356),
.B(n_5363),
.Y(n_5465)
);

BUFx2_ASAP7_75t_L g5466 ( 
.A(n_5255),
.Y(n_5466)
);

AOI22xp5_ASAP7_75t_L g5467 ( 
.A1(n_5289),
.A2(n_5121),
.B1(n_5129),
.B2(n_5059),
.Y(n_5467)
);

BUFx6f_ASAP7_75t_L g5468 ( 
.A(n_5221),
.Y(n_5468)
);

AOI22xp5_ASAP7_75t_L g5469 ( 
.A1(n_5236),
.A2(n_5127),
.B1(n_5016),
.B2(n_4995),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_5277),
.Y(n_5470)
);

INVx6_ASAP7_75t_L g5471 ( 
.A(n_5259),
.Y(n_5471)
);

INVx2_ASAP7_75t_L g5472 ( 
.A(n_5384),
.Y(n_5472)
);

CKINVDCx20_ASAP7_75t_R g5473 ( 
.A(n_5333),
.Y(n_5473)
);

OAI22xp5_ASAP7_75t_L g5474 ( 
.A1(n_5228),
.A2(n_5151),
.B1(n_5139),
.B2(n_5091),
.Y(n_5474)
);

CKINVDCx11_ASAP7_75t_R g5475 ( 
.A(n_5366),
.Y(n_5475)
);

BUFx8_ASAP7_75t_SL g5476 ( 
.A(n_5366),
.Y(n_5476)
);

CKINVDCx11_ASAP7_75t_R g5477 ( 
.A(n_5362),
.Y(n_5477)
);

OAI22xp5_ASAP7_75t_L g5478 ( 
.A1(n_5219),
.A2(n_5151),
.B1(n_5139),
.B2(n_5091),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5279),
.Y(n_5479)
);

INVx2_ASAP7_75t_L g5480 ( 
.A(n_5306),
.Y(n_5480)
);

INVx1_ASAP7_75t_SL g5481 ( 
.A(n_5200),
.Y(n_5481)
);

AOI22xp33_ASAP7_75t_L g5482 ( 
.A1(n_5340),
.A2(n_2009),
.B1(n_2033),
.B2(n_2032),
.Y(n_5482)
);

CKINVDCx20_ASAP7_75t_R g5483 ( 
.A(n_5386),
.Y(n_5483)
);

INVx2_ASAP7_75t_SL g5484 ( 
.A(n_5190),
.Y(n_5484)
);

BUFx3_ASAP7_75t_L g5485 ( 
.A(n_5377),
.Y(n_5485)
);

INVx2_ASAP7_75t_SL g5486 ( 
.A(n_5197),
.Y(n_5486)
);

AND2x2_ASAP7_75t_L g5487 ( 
.A(n_5319),
.B(n_5084),
.Y(n_5487)
);

OAI22xp5_ASAP7_75t_L g5488 ( 
.A1(n_5345),
.A2(n_5151),
.B1(n_5139),
.B2(n_5091),
.Y(n_5488)
);

BUFx2_ASAP7_75t_L g5489 ( 
.A(n_5387),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5281),
.Y(n_5490)
);

AOI22xp33_ASAP7_75t_SL g5491 ( 
.A1(n_5250),
.A2(n_3343),
.B1(n_55),
.B2(n_57),
.Y(n_5491)
);

INVx3_ASAP7_75t_SL g5492 ( 
.A(n_5393),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5285),
.Y(n_5493)
);

AOI22xp33_ASAP7_75t_SL g5494 ( 
.A1(n_5265),
.A2(n_3343),
.B1(n_57),
.B2(n_58),
.Y(n_5494)
);

INVx11_ASAP7_75t_L g5495 ( 
.A(n_5194),
.Y(n_5495)
);

CKINVDCx11_ASAP7_75t_R g5496 ( 
.A(n_5271),
.Y(n_5496)
);

AOI22xp5_ASAP7_75t_L g5497 ( 
.A1(n_5265),
.A2(n_58),
.B1(n_59),
.B2(n_54),
.Y(n_5497)
);

CKINVDCx5p33_ASAP7_75t_R g5498 ( 
.A(n_5271),
.Y(n_5498)
);

INVx8_ASAP7_75t_L g5499 ( 
.A(n_5361),
.Y(n_5499)
);

CKINVDCx5p33_ASAP7_75t_R g5500 ( 
.A(n_5271),
.Y(n_5500)
);

CKINVDCx14_ASAP7_75t_R g5501 ( 
.A(n_5232),
.Y(n_5501)
);

CKINVDCx11_ASAP7_75t_R g5502 ( 
.A(n_5278),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5295),
.Y(n_5503)
);

BUFx2_ASAP7_75t_R g5504 ( 
.A(n_5245),
.Y(n_5504)
);

OAI22xp5_ASAP7_75t_SL g5505 ( 
.A1(n_5253),
.A2(n_32),
.B1(n_33),
.B2(n_60),
.Y(n_5505)
);

INVx4_ASAP7_75t_L g5506 ( 
.A(n_5253),
.Y(n_5506)
);

NAND2x1p5_ASAP7_75t_L g5507 ( 
.A(n_5324),
.B(n_5084),
.Y(n_5507)
);

INVx6_ASAP7_75t_L g5508 ( 
.A(n_5278),
.Y(n_5508)
);

INVx2_ASAP7_75t_L g5509 ( 
.A(n_5286),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_5305),
.Y(n_5510)
);

CKINVDCx6p67_ASAP7_75t_R g5511 ( 
.A(n_5233),
.Y(n_5511)
);

BUFx4_ASAP7_75t_SL g5512 ( 
.A(n_5252),
.Y(n_5512)
);

INVx1_ASAP7_75t_SL g5513 ( 
.A(n_5368),
.Y(n_5513)
);

OAI22xp5_ASAP7_75t_L g5514 ( 
.A1(n_5218),
.A2(n_2919),
.B1(n_2927),
.B2(n_2920),
.Y(n_5514)
);

CKINVDCx5p33_ASAP7_75t_R g5515 ( 
.A(n_5278),
.Y(n_5515)
);

INVx2_ASAP7_75t_L g5516 ( 
.A(n_5305),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_5367),
.B(n_60),
.Y(n_5517)
);

CKINVDCx11_ASAP7_75t_R g5518 ( 
.A(n_5282),
.Y(n_5518)
);

AOI22xp33_ASAP7_75t_L g5519 ( 
.A1(n_5376),
.A2(n_2009),
.B1(n_2033),
.B2(n_2032),
.Y(n_5519)
);

AOI22xp33_ASAP7_75t_SL g5520 ( 
.A1(n_5237),
.A2(n_62),
.B1(n_63),
.B2(n_61),
.Y(n_5520)
);

INVx6_ASAP7_75t_L g5521 ( 
.A(n_5296),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_5304),
.Y(n_5522)
);

CKINVDCx5p33_ASAP7_75t_R g5523 ( 
.A(n_5296),
.Y(n_5523)
);

AOI22xp33_ASAP7_75t_L g5524 ( 
.A1(n_5339),
.A2(n_5352),
.B1(n_5240),
.B2(n_5357),
.Y(n_5524)
);

AOI21xp5_ASAP7_75t_L g5525 ( 
.A1(n_5225),
.A2(n_2042),
.B(n_1960),
.Y(n_5525)
);

BUFx3_ASAP7_75t_L g5526 ( 
.A(n_5396),
.Y(n_5526)
);

AOI21xp5_ASAP7_75t_L g5527 ( 
.A1(n_5331),
.A2(n_2042),
.B(n_1960),
.Y(n_5527)
);

INVx6_ASAP7_75t_L g5528 ( 
.A(n_5296),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_5313),
.Y(n_5529)
);

CKINVDCx20_ASAP7_75t_R g5530 ( 
.A(n_5199),
.Y(n_5530)
);

OAI22xp5_ASAP7_75t_L g5531 ( 
.A1(n_5329),
.A2(n_2919),
.B1(n_2927),
.B2(n_2920),
.Y(n_5531)
);

OAI22xp33_ASAP7_75t_SL g5532 ( 
.A1(n_5266),
.A2(n_33),
.B1(n_62),
.B2(n_61),
.Y(n_5532)
);

BUFx3_ASAP7_75t_L g5533 ( 
.A(n_5294),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5321),
.Y(n_5534)
);

AOI22xp5_ASAP7_75t_L g5535 ( 
.A1(n_5394),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_5328),
.Y(n_5536)
);

INVx2_ASAP7_75t_L g5537 ( 
.A(n_5326),
.Y(n_5537)
);

AOI22xp5_ASAP7_75t_L g5538 ( 
.A1(n_5268),
.A2(n_70),
.B1(n_64),
.B2(n_69),
.Y(n_5538)
);

NAND2xp5_ASAP7_75t_L g5539 ( 
.A(n_5215),
.B(n_70),
.Y(n_5539)
);

INVx2_ASAP7_75t_L g5540 ( 
.A(n_5326),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5330),
.Y(n_5541)
);

AND2x2_ASAP7_75t_L g5542 ( 
.A(n_5189),
.B(n_72),
.Y(n_5542)
);

AOI22xp33_ASAP7_75t_L g5543 ( 
.A1(n_5270),
.A2(n_2035),
.B1(n_2044),
.B2(n_2039),
.Y(n_5543)
);

CKINVDCx12_ASAP7_75t_R g5544 ( 
.A(n_5292),
.Y(n_5544)
);

OAI22xp5_ASAP7_75t_L g5545 ( 
.A1(n_5329),
.A2(n_2939),
.B1(n_2940),
.B2(n_2931),
.Y(n_5545)
);

CKINVDCx11_ASAP7_75t_R g5546 ( 
.A(n_5303),
.Y(n_5546)
);

AOI22xp33_ASAP7_75t_L g5547 ( 
.A1(n_5355),
.A2(n_2035),
.B1(n_2044),
.B2(n_2039),
.Y(n_5547)
);

BUFx12f_ASAP7_75t_L g5548 ( 
.A(n_5342),
.Y(n_5548)
);

AOI22xp33_ASAP7_75t_L g5549 ( 
.A1(n_5205),
.A2(n_2035),
.B1(n_2044),
.B2(n_2039),
.Y(n_5549)
);

BUFx6f_ASAP7_75t_L g5550 ( 
.A(n_5303),
.Y(n_5550)
);

INVx2_ASAP7_75t_SL g5551 ( 
.A(n_5189),
.Y(n_5551)
);

CKINVDCx14_ASAP7_75t_R g5552 ( 
.A(n_5263),
.Y(n_5552)
);

BUFx3_ASAP7_75t_L g5553 ( 
.A(n_5343),
.Y(n_5553)
);

OAI22xp33_ASAP7_75t_L g5554 ( 
.A1(n_5324),
.A2(n_5212),
.B1(n_5204),
.B2(n_5213),
.Y(n_5554)
);

BUFx3_ASAP7_75t_L g5555 ( 
.A(n_5268),
.Y(n_5555)
);

OAI22xp33_ASAP7_75t_L g5556 ( 
.A1(n_5216),
.A2(n_77),
.B1(n_74),
.B2(n_75),
.Y(n_5556)
);

INVx2_ASAP7_75t_L g5557 ( 
.A(n_5244),
.Y(n_5557)
);

BUFx10_ASAP7_75t_L g5558 ( 
.A(n_5280),
.Y(n_5558)
);

CKINVDCx5p33_ASAP7_75t_R g5559 ( 
.A(n_5323),
.Y(n_5559)
);

INVx6_ASAP7_75t_L g5560 ( 
.A(n_5323),
.Y(n_5560)
);

AOI22xp33_ASAP7_75t_L g5561 ( 
.A1(n_5196),
.A2(n_2064),
.B1(n_2067),
.B2(n_2047),
.Y(n_5561)
);

AOI22xp33_ASAP7_75t_SL g5562 ( 
.A1(n_5243),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_5562)
);

INVxp67_ASAP7_75t_SL g5563 ( 
.A(n_5392),
.Y(n_5563)
);

AOI22xp33_ASAP7_75t_SL g5564 ( 
.A1(n_5399),
.A2(n_84),
.B1(n_80),
.B2(n_82),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_5203),
.B(n_84),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_5298),
.Y(n_5566)
);

CKINVDCx20_ASAP7_75t_R g5567 ( 
.A(n_5365),
.Y(n_5567)
);

AND2x2_ASAP7_75t_L g5568 ( 
.A(n_5287),
.B(n_85),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_5288),
.Y(n_5569)
);

BUFx12f_ASAP7_75t_L g5570 ( 
.A(n_5311),
.Y(n_5570)
);

INVx6_ASAP7_75t_L g5571 ( 
.A(n_5346),
.Y(n_5571)
);

INVx2_ASAP7_75t_SL g5572 ( 
.A(n_5226),
.Y(n_5572)
);

HB1xp67_ASAP7_75t_L g5573 ( 
.A(n_5385),
.Y(n_5573)
);

AOI22xp33_ASAP7_75t_SL g5574 ( 
.A1(n_5280),
.A2(n_89),
.B1(n_86),
.B2(n_87),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5378),
.Y(n_5575)
);

BUFx3_ASAP7_75t_L g5576 ( 
.A(n_5290),
.Y(n_5576)
);

CKINVDCx5p33_ASAP7_75t_R g5577 ( 
.A(n_5346),
.Y(n_5577)
);

INVx6_ASAP7_75t_L g5578 ( 
.A(n_5346),
.Y(n_5578)
);

CKINVDCx11_ASAP7_75t_R g5579 ( 
.A(n_5358),
.Y(n_5579)
);

AOI22xp5_ASAP7_75t_SL g5580 ( 
.A1(n_5290),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5388),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_5395),
.Y(n_5582)
);

BUFx12f_ASAP7_75t_L g5583 ( 
.A(n_5238),
.Y(n_5583)
);

AOI22xp5_ASAP7_75t_L g5584 ( 
.A1(n_5383),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_5584)
);

AOI22xp33_ASAP7_75t_L g5585 ( 
.A1(n_5230),
.A2(n_2064),
.B1(n_2067),
.B2(n_2047),
.Y(n_5585)
);

NOR2xp33_ASAP7_75t_L g5586 ( 
.A(n_5412),
.B(n_5241),
.Y(n_5586)
);

NAND2xp5_ASAP7_75t_L g5587 ( 
.A(n_5421),
.B(n_5322),
.Y(n_5587)
);

CKINVDCx8_ASAP7_75t_R g5588 ( 
.A(n_5451),
.Y(n_5588)
);

OAI22xp33_ASAP7_75t_L g5589 ( 
.A1(n_5492),
.A2(n_5382),
.B1(n_5224),
.B2(n_5360),
.Y(n_5589)
);

AOI22xp33_ASAP7_75t_L g5590 ( 
.A1(n_5405),
.A2(n_5201),
.B1(n_5272),
.B2(n_5351),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5400),
.Y(n_5591)
);

AND2x4_ASAP7_75t_L g5592 ( 
.A(n_5411),
.B(n_5337),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_5446),
.B(n_5293),
.Y(n_5593)
);

AOI22xp33_ASAP7_75t_L g5594 ( 
.A1(n_5427),
.A2(n_5214),
.B1(n_5206),
.B2(n_5301),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5414),
.Y(n_5595)
);

CKINVDCx16_ASAP7_75t_R g5596 ( 
.A(n_5473),
.Y(n_5596)
);

AO31x2_ASAP7_75t_L g5597 ( 
.A1(n_5506),
.A2(n_5314),
.A3(n_5336),
.B(n_5332),
.Y(n_5597)
);

BUFx12f_ASAP7_75t_L g5598 ( 
.A(n_5437),
.Y(n_5598)
);

AOI21xp33_ASAP7_75t_L g5599 ( 
.A1(n_5554),
.A2(n_5338),
.B(n_5369),
.Y(n_5599)
);

OAI21x1_ASAP7_75t_L g5600 ( 
.A1(n_5420),
.A2(n_5371),
.B(n_5359),
.Y(n_5600)
);

OAI22xp33_ASAP7_75t_L g5601 ( 
.A1(n_5443),
.A2(n_5360),
.B1(n_5262),
.B2(n_5283),
.Y(n_5601)
);

AOI21xp33_ASAP7_75t_L g5602 ( 
.A1(n_5442),
.A2(n_5372),
.B(n_5251),
.Y(n_5602)
);

OR2x2_ASAP7_75t_L g5603 ( 
.A(n_5445),
.B(n_5220),
.Y(n_5603)
);

AOI21xp33_ASAP7_75t_L g5604 ( 
.A1(n_5438),
.A2(n_5406),
.B(n_5423),
.Y(n_5604)
);

BUFx2_ASAP7_75t_L g5605 ( 
.A(n_5501),
.Y(n_5605)
);

NAND2x1_ASAP7_75t_L g5606 ( 
.A(n_5466),
.B(n_5359),
.Y(n_5606)
);

BUFx8_ASAP7_75t_L g5607 ( 
.A(n_5451),
.Y(n_5607)
);

NAND2xp5_ASAP7_75t_SL g5608 ( 
.A(n_5433),
.B(n_5425),
.Y(n_5608)
);

CKINVDCx16_ASAP7_75t_R g5609 ( 
.A(n_5407),
.Y(n_5609)
);

INVx2_ASAP7_75t_SL g5610 ( 
.A(n_5558),
.Y(n_5610)
);

AOI22xp33_ASAP7_75t_SL g5611 ( 
.A1(n_5505),
.A2(n_5264),
.B1(n_5262),
.B2(n_5347),
.Y(n_5611)
);

OAI22xp33_ASAP7_75t_L g5612 ( 
.A1(n_5511),
.A2(n_5325),
.B1(n_5334),
.B2(n_5308),
.Y(n_5612)
);

CKINVDCx5p33_ASAP7_75t_R g5613 ( 
.A(n_5441),
.Y(n_5613)
);

INVx4_ASAP7_75t_L g5614 ( 
.A(n_5451),
.Y(n_5614)
);

AND2x6_ASAP7_75t_L g5615 ( 
.A(n_5468),
.B(n_5391),
.Y(n_5615)
);

AND2x6_ASAP7_75t_L g5616 ( 
.A(n_5468),
.B(n_5358),
.Y(n_5616)
);

INVx3_ASAP7_75t_L g5617 ( 
.A(n_5403),
.Y(n_5617)
);

OAI22xp5_ASAP7_75t_L g5618 ( 
.A1(n_5413),
.A2(n_5422),
.B1(n_5401),
.B2(n_5504),
.Y(n_5618)
);

AND2x2_ASAP7_75t_L g5619 ( 
.A(n_5489),
.B(n_5371),
.Y(n_5619)
);

HB1xp67_ASAP7_75t_L g5620 ( 
.A(n_5448),
.Y(n_5620)
);

INVx3_ASAP7_75t_L g5621 ( 
.A(n_5403),
.Y(n_5621)
);

CKINVDCx5p33_ASAP7_75t_R g5622 ( 
.A(n_5449),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_5444),
.Y(n_5623)
);

INVx2_ASAP7_75t_SL g5624 ( 
.A(n_5558),
.Y(n_5624)
);

AOI22xp33_ASAP7_75t_SL g5625 ( 
.A1(n_5505),
.A2(n_5350),
.B1(n_5335),
.B2(n_5211),
.Y(n_5625)
);

BUFx3_ASAP7_75t_L g5626 ( 
.A(n_5476),
.Y(n_5626)
);

CKINVDCx6p67_ASAP7_75t_R g5627 ( 
.A(n_5477),
.Y(n_5627)
);

OR2x2_ASAP7_75t_L g5628 ( 
.A(n_5486),
.B(n_5302),
.Y(n_5628)
);

AND2x4_ASAP7_75t_L g5629 ( 
.A(n_5506),
.B(n_5341),
.Y(n_5629)
);

INVx4_ASAP7_75t_SL g5630 ( 
.A(n_5410),
.Y(n_5630)
);

INVx6_ASAP7_75t_L g5631 ( 
.A(n_5468),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_5453),
.Y(n_5632)
);

INVx1_ASAP7_75t_SL g5633 ( 
.A(n_5475),
.Y(n_5633)
);

BUFx4f_ASAP7_75t_L g5634 ( 
.A(n_5410),
.Y(n_5634)
);

OR2x6_ASAP7_75t_L g5635 ( 
.A(n_5424),
.B(n_5299),
.Y(n_5635)
);

NAND2xp5_ASAP7_75t_L g5636 ( 
.A(n_5465),
.B(n_5310),
.Y(n_5636)
);

OAI22xp33_ASAP7_75t_L g5637 ( 
.A1(n_5481),
.A2(n_5430),
.B1(n_5459),
.B2(n_5513),
.Y(n_5637)
);

NAND2xp5_ASAP7_75t_L g5638 ( 
.A(n_5517),
.B(n_5214),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5456),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_5470),
.Y(n_5640)
);

OA21x2_ASAP7_75t_L g5641 ( 
.A1(n_5563),
.A2(n_5426),
.B(n_5569),
.Y(n_5641)
);

INVx2_ASAP7_75t_SL g5642 ( 
.A(n_5424),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_5479),
.Y(n_5643)
);

NAND2xp5_ASAP7_75t_L g5644 ( 
.A(n_5524),
.B(n_5335),
.Y(n_5644)
);

BUFx2_ASAP7_75t_L g5645 ( 
.A(n_5567),
.Y(n_5645)
);

CKINVDCx16_ASAP7_75t_R g5646 ( 
.A(n_5485),
.Y(n_5646)
);

NAND2xp5_ASAP7_75t_L g5647 ( 
.A(n_5566),
.B(n_5358),
.Y(n_5647)
);

OAI22xp33_ASAP7_75t_L g5648 ( 
.A1(n_5459),
.A2(n_5307),
.B1(n_5211),
.B2(n_5274),
.Y(n_5648)
);

AO21x2_ASAP7_75t_L g5649 ( 
.A1(n_5415),
.A2(n_5297),
.B(n_5231),
.Y(n_5649)
);

AOI22xp33_ASAP7_75t_L g5650 ( 
.A1(n_5418),
.A2(n_5256),
.B1(n_5320),
.B2(n_5229),
.Y(n_5650)
);

OAI22xp5_ASAP7_75t_L g5651 ( 
.A1(n_5404),
.A2(n_5375),
.B1(n_5379),
.B2(n_5207),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_5490),
.Y(n_5652)
);

NOR2xp33_ASAP7_75t_L g5653 ( 
.A(n_5495),
.B(n_92),
.Y(n_5653)
);

AND2x2_ASAP7_75t_L g5654 ( 
.A(n_5572),
.B(n_5249),
.Y(n_5654)
);

AO31x2_ASAP7_75t_L g5655 ( 
.A1(n_5575),
.A2(n_5284),
.A3(n_5249),
.B(n_98),
.Y(n_5655)
);

A2O1A1Ixp33_ASAP7_75t_L g5656 ( 
.A1(n_5580),
.A2(n_98),
.B(n_93),
.C(n_97),
.Y(n_5656)
);

OA21x2_ASAP7_75t_L g5657 ( 
.A1(n_5581),
.A2(n_5582),
.B(n_5472),
.Y(n_5657)
);

OAI22xp5_ASAP7_75t_L g5658 ( 
.A1(n_5431),
.A2(n_5249),
.B1(n_102),
.B2(n_99),
.Y(n_5658)
);

BUFx6f_ASAP7_75t_L g5659 ( 
.A(n_5496),
.Y(n_5659)
);

OAI22xp5_ASAP7_75t_L g5660 ( 
.A1(n_5552),
.A2(n_102),
.B1(n_99),
.B2(n_101),
.Y(n_5660)
);

OAI22xp5_ASAP7_75t_L g5661 ( 
.A1(n_5409),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_5661)
);

OR2x6_ASAP7_75t_L g5662 ( 
.A(n_5428),
.B(n_1221),
.Y(n_5662)
);

NAND2xp33_ASAP7_75t_R g5663 ( 
.A(n_5434),
.B(n_106),
.Y(n_5663)
);

AND2x2_ASAP7_75t_L g5664 ( 
.A(n_5480),
.B(n_108),
.Y(n_5664)
);

OAI22xp5_ASAP7_75t_L g5665 ( 
.A1(n_5452),
.A2(n_114),
.B1(n_108),
.B2(n_113),
.Y(n_5665)
);

OAI22xp5_ASAP7_75t_L g5666 ( 
.A1(n_5564),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_5503),
.Y(n_5667)
);

OAI22xp5_ASAP7_75t_L g5668 ( 
.A1(n_5458),
.A2(n_118),
.B1(n_115),
.B2(n_116),
.Y(n_5668)
);

BUFx3_ASAP7_75t_L g5669 ( 
.A(n_5483),
.Y(n_5669)
);

AND2x2_ASAP7_75t_L g5670 ( 
.A(n_5551),
.B(n_119),
.Y(n_5670)
);

OAI22xp5_ASAP7_75t_L g5671 ( 
.A1(n_5535),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_5671)
);

AOI21xp33_ASAP7_75t_L g5672 ( 
.A1(n_5450),
.A2(n_120),
.B(n_122),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5522),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_5529),
.Y(n_5674)
);

AOI22xp33_ASAP7_75t_SL g5675 ( 
.A1(n_5580),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5534),
.Y(n_5676)
);

INVx3_ASAP7_75t_L g5677 ( 
.A(n_5440),
.Y(n_5677)
);

OAI211xp5_ASAP7_75t_L g5678 ( 
.A1(n_5520),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_5678)
);

OAI22xp33_ASAP7_75t_L g5679 ( 
.A1(n_5535),
.A2(n_5484),
.B1(n_5584),
.B2(n_5497),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5536),
.Y(n_5680)
);

INVx3_ASAP7_75t_L g5681 ( 
.A(n_5440),
.Y(n_5681)
);

OAI22xp33_ASAP7_75t_L g5682 ( 
.A1(n_5584),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_5682)
);

NAND2xp33_ASAP7_75t_R g5683 ( 
.A(n_5498),
.B(n_129),
.Y(n_5683)
);

OAI21x1_ASAP7_75t_SL g5684 ( 
.A1(n_5432),
.A2(n_130),
.B(n_131),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_5541),
.Y(n_5685)
);

INVx3_ASAP7_75t_L g5686 ( 
.A(n_5550),
.Y(n_5686)
);

AND2x4_ASAP7_75t_L g5687 ( 
.A(n_5436),
.B(n_132),
.Y(n_5687)
);

AO31x2_ASAP7_75t_L g5688 ( 
.A1(n_5455),
.A2(n_134),
.A3(n_130),
.B(n_132),
.Y(n_5688)
);

O2A1O1Ixp33_ASAP7_75t_SL g5689 ( 
.A1(n_5408),
.A2(n_137),
.B(n_139),
.C(n_136),
.Y(n_5689)
);

OAI22xp5_ASAP7_75t_L g5690 ( 
.A1(n_5491),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_5690)
);

OR2x6_ASAP7_75t_L g5691 ( 
.A(n_5428),
.B(n_1221),
.Y(n_5691)
);

NAND2xp5_ASAP7_75t_L g5692 ( 
.A(n_5565),
.B(n_135),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_5550),
.Y(n_5693)
);

AND2x2_ASAP7_75t_L g5694 ( 
.A(n_5454),
.B(n_140),
.Y(n_5694)
);

OAI22xp5_ASAP7_75t_L g5695 ( 
.A1(n_5462),
.A2(n_144),
.B1(n_141),
.B2(n_142),
.Y(n_5695)
);

OAI222xp33_ASAP7_75t_L g5696 ( 
.A1(n_5538),
.A2(n_145),
.B1(n_147),
.B2(n_141),
.C1(n_142),
.C2(n_146),
.Y(n_5696)
);

AOI22xp33_ASAP7_75t_L g5697 ( 
.A1(n_5583),
.A2(n_2064),
.B1(n_2067),
.B2(n_2047),
.Y(n_5697)
);

INVxp67_ASAP7_75t_SL g5698 ( 
.A(n_5416),
.Y(n_5698)
);

CKINVDCx11_ASAP7_75t_R g5699 ( 
.A(n_5402),
.Y(n_5699)
);

AOI21xp33_ASAP7_75t_L g5700 ( 
.A1(n_5556),
.A2(n_145),
.B(n_146),
.Y(n_5700)
);

OAI22xp33_ASAP7_75t_L g5701 ( 
.A1(n_5497),
.A2(n_5555),
.B1(n_5576),
.B2(n_5538),
.Y(n_5701)
);

OAI21x1_ASAP7_75t_L g5702 ( 
.A1(n_5507),
.A2(n_2955),
.B(n_2952),
.Y(n_5702)
);

AOI21xp33_ASAP7_75t_L g5703 ( 
.A1(n_5532),
.A2(n_148),
.B(n_149),
.Y(n_5703)
);

INVx4_ASAP7_75t_L g5704 ( 
.A(n_5428),
.Y(n_5704)
);

BUFx2_ASAP7_75t_L g5705 ( 
.A(n_5419),
.Y(n_5705)
);

BUFx3_ASAP7_75t_L g5706 ( 
.A(n_5570),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5487),
.Y(n_5707)
);

BUFx3_ASAP7_75t_L g5708 ( 
.A(n_5526),
.Y(n_5708)
);

AOI22xp33_ASAP7_75t_L g5709 ( 
.A1(n_5562),
.A2(n_2090),
.B1(n_2099),
.B2(n_2068),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_5573),
.Y(n_5710)
);

INVx2_ASAP7_75t_L g5711 ( 
.A(n_5471),
.Y(n_5711)
);

CKINVDCx5p33_ASAP7_75t_R g5712 ( 
.A(n_5502),
.Y(n_5712)
);

CKINVDCx20_ASAP7_75t_R g5713 ( 
.A(n_5530),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5454),
.B(n_5461),
.Y(n_5714)
);

OAI22xp5_ASAP7_75t_L g5715 ( 
.A1(n_5547),
.A2(n_152),
.B1(n_149),
.B2(n_151),
.Y(n_5715)
);

BUFx3_ASAP7_75t_L g5716 ( 
.A(n_5429),
.Y(n_5716)
);

A2O1A1Ixp33_ASAP7_75t_L g5717 ( 
.A1(n_5574),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_5717)
);

NOR4xp25_ASAP7_75t_L g5718 ( 
.A(n_5539),
.B(n_158),
.C(n_156),
.D(n_157),
.Y(n_5718)
);

AND2x4_ASAP7_75t_L g5719 ( 
.A(n_5461),
.B(n_159),
.Y(n_5719)
);

INVx2_ASAP7_75t_L g5720 ( 
.A(n_5471),
.Y(n_5720)
);

AOI221xp5_ASAP7_75t_L g5721 ( 
.A1(n_5494),
.A2(n_5460),
.B1(n_5447),
.B2(n_5568),
.C(n_5585),
.Y(n_5721)
);

OAI22xp5_ASAP7_75t_L g5722 ( 
.A1(n_5500),
.A2(n_5523),
.B1(n_5559),
.B2(n_5515),
.Y(n_5722)
);

AO21x2_ASAP7_75t_L g5723 ( 
.A1(n_5493),
.A2(n_158),
.B(n_159),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5557),
.Y(n_5724)
);

CKINVDCx5p33_ASAP7_75t_R g5725 ( 
.A(n_5518),
.Y(n_5725)
);

BUFx3_ASAP7_75t_L g5726 ( 
.A(n_5546),
.Y(n_5726)
);

AND2x2_ASAP7_75t_L g5727 ( 
.A(n_5533),
.B(n_161),
.Y(n_5727)
);

AND2x2_ASAP7_75t_L g5728 ( 
.A(n_5553),
.B(n_162),
.Y(n_5728)
);

AOI21xp33_ASAP7_75t_L g5729 ( 
.A1(n_5439),
.A2(n_162),
.B(n_163),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_5508),
.Y(n_5730)
);

NAND2xp5_ASAP7_75t_L g5731 ( 
.A(n_5542),
.B(n_164),
.Y(n_5731)
);

INVx1_ASAP7_75t_SL g5732 ( 
.A(n_5579),
.Y(n_5732)
);

NOR2xp33_ASAP7_75t_L g5733 ( 
.A(n_5548),
.B(n_165),
.Y(n_5733)
);

BUFx2_ASAP7_75t_L g5734 ( 
.A(n_5464),
.Y(n_5734)
);

AOI22xp33_ASAP7_75t_L g5735 ( 
.A1(n_5464),
.A2(n_2140),
.B1(n_2100),
.B2(n_2042),
.Y(n_5735)
);

OAI21x1_ASAP7_75t_L g5736 ( 
.A1(n_5509),
.A2(n_3010),
.B(n_3008),
.Y(n_5736)
);

NAND2xp5_ASAP7_75t_L g5737 ( 
.A(n_5510),
.B(n_166),
.Y(n_5737)
);

NAND2x1_ASAP7_75t_L g5738 ( 
.A(n_5417),
.B(n_1221),
.Y(n_5738)
);

AOI21xp5_ASAP7_75t_L g5739 ( 
.A1(n_5464),
.A2(n_166),
.B(n_167),
.Y(n_5739)
);

AND2x4_ASAP7_75t_L g5740 ( 
.A(n_5516),
.B(n_168),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5508),
.Y(n_5741)
);

AND2x2_ASAP7_75t_L g5742 ( 
.A(n_5537),
.B(n_167),
.Y(n_5742)
);

OAI21x1_ASAP7_75t_L g5743 ( 
.A1(n_5540),
.A2(n_3019),
.B(n_3017),
.Y(n_5743)
);

OAI22xp5_ASAP7_75t_L g5744 ( 
.A1(n_5577),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_5744)
);

AOI22xp33_ASAP7_75t_L g5745 ( 
.A1(n_5499),
.A2(n_2100),
.B1(n_2140),
.B2(n_1960),
.Y(n_5745)
);

AOI22xp33_ASAP7_75t_L g5746 ( 
.A1(n_5499),
.A2(n_2140),
.B1(n_2100),
.B2(n_2678),
.Y(n_5746)
);

AND2x6_ASAP7_75t_L g5747 ( 
.A(n_5467),
.B(n_170),
.Y(n_5747)
);

NAND2xp33_ASAP7_75t_R g5748 ( 
.A(n_5512),
.B(n_171),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5521),
.Y(n_5749)
);

AND2x4_ASAP7_75t_L g5750 ( 
.A(n_5463),
.B(n_174),
.Y(n_5750)
);

OAI22xp33_ASAP7_75t_L g5751 ( 
.A1(n_5528),
.A2(n_176),
.B1(n_173),
.B2(n_175),
.Y(n_5751)
);

INVx3_ASAP7_75t_L g5752 ( 
.A(n_5560),
.Y(n_5752)
);

AND2x6_ASAP7_75t_SL g5753 ( 
.A(n_5544),
.B(n_175),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5560),
.Y(n_5754)
);

BUFx12f_ASAP7_75t_L g5755 ( 
.A(n_5578),
.Y(n_5755)
);

INVx6_ASAP7_75t_L g5756 ( 
.A(n_5571),
.Y(n_5756)
);

AOI22xp33_ASAP7_75t_L g5757 ( 
.A1(n_5578),
.A2(n_2713),
.B1(n_2741),
.B2(n_2694),
.Y(n_5757)
);

OR2x6_ASAP7_75t_L g5758 ( 
.A(n_5527),
.B(n_1270),
.Y(n_5758)
);

AOI22xp33_ASAP7_75t_L g5759 ( 
.A1(n_5549),
.A2(n_2741),
.B1(n_2744),
.B2(n_2713),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5474),
.Y(n_5760)
);

OAI221xp5_ASAP7_75t_L g5761 ( 
.A1(n_5435),
.A2(n_182),
.B1(n_178),
.B2(n_181),
.C(n_183),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5705),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5591),
.Y(n_5763)
);

AOI211xp5_ASAP7_75t_L g5764 ( 
.A1(n_5618),
.A2(n_5457),
.B(n_5478),
.C(n_5488),
.Y(n_5764)
);

INVx5_ASAP7_75t_L g5765 ( 
.A(n_5598),
.Y(n_5765)
);

AND2x2_ASAP7_75t_L g5766 ( 
.A(n_5605),
.B(n_5561),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5595),
.Y(n_5767)
);

OAI21xp5_ASAP7_75t_SL g5768 ( 
.A1(n_5701),
.A2(n_5482),
.B(n_5543),
.Y(n_5768)
);

AOI22xp33_ASAP7_75t_L g5769 ( 
.A1(n_5747),
.A2(n_5519),
.B1(n_5469),
.B2(n_5514),
.Y(n_5769)
);

INVxp67_ASAP7_75t_L g5770 ( 
.A(n_5748),
.Y(n_5770)
);

OAI21xp5_ASAP7_75t_SL g5771 ( 
.A1(n_5604),
.A2(n_5545),
.B(n_5531),
.Y(n_5771)
);

NOR2xp33_ASAP7_75t_L g5772 ( 
.A(n_5627),
.B(n_182),
.Y(n_5772)
);

AOI22xp33_ASAP7_75t_L g5773 ( 
.A1(n_5747),
.A2(n_5525),
.B1(n_2741),
.B2(n_2744),
.Y(n_5773)
);

AOI22xp33_ASAP7_75t_L g5774 ( 
.A1(n_5747),
.A2(n_2744),
.B1(n_2750),
.B2(n_2713),
.Y(n_5774)
);

OAI21xp5_ASAP7_75t_L g5775 ( 
.A1(n_5739),
.A2(n_183),
.B(n_185),
.Y(n_5775)
);

INVx5_ASAP7_75t_SL g5776 ( 
.A(n_5659),
.Y(n_5776)
);

NAND2xp5_ASAP7_75t_L g5777 ( 
.A(n_5687),
.B(n_187),
.Y(n_5777)
);

INVx2_ASAP7_75t_L g5778 ( 
.A(n_5631),
.Y(n_5778)
);

OAI22xp5_ASAP7_75t_L g5779 ( 
.A1(n_5594),
.A2(n_191),
.B1(n_188),
.B2(n_189),
.Y(n_5779)
);

OAI22xp5_ASAP7_75t_L g5780 ( 
.A1(n_5611),
.A2(n_192),
.B1(n_188),
.B2(n_189),
.Y(n_5780)
);

AOI22xp33_ASAP7_75t_L g5781 ( 
.A1(n_5608),
.A2(n_2757),
.B1(n_2750),
.B2(n_1288),
.Y(n_5781)
);

CKINVDCx20_ASAP7_75t_R g5782 ( 
.A(n_5713),
.Y(n_5782)
);

HB1xp67_ASAP7_75t_L g5783 ( 
.A(n_5620),
.Y(n_5783)
);

OAI22xp5_ASAP7_75t_SL g5784 ( 
.A1(n_5646),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_5784)
);

AOI22xp33_ASAP7_75t_L g5785 ( 
.A1(n_5679),
.A2(n_2757),
.B1(n_2750),
.B2(n_1288),
.Y(n_5785)
);

OAI21xp5_ASAP7_75t_SL g5786 ( 
.A1(n_5675),
.A2(n_193),
.B(n_194),
.Y(n_5786)
);

OAI22xp5_ASAP7_75t_L g5787 ( 
.A1(n_5650),
.A2(n_198),
.B1(n_195),
.B2(n_196),
.Y(n_5787)
);

OAI22xp33_ASAP7_75t_L g5788 ( 
.A1(n_5593),
.A2(n_199),
.B1(n_195),
.B2(n_198),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5631),
.Y(n_5789)
);

OAI22xp5_ASAP7_75t_L g5790 ( 
.A1(n_5625),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_5790)
);

NOR2xp33_ASAP7_75t_L g5791 ( 
.A(n_5609),
.B(n_203),
.Y(n_5791)
);

INVx5_ASAP7_75t_SL g5792 ( 
.A(n_5659),
.Y(n_5792)
);

AND2x2_ASAP7_75t_L g5793 ( 
.A(n_5752),
.B(n_203),
.Y(n_5793)
);

NAND2x1p5_ASAP7_75t_L g5794 ( 
.A(n_5606),
.B(n_1289),
.Y(n_5794)
);

HB1xp67_ASAP7_75t_L g5795 ( 
.A(n_5597),
.Y(n_5795)
);

OR2x2_ASAP7_75t_SL g5796 ( 
.A(n_5596),
.B(n_208),
.Y(n_5796)
);

AOI22xp33_ASAP7_75t_L g5797 ( 
.A1(n_5760),
.A2(n_1289),
.B1(n_1318),
.B2(n_1307),
.Y(n_5797)
);

AOI22xp33_ASAP7_75t_L g5798 ( 
.A1(n_5637),
.A2(n_1289),
.B1(n_1318),
.B2(n_1307),
.Y(n_5798)
);

AND2x2_ASAP7_75t_L g5799 ( 
.A(n_5714),
.B(n_210),
.Y(n_5799)
);

OAI21xp5_ASAP7_75t_L g5800 ( 
.A1(n_5656),
.A2(n_211),
.B(n_214),
.Y(n_5800)
);

AOI22xp33_ASAP7_75t_L g5801 ( 
.A1(n_5672),
.A2(n_5721),
.B1(n_5729),
.B2(n_5658),
.Y(n_5801)
);

AOI22xp33_ASAP7_75t_L g5802 ( 
.A1(n_5750),
.A2(n_1318),
.B1(n_1338),
.B2(n_1325),
.Y(n_5802)
);

AOI22xp33_ASAP7_75t_L g5803 ( 
.A1(n_5750),
.A2(n_1325),
.B1(n_1354),
.B2(n_1338),
.Y(n_5803)
);

AOI21xp5_ASAP7_75t_L g5804 ( 
.A1(n_5668),
.A2(n_211),
.B(n_214),
.Y(n_5804)
);

OAI22xp33_ASAP7_75t_L g5805 ( 
.A1(n_5683),
.A2(n_218),
.B1(n_215),
.B2(n_216),
.Y(n_5805)
);

AOI22xp33_ASAP7_75t_L g5806 ( 
.A1(n_5695),
.A2(n_1325),
.B1(n_1354),
.B2(n_1338),
.Y(n_5806)
);

OAI22xp33_ASAP7_75t_L g5807 ( 
.A1(n_5663),
.A2(n_218),
.B1(n_215),
.B2(n_216),
.Y(n_5807)
);

AOI22xp33_ASAP7_75t_L g5808 ( 
.A1(n_5665),
.A2(n_1325),
.B1(n_1354),
.B2(n_1338),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5756),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5623),
.Y(n_5810)
);

CKINVDCx6p67_ASAP7_75t_R g5811 ( 
.A(n_5626),
.Y(n_5811)
);

AOI22xp33_ASAP7_75t_L g5812 ( 
.A1(n_5734),
.A2(n_1355),
.B1(n_1988),
.B2(n_1984),
.Y(n_5812)
);

AOI22xp33_ASAP7_75t_SL g5813 ( 
.A1(n_5761),
.A2(n_224),
.B1(n_220),
.B2(n_222),
.Y(n_5813)
);

INVx4_ASAP7_75t_L g5814 ( 
.A(n_5614),
.Y(n_5814)
);

INVx6_ASAP7_75t_L g5815 ( 
.A(n_5607),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5632),
.Y(n_5816)
);

AND2x2_ASAP7_75t_L g5817 ( 
.A(n_5619),
.B(n_225),
.Y(n_5817)
);

AOI22xp33_ASAP7_75t_L g5818 ( 
.A1(n_5617),
.A2(n_1355),
.B1(n_1997),
.B2(n_1988),
.Y(n_5818)
);

AOI22xp33_ASAP7_75t_SL g5819 ( 
.A1(n_5678),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_L g5820 ( 
.A(n_5610),
.B(n_228),
.Y(n_5820)
);

INVx2_ASAP7_75t_L g5821 ( 
.A(n_5756),
.Y(n_5821)
);

INVx4_ASAP7_75t_SL g5822 ( 
.A(n_5616),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_5639),
.Y(n_5823)
);

OAI22xp5_ASAP7_75t_L g5824 ( 
.A1(n_5717),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_5824)
);

BUFx4f_ASAP7_75t_SL g5825 ( 
.A(n_5633),
.Y(n_5825)
);

CKINVDCx11_ASAP7_75t_R g5826 ( 
.A(n_5588),
.Y(n_5826)
);

OAI22xp5_ASAP7_75t_L g5827 ( 
.A1(n_5590),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_5827)
);

BUFx3_ASAP7_75t_L g5828 ( 
.A(n_5726),
.Y(n_5828)
);

OAI21xp33_ASAP7_75t_L g5829 ( 
.A1(n_5718),
.A2(n_233),
.B(n_234),
.Y(n_5829)
);

AOI222xp33_ASAP7_75t_L g5830 ( 
.A1(n_5696),
.A2(n_238),
.B1(n_240),
.B2(n_235),
.C1(n_237),
.C2(n_239),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_5640),
.Y(n_5831)
);

BUFx6f_ASAP7_75t_L g5832 ( 
.A(n_5699),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5686),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5643),
.Y(n_5834)
);

INVx2_ASAP7_75t_L g5835 ( 
.A(n_5686),
.Y(n_5835)
);

OAI22xp5_ASAP7_75t_L g5836 ( 
.A1(n_5634),
.A2(n_5612),
.B1(n_5624),
.B2(n_5635),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5652),
.Y(n_5837)
);

OAI21xp5_ASAP7_75t_SL g5838 ( 
.A1(n_5700),
.A2(n_241),
.B(n_243),
.Y(n_5838)
);

INVx2_ASAP7_75t_L g5839 ( 
.A(n_5629),
.Y(n_5839)
);

BUFx2_ASAP7_75t_L g5840 ( 
.A(n_5755),
.Y(n_5840)
);

AOI22xp33_ASAP7_75t_SL g5841 ( 
.A1(n_5661),
.A2(n_244),
.B1(n_241),
.B2(n_243),
.Y(n_5841)
);

AOI22xp33_ASAP7_75t_L g5842 ( 
.A1(n_5621),
.A2(n_1355),
.B1(n_1998),
.B2(n_1997),
.Y(n_5842)
);

AND2x4_ASAP7_75t_L g5843 ( 
.A(n_5630),
.B(n_246),
.Y(n_5843)
);

AOI22xp33_ASAP7_75t_L g5844 ( 
.A1(n_5642),
.A2(n_2004),
.B1(n_1998),
.B2(n_2504),
.Y(n_5844)
);

NAND2xp5_ASAP7_75t_L g5845 ( 
.A(n_5740),
.B(n_246),
.Y(n_5845)
);

NAND2xp5_ASAP7_75t_L g5846 ( 
.A(n_5740),
.B(n_247),
.Y(n_5846)
);

AND2x2_ASAP7_75t_L g5847 ( 
.A(n_5677),
.B(n_248),
.Y(n_5847)
);

AOI22xp33_ASAP7_75t_SL g5848 ( 
.A1(n_5671),
.A2(n_251),
.B1(n_248),
.B2(n_250),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5667),
.Y(n_5849)
);

AOI22xp33_ASAP7_75t_L g5850 ( 
.A1(n_5599),
.A2(n_2004),
.B1(n_2513),
.B2(n_2504),
.Y(n_5850)
);

INVx5_ASAP7_75t_SL g5851 ( 
.A(n_5723),
.Y(n_5851)
);

AOI22xp33_ASAP7_75t_L g5852 ( 
.A1(n_5602),
.A2(n_2513),
.B1(n_2521),
.B2(n_2504),
.Y(n_5852)
);

OAI22xp5_ASAP7_75t_L g5853 ( 
.A1(n_5682),
.A2(n_253),
.B1(n_250),
.B2(n_252),
.Y(n_5853)
);

BUFx4f_ASAP7_75t_SL g5854 ( 
.A(n_5732),
.Y(n_5854)
);

OAI22xp5_ASAP7_75t_L g5855 ( 
.A1(n_5635),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_5855)
);

AOI22xp33_ASAP7_75t_L g5856 ( 
.A1(n_5651),
.A2(n_2513),
.B1(n_2521),
.B2(n_2504),
.Y(n_5856)
);

CKINVDCx20_ASAP7_75t_R g5857 ( 
.A(n_5613),
.Y(n_5857)
);

AOI22xp33_ASAP7_75t_SL g5858 ( 
.A1(n_5690),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_5858)
);

AOI22xp33_ASAP7_75t_SL g5859 ( 
.A1(n_5666),
.A2(n_260),
.B1(n_257),
.B2(n_259),
.Y(n_5859)
);

AOI22xp33_ASAP7_75t_SL g5860 ( 
.A1(n_5677),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_5860)
);

INVx1_ASAP7_75t_SL g5861 ( 
.A(n_5753),
.Y(n_5861)
);

CKINVDCx5p33_ASAP7_75t_R g5862 ( 
.A(n_5712),
.Y(n_5862)
);

BUFx12f_ASAP7_75t_L g5863 ( 
.A(n_5725),
.Y(n_5863)
);

INVx3_ASAP7_75t_L g5864 ( 
.A(n_5614),
.Y(n_5864)
);

BUFx2_ASAP7_75t_L g5865 ( 
.A(n_5616),
.Y(n_5865)
);

CKINVDCx5p33_ASAP7_75t_R g5866 ( 
.A(n_5622),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5673),
.Y(n_5867)
);

AOI222xp33_ASAP7_75t_L g5868 ( 
.A1(n_5660),
.A2(n_264),
.B1(n_267),
.B2(n_261),
.C1(n_263),
.C2(n_266),
.Y(n_5868)
);

AOI22xp33_ASAP7_75t_L g5869 ( 
.A1(n_5644),
.A2(n_2521),
.B1(n_2568),
.B2(n_2513),
.Y(n_5869)
);

NAND2xp5_ASAP7_75t_L g5870 ( 
.A(n_5711),
.B(n_266),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5674),
.Y(n_5871)
);

NAND2xp5_ASAP7_75t_L g5872 ( 
.A(n_5720),
.B(n_270),
.Y(n_5872)
);

AOI22xp33_ASAP7_75t_SL g5873 ( 
.A1(n_5681),
.A2(n_275),
.B1(n_270),
.B2(n_272),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5676),
.Y(n_5874)
);

OAI22xp5_ASAP7_75t_SL g5875 ( 
.A1(n_5653),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5680),
.Y(n_5876)
);

AOI22xp5_ASAP7_75t_L g5877 ( 
.A1(n_5681),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_5877)
);

BUFx2_ASAP7_75t_L g5878 ( 
.A(n_5616),
.Y(n_5878)
);

AND2x2_ASAP7_75t_L g5879 ( 
.A(n_5730),
.B(n_280),
.Y(n_5879)
);

OAI222xp33_ASAP7_75t_L g5880 ( 
.A1(n_5648),
.A2(n_283),
.B1(n_288),
.B2(n_280),
.C1(n_282),
.C2(n_286),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_5685),
.Y(n_5881)
);

AOI22xp33_ASAP7_75t_L g5882 ( 
.A1(n_5703),
.A2(n_2568),
.B1(n_2580),
.B2(n_2521),
.Y(n_5882)
);

AOI22xp33_ASAP7_75t_L g5883 ( 
.A1(n_5589),
.A2(n_2580),
.B1(n_2568),
.B2(n_1916),
.Y(n_5883)
);

AOI22xp33_ASAP7_75t_L g5884 ( 
.A1(n_5645),
.A2(n_2580),
.B1(n_2568),
.B2(n_1916),
.Y(n_5884)
);

NOR2xp33_ASAP7_75t_L g5885 ( 
.A(n_5706),
.B(n_5708),
.Y(n_5885)
);

AOI22xp33_ASAP7_75t_SL g5886 ( 
.A1(n_5649),
.A2(n_288),
.B1(n_283),
.B2(n_286),
.Y(n_5886)
);

AOI22xp33_ASAP7_75t_L g5887 ( 
.A1(n_5741),
.A2(n_1916),
.B1(n_1928),
.B2(n_1926),
.Y(n_5887)
);

NOR2xp33_ASAP7_75t_L g5888 ( 
.A(n_5722),
.B(n_292),
.Y(n_5888)
);

AOI22xp33_ASAP7_75t_L g5889 ( 
.A1(n_5749),
.A2(n_1916),
.B1(n_1928),
.B2(n_1926),
.Y(n_5889)
);

OAI21xp5_ASAP7_75t_SL g5890 ( 
.A1(n_5733),
.A2(n_295),
.B(n_296),
.Y(n_5890)
);

BUFx4f_ASAP7_75t_SL g5891 ( 
.A(n_5669),
.Y(n_5891)
);

CKINVDCx5p33_ASAP7_75t_R g5892 ( 
.A(n_5716),
.Y(n_5892)
);

BUFx4f_ASAP7_75t_SL g5893 ( 
.A(n_5704),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5688),
.Y(n_5894)
);

OAI22xp5_ASAP7_75t_L g5895 ( 
.A1(n_5754),
.A2(n_300),
.B1(n_297),
.B2(n_298),
.Y(n_5895)
);

AOI22xp33_ASAP7_75t_L g5896 ( 
.A1(n_5592),
.A2(n_1928),
.B1(n_1938),
.B2(n_1926),
.Y(n_5896)
);

AOI22xp33_ASAP7_75t_L g5897 ( 
.A1(n_5592),
.A2(n_1928),
.B1(n_1938),
.B2(n_1926),
.Y(n_5897)
);

AOI222xp33_ASAP7_75t_L g5898 ( 
.A1(n_5744),
.A2(n_307),
.B1(n_309),
.B2(n_301),
.C1(n_306),
.C2(n_308),
.Y(n_5898)
);

AOI22xp33_ASAP7_75t_L g5899 ( 
.A1(n_5704),
.A2(n_1938),
.B1(n_1941),
.B2(n_1926),
.Y(n_5899)
);

OAI21xp5_ASAP7_75t_SL g5900 ( 
.A1(n_5586),
.A2(n_307),
.B(n_308),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_5693),
.B(n_310),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5688),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5688),
.Y(n_5903)
);

AOI22xp33_ASAP7_75t_L g5904 ( 
.A1(n_5601),
.A2(n_1941),
.B1(n_1942),
.B2(n_1938),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5630),
.B(n_310),
.Y(n_5905)
);

BUFx2_ASAP7_75t_L g5906 ( 
.A(n_5615),
.Y(n_5906)
);

HB1xp67_ASAP7_75t_L g5907 ( 
.A(n_5597),
.Y(n_5907)
);

OAI22xp5_ASAP7_75t_L g5908 ( 
.A1(n_5738),
.A2(n_315),
.B1(n_311),
.B2(n_314),
.Y(n_5908)
);

AND2x2_ASAP7_75t_L g5909 ( 
.A(n_5707),
.B(n_314),
.Y(n_5909)
);

HB1xp67_ASAP7_75t_L g5910 ( 
.A(n_5641),
.Y(n_5910)
);

AOI22xp33_ASAP7_75t_SL g5911 ( 
.A1(n_5684),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_5911)
);

CKINVDCx6p67_ASAP7_75t_R g5912 ( 
.A(n_5727),
.Y(n_5912)
);

OAI22xp33_ASAP7_75t_L g5913 ( 
.A1(n_5647),
.A2(n_321),
.B1(n_317),
.B2(n_319),
.Y(n_5913)
);

HB1xp67_ASAP7_75t_L g5914 ( 
.A(n_5641),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5724),
.Y(n_5915)
);

INVx2_ASAP7_75t_SL g5916 ( 
.A(n_5719),
.Y(n_5916)
);

AOI22xp33_ASAP7_75t_L g5917 ( 
.A1(n_5615),
.A2(n_5587),
.B1(n_5638),
.B2(n_5603),
.Y(n_5917)
);

AOI22xp33_ASAP7_75t_L g5918 ( 
.A1(n_5615),
.A2(n_1941),
.B1(n_1942),
.B2(n_1938),
.Y(n_5918)
);

AND2x2_ASAP7_75t_L g5919 ( 
.A(n_5698),
.B(n_325),
.Y(n_5919)
);

NAND2xp5_ASAP7_75t_L g5920 ( 
.A(n_5742),
.B(n_326),
.Y(n_5920)
);

CKINVDCx5p33_ASAP7_75t_R g5921 ( 
.A(n_5719),
.Y(n_5921)
);

AOI22xp33_ASAP7_75t_L g5922 ( 
.A1(n_5715),
.A2(n_1942),
.B1(n_1941),
.B2(n_1920),
.Y(n_5922)
);

AOI22xp33_ASAP7_75t_SL g5923 ( 
.A1(n_5654),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_5923)
);

AOI22xp33_ASAP7_75t_L g5924 ( 
.A1(n_5709),
.A2(n_1942),
.B1(n_1920),
.B2(n_1908),
.Y(n_5924)
);

HB1xp67_ASAP7_75t_L g5925 ( 
.A(n_5910),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5783),
.Y(n_5926)
);

AO21x2_ASAP7_75t_L g5927 ( 
.A1(n_5914),
.A2(n_5692),
.B(n_5710),
.Y(n_5927)
);

INVx3_ASAP7_75t_L g5928 ( 
.A(n_5832),
.Y(n_5928)
);

OR2x2_ASAP7_75t_L g5929 ( 
.A(n_5762),
.B(n_5737),
.Y(n_5929)
);

AND2x2_ASAP7_75t_L g5930 ( 
.A(n_5840),
.B(n_5664),
.Y(n_5930)
);

BUFx2_ASAP7_75t_L g5931 ( 
.A(n_5832),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_5894),
.B(n_5694),
.Y(n_5932)
);

AND2x2_ASAP7_75t_L g5933 ( 
.A(n_5809),
.B(n_5670),
.Y(n_5933)
);

INVx2_ASAP7_75t_SL g5934 ( 
.A(n_5765),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5763),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5767),
.Y(n_5936)
);

NAND2xp5_ASAP7_75t_L g5937 ( 
.A(n_5902),
.B(n_5657),
.Y(n_5937)
);

BUFx3_ASAP7_75t_L g5938 ( 
.A(n_5832),
.Y(n_5938)
);

NAND2xp5_ASAP7_75t_L g5939 ( 
.A(n_5903),
.B(n_5657),
.Y(n_5939)
);

AND2x2_ASAP7_75t_L g5940 ( 
.A(n_5821),
.B(n_5728),
.Y(n_5940)
);

AND2x4_ASAP7_75t_L g5941 ( 
.A(n_5822),
.B(n_5662),
.Y(n_5941)
);

AND2x2_ASAP7_75t_L g5942 ( 
.A(n_5778),
.B(n_5628),
.Y(n_5942)
);

AND2x2_ASAP7_75t_L g5943 ( 
.A(n_5789),
.B(n_5691),
.Y(n_5943)
);

AND2x2_ASAP7_75t_L g5944 ( 
.A(n_5912),
.B(n_5691),
.Y(n_5944)
);

AOI22xp33_ASAP7_75t_L g5945 ( 
.A1(n_5801),
.A2(n_5751),
.B1(n_5758),
.B2(n_5731),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5916),
.B(n_5636),
.Y(n_5946)
);

OAI22xp5_ASAP7_75t_L g5947 ( 
.A1(n_5886),
.A2(n_5697),
.B1(n_5689),
.B2(n_5746),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5839),
.B(n_5600),
.Y(n_5948)
);

HB1xp67_ASAP7_75t_L g5949 ( 
.A(n_5795),
.Y(n_5949)
);

NAND2xp5_ASAP7_75t_L g5950 ( 
.A(n_5915),
.B(n_5655),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5810),
.Y(n_5951)
);

INVx2_ASAP7_75t_L g5952 ( 
.A(n_5843),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5816),
.Y(n_5953)
);

OAI22xp5_ASAP7_75t_L g5954 ( 
.A1(n_5770),
.A2(n_5759),
.B1(n_5735),
.B2(n_5745),
.Y(n_5954)
);

INVx1_ASAP7_75t_L g5955 ( 
.A(n_5823),
.Y(n_5955)
);

AND2x2_ASAP7_75t_L g5956 ( 
.A(n_5864),
.B(n_5702),
.Y(n_5956)
);

INVx2_ASAP7_75t_L g5957 ( 
.A(n_5828),
.Y(n_5957)
);

BUFx3_ASAP7_75t_L g5958 ( 
.A(n_5815),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5843),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5831),
.Y(n_5960)
);

AND2x2_ASAP7_75t_L g5961 ( 
.A(n_5864),
.B(n_5736),
.Y(n_5961)
);

AND2x2_ASAP7_75t_L g5962 ( 
.A(n_5766),
.B(n_5743),
.Y(n_5962)
);

INVx2_ASAP7_75t_SL g5963 ( 
.A(n_5815),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5834),
.Y(n_5964)
);

AND2x4_ASAP7_75t_L g5965 ( 
.A(n_5822),
.B(n_5757),
.Y(n_5965)
);

INVxp67_ASAP7_75t_SL g5966 ( 
.A(n_5907),
.Y(n_5966)
);

BUFx3_ASAP7_75t_L g5967 ( 
.A(n_5863),
.Y(n_5967)
);

AND2x2_ASAP7_75t_L g5968 ( 
.A(n_5906),
.B(n_331),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5837),
.Y(n_5969)
);

AOI22xp33_ASAP7_75t_L g5970 ( 
.A1(n_5790),
.A2(n_336),
.B1(n_332),
.B2(n_335),
.Y(n_5970)
);

AND2x2_ASAP7_75t_L g5971 ( 
.A(n_5885),
.B(n_332),
.Y(n_5971)
);

AO31x2_ASAP7_75t_L g5972 ( 
.A1(n_5865),
.A2(n_338),
.A3(n_336),
.B(n_337),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5849),
.Y(n_5973)
);

AND2x2_ASAP7_75t_L g5974 ( 
.A(n_5878),
.B(n_337),
.Y(n_5974)
);

INVx2_ASAP7_75t_L g5975 ( 
.A(n_5814),
.Y(n_5975)
);

INVx2_ASAP7_75t_SL g5976 ( 
.A(n_5825),
.Y(n_5976)
);

AOI22xp33_ASAP7_75t_L g5977 ( 
.A1(n_5829),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_5977)
);

HB1xp67_ASAP7_75t_L g5978 ( 
.A(n_5919),
.Y(n_5978)
);

NAND2xp5_ASAP7_75t_L g5979 ( 
.A(n_5867),
.B(n_342),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5871),
.Y(n_5980)
);

AND2x4_ASAP7_75t_L g5981 ( 
.A(n_5833),
.B(n_342),
.Y(n_5981)
);

AND2x2_ASAP7_75t_L g5982 ( 
.A(n_5811),
.B(n_343),
.Y(n_5982)
);

AOI22xp33_ASAP7_75t_L g5983 ( 
.A1(n_5780),
.A2(n_346),
.B1(n_343),
.B2(n_345),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5874),
.Y(n_5984)
);

BUFx3_ASAP7_75t_L g5985 ( 
.A(n_5854),
.Y(n_5985)
);

OR2x2_ASAP7_75t_L g5986 ( 
.A(n_5835),
.B(n_5917),
.Y(n_5986)
);

INVx2_ASAP7_75t_L g5987 ( 
.A(n_5921),
.Y(n_5987)
);

NAND2xp5_ASAP7_75t_L g5988 ( 
.A(n_5876),
.B(n_5881),
.Y(n_5988)
);

BUFx2_ASAP7_75t_L g5989 ( 
.A(n_5893),
.Y(n_5989)
);

BUFx2_ASAP7_75t_L g5990 ( 
.A(n_5796),
.Y(n_5990)
);

BUFx3_ASAP7_75t_L g5991 ( 
.A(n_5826),
.Y(n_5991)
);

AND2x2_ASAP7_75t_L g5992 ( 
.A(n_5776),
.B(n_348),
.Y(n_5992)
);

INVxp33_ASAP7_75t_L g5993 ( 
.A(n_5836),
.Y(n_5993)
);

INVx2_ASAP7_75t_L g5994 ( 
.A(n_5891),
.Y(n_5994)
);

BUFx3_ASAP7_75t_L g5995 ( 
.A(n_5857),
.Y(n_5995)
);

INVx2_ASAP7_75t_L g5996 ( 
.A(n_5905),
.Y(n_5996)
);

AND2x2_ASAP7_75t_L g5997 ( 
.A(n_5776),
.B(n_349),
.Y(n_5997)
);

HB1xp67_ASAP7_75t_L g5998 ( 
.A(n_5851),
.Y(n_5998)
);

HB1xp67_ASAP7_75t_L g5999 ( 
.A(n_5851),
.Y(n_5999)
);

HB1xp67_ASAP7_75t_L g6000 ( 
.A(n_5851),
.Y(n_6000)
);

BUFx3_ASAP7_75t_L g6001 ( 
.A(n_5782),
.Y(n_6001)
);

INVx1_ASAP7_75t_L g6002 ( 
.A(n_5909),
.Y(n_6002)
);

AND2x2_ASAP7_75t_L g6003 ( 
.A(n_5776),
.B(n_350),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_L g6004 ( 
.A(n_5856),
.B(n_351),
.Y(n_6004)
);

INVx1_ASAP7_75t_L g6005 ( 
.A(n_5870),
.Y(n_6005)
);

INVx2_ASAP7_75t_L g6006 ( 
.A(n_5792),
.Y(n_6006)
);

NAND2xp5_ASAP7_75t_L g6007 ( 
.A(n_5923),
.B(n_351),
.Y(n_6007)
);

AND2x2_ASAP7_75t_L g6008 ( 
.A(n_5792),
.B(n_352),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5872),
.Y(n_6009)
);

OAI22xp5_ASAP7_75t_L g6010 ( 
.A1(n_5861),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_6010)
);

INVx2_ASAP7_75t_L g6011 ( 
.A(n_5792),
.Y(n_6011)
);

BUFx6f_ASAP7_75t_L g6012 ( 
.A(n_5847),
.Y(n_6012)
);

AND2x2_ASAP7_75t_L g6013 ( 
.A(n_5799),
.B(n_355),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5901),
.Y(n_6014)
);

AND2x2_ASAP7_75t_L g6015 ( 
.A(n_5817),
.B(n_356),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5820),
.Y(n_6016)
);

AOI22xp33_ASAP7_75t_L g6017 ( 
.A1(n_5827),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5879),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5794),
.Y(n_6019)
);

INVx2_ASAP7_75t_L g6020 ( 
.A(n_5794),
.Y(n_6020)
);

INVx2_ASAP7_75t_L g6021 ( 
.A(n_5892),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5793),
.Y(n_6022)
);

NOR2xp33_ASAP7_75t_L g6023 ( 
.A(n_5861),
.B(n_363),
.Y(n_6023)
);

AOI22xp33_ASAP7_75t_SL g6024 ( 
.A1(n_5784),
.A2(n_367),
.B1(n_364),
.B2(n_365),
.Y(n_6024)
);

AND2x2_ASAP7_75t_L g6025 ( 
.A(n_5883),
.B(n_364),
.Y(n_6025)
);

INVx2_ASAP7_75t_L g6026 ( 
.A(n_5777),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5862),
.B(n_365),
.Y(n_6027)
);

INVx2_ASAP7_75t_L g6028 ( 
.A(n_5845),
.Y(n_6028)
);

NAND2xp5_ASAP7_75t_L g6029 ( 
.A(n_5785),
.B(n_369),
.Y(n_6029)
);

INVx3_ASAP7_75t_L g6030 ( 
.A(n_5866),
.Y(n_6030)
);

BUFx3_ASAP7_75t_L g6031 ( 
.A(n_5772),
.Y(n_6031)
);

INVx3_ASAP7_75t_L g6032 ( 
.A(n_5846),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5920),
.Y(n_6033)
);

BUFx3_ASAP7_75t_L g6034 ( 
.A(n_5791),
.Y(n_6034)
);

AND2x4_ASAP7_75t_L g6035 ( 
.A(n_5775),
.B(n_370),
.Y(n_6035)
);

INVx1_ASAP7_75t_SL g6036 ( 
.A(n_5875),
.Y(n_6036)
);

AOI22xp33_ASAP7_75t_L g6037 ( 
.A1(n_5827),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_6037)
);

HB1xp67_ASAP7_75t_L g6038 ( 
.A(n_5880),
.Y(n_6038)
);

BUFx6f_ASAP7_75t_L g6039 ( 
.A(n_5888),
.Y(n_6039)
);

AND2x4_ASAP7_75t_L g6040 ( 
.A(n_5775),
.B(n_372),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5855),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5904),
.B(n_374),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_5853),
.Y(n_6043)
);

AOI22xp33_ASAP7_75t_L g6044 ( 
.A1(n_5813),
.A2(n_379),
.B1(n_375),
.B2(n_377),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5781),
.B(n_375),
.Y(n_6045)
);

AND2x2_ASAP7_75t_L g6046 ( 
.A(n_5764),
.B(n_377),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5853),
.Y(n_6047)
);

BUFx2_ASAP7_75t_L g6048 ( 
.A(n_5800),
.Y(n_6048)
);

AND2x2_ASAP7_75t_L g6049 ( 
.A(n_5869),
.B(n_379),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5925),
.Y(n_6050)
);

INVx3_ASAP7_75t_L g6051 ( 
.A(n_5985),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5925),
.Y(n_6052)
);

INVx2_ASAP7_75t_L g6053 ( 
.A(n_5985),
.Y(n_6053)
);

AND2x4_ASAP7_75t_L g6054 ( 
.A(n_5991),
.B(n_5800),
.Y(n_6054)
);

NOR2x2_ASAP7_75t_L g6055 ( 
.A(n_6006),
.B(n_5900),
.Y(n_6055)
);

AND2x2_ASAP7_75t_L g6056 ( 
.A(n_5931),
.B(n_5976),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5949),
.Y(n_6057)
);

NAND2xp5_ASAP7_75t_L g6058 ( 
.A(n_6038),
.B(n_5805),
.Y(n_6058)
);

AND2x2_ASAP7_75t_L g6059 ( 
.A(n_5989),
.B(n_5852),
.Y(n_6059)
);

NAND2xp5_ASAP7_75t_L g6060 ( 
.A(n_6038),
.B(n_5807),
.Y(n_6060)
);

AND2x2_ASAP7_75t_L g6061 ( 
.A(n_5928),
.B(n_5768),
.Y(n_6061)
);

BUFx2_ASAP7_75t_L g6062 ( 
.A(n_5938),
.Y(n_6062)
);

CKINVDCx5p33_ASAP7_75t_R g6063 ( 
.A(n_5938),
.Y(n_6063)
);

HB1xp67_ASAP7_75t_L g6064 ( 
.A(n_5978),
.Y(n_6064)
);

AND2x2_ASAP7_75t_L g6065 ( 
.A(n_5928),
.B(n_5890),
.Y(n_6065)
);

NAND2xp5_ASAP7_75t_L g6066 ( 
.A(n_6048),
.B(n_5788),
.Y(n_6066)
);

BUFx4f_ASAP7_75t_L g6067 ( 
.A(n_5992),
.Y(n_6067)
);

OAI22xp5_ASAP7_75t_L g6068 ( 
.A1(n_5977),
.A2(n_5786),
.B1(n_5911),
.B2(n_5890),
.Y(n_6068)
);

INVx2_ASAP7_75t_L g6069 ( 
.A(n_5958),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_5966),
.Y(n_6070)
);

AOI22xp33_ASAP7_75t_L g6071 ( 
.A1(n_5990),
.A2(n_5779),
.B1(n_5787),
.B2(n_5830),
.Y(n_6071)
);

AND2x2_ASAP7_75t_L g6072 ( 
.A(n_6011),
.B(n_5771),
.Y(n_6072)
);

NAND2xp5_ASAP7_75t_L g6073 ( 
.A(n_6046),
.B(n_5786),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5926),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_5988),
.Y(n_6075)
);

AND2x2_ASAP7_75t_L g6076 ( 
.A(n_5930),
.B(n_5963),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_5994),
.B(n_5771),
.Y(n_6077)
);

AND2x2_ASAP7_75t_L g6078 ( 
.A(n_5996),
.B(n_5769),
.Y(n_6078)
);

AND2x2_ASAP7_75t_L g6079 ( 
.A(n_5996),
.B(n_5850),
.Y(n_6079)
);

BUFx2_ASAP7_75t_SL g6080 ( 
.A(n_5995),
.Y(n_6080)
);

BUFx2_ASAP7_75t_L g6081 ( 
.A(n_5952),
.Y(n_6081)
);

HB1xp67_ASAP7_75t_L g6082 ( 
.A(n_5927),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5988),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_6002),
.Y(n_6084)
);

INVx2_ASAP7_75t_L g6085 ( 
.A(n_6001),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5935),
.Y(n_6086)
);

AND2x4_ASAP7_75t_L g6087 ( 
.A(n_5934),
.B(n_5877),
.Y(n_6087)
);

BUFx2_ASAP7_75t_L g6088 ( 
.A(n_5952),
.Y(n_6088)
);

BUFx3_ASAP7_75t_L g6089 ( 
.A(n_5995),
.Y(n_6089)
);

NAND2xp5_ASAP7_75t_L g6090 ( 
.A(n_6036),
.B(n_5838),
.Y(n_6090)
);

NAND2xp5_ASAP7_75t_L g6091 ( 
.A(n_6036),
.B(n_5830),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_5936),
.Y(n_6092)
);

AND2x2_ASAP7_75t_L g6093 ( 
.A(n_5957),
.B(n_5774),
.Y(n_6093)
);

AND2x2_ASAP7_75t_L g6094 ( 
.A(n_5959),
.B(n_5798),
.Y(n_6094)
);

AND2x2_ASAP7_75t_L g6095 ( 
.A(n_5940),
.B(n_5884),
.Y(n_6095)
);

NAND2xp5_ASAP7_75t_L g6096 ( 
.A(n_6043),
.B(n_5913),
.Y(n_6096)
);

HB1xp67_ASAP7_75t_L g6097 ( 
.A(n_5927),
.Y(n_6097)
);

BUFx6f_ASAP7_75t_SL g6098 ( 
.A(n_5967),
.Y(n_6098)
);

BUFx2_ASAP7_75t_L g6099 ( 
.A(n_6031),
.Y(n_6099)
);

BUFx2_ASAP7_75t_L g6100 ( 
.A(n_6031),
.Y(n_6100)
);

INVx2_ASAP7_75t_L g6101 ( 
.A(n_6012),
.Y(n_6101)
);

HB1xp67_ASAP7_75t_L g6102 ( 
.A(n_5998),
.Y(n_6102)
);

NOR2x1_ASAP7_75t_SL g6103 ( 
.A(n_6012),
.B(n_5908),
.Y(n_6103)
);

BUFx2_ASAP7_75t_L g6104 ( 
.A(n_6012),
.Y(n_6104)
);

INVx2_ASAP7_75t_SL g6105 ( 
.A(n_6012),
.Y(n_6105)
);

AND2x2_ASAP7_75t_L g6106 ( 
.A(n_6030),
.B(n_5882),
.Y(n_6106)
);

BUFx3_ASAP7_75t_L g6107 ( 
.A(n_5997),
.Y(n_6107)
);

AND2x2_ASAP7_75t_L g6108 ( 
.A(n_6030),
.B(n_5933),
.Y(n_6108)
);

HB1xp67_ASAP7_75t_L g6109 ( 
.A(n_5998),
.Y(n_6109)
);

BUFx6f_ASAP7_75t_L g6110 ( 
.A(n_6003),
.Y(n_6110)
);

NAND2xp5_ASAP7_75t_L g6111 ( 
.A(n_6047),
.B(n_5868),
.Y(n_6111)
);

INVx2_ASAP7_75t_SL g6112 ( 
.A(n_6008),
.Y(n_6112)
);

BUFx3_ASAP7_75t_L g6113 ( 
.A(n_5982),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_5951),
.Y(n_6114)
);

OR2x2_ASAP7_75t_L g6115 ( 
.A(n_6018),
.B(n_5895),
.Y(n_6115)
);

BUFx3_ASAP7_75t_L g6116 ( 
.A(n_5981),
.Y(n_6116)
);

BUFx3_ASAP7_75t_L g6117 ( 
.A(n_5981),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5953),
.Y(n_6118)
);

AND2x2_ASAP7_75t_L g6119 ( 
.A(n_5987),
.B(n_6021),
.Y(n_6119)
);

AND2x2_ASAP7_75t_L g6120 ( 
.A(n_5944),
.B(n_5896),
.Y(n_6120)
);

INVxp67_ASAP7_75t_SL g6121 ( 
.A(n_6023),
.Y(n_6121)
);

BUFx6f_ASAP7_75t_L g6122 ( 
.A(n_6027),
.Y(n_6122)
);

AND2x4_ASAP7_75t_SL g6123 ( 
.A(n_5941),
.B(n_5773),
.Y(n_6123)
);

NAND2xp5_ASAP7_75t_L g6124 ( 
.A(n_6032),
.B(n_5868),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_6032),
.B(n_5819),
.Y(n_6125)
);

AND2x2_ASAP7_75t_L g6126 ( 
.A(n_5942),
.B(n_5897),
.Y(n_6126)
);

AOI22xp33_ASAP7_75t_L g6127 ( 
.A1(n_5993),
.A2(n_5824),
.B1(n_5858),
.B2(n_5859),
.Y(n_6127)
);

NOR2x1_ASAP7_75t_R g6128 ( 
.A(n_6034),
.B(n_5860),
.Y(n_6128)
);

INVx2_ASAP7_75t_L g6129 ( 
.A(n_5975),
.Y(n_6129)
);

INVx1_ASAP7_75t_SL g6130 ( 
.A(n_5968),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5955),
.Y(n_6131)
);

AND2x2_ASAP7_75t_L g6132 ( 
.A(n_6034),
.B(n_5873),
.Y(n_6132)
);

INVx2_ASAP7_75t_L g6133 ( 
.A(n_6022),
.Y(n_6133)
);

NAND2xp5_ASAP7_75t_L g6134 ( 
.A(n_6041),
.B(n_5804),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_5943),
.B(n_5844),
.Y(n_6135)
);

AND2x2_ASAP7_75t_L g6136 ( 
.A(n_6014),
.B(n_5802),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5960),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_5964),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_5969),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_5973),
.Y(n_6140)
);

INVx5_ASAP7_75t_L g6141 ( 
.A(n_6039),
.Y(n_6141)
);

AND2x2_ASAP7_75t_L g6142 ( 
.A(n_5946),
.B(n_5803),
.Y(n_6142)
);

NAND2xp5_ASAP7_75t_L g6143 ( 
.A(n_6033),
.B(n_5824),
.Y(n_6143)
);

HB1xp67_ASAP7_75t_L g6144 ( 
.A(n_5999),
.Y(n_6144)
);

INVx2_ASAP7_75t_L g6145 ( 
.A(n_6019),
.Y(n_6145)
);

OAI21xp33_ASAP7_75t_L g6146 ( 
.A1(n_5993),
.A2(n_5841),
.B(n_5848),
.Y(n_6146)
);

NAND2xp5_ASAP7_75t_L g6147 ( 
.A(n_6064),
.B(n_6023),
.Y(n_6147)
);

NAND2xp5_ASAP7_75t_L g6148 ( 
.A(n_6071),
.B(n_6026),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_6082),
.Y(n_6149)
);

OR2x2_ASAP7_75t_L g6150 ( 
.A(n_6130),
.B(n_5932),
.Y(n_6150)
);

INVx2_ASAP7_75t_SL g6151 ( 
.A(n_6141),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_6082),
.Y(n_6152)
);

NAND2xp5_ASAP7_75t_L g6153 ( 
.A(n_6071),
.B(n_6028),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_6097),
.Y(n_6154)
);

INVx1_ASAP7_75t_L g6155 ( 
.A(n_6097),
.Y(n_6155)
);

HB1xp67_ASAP7_75t_L g6156 ( 
.A(n_6102),
.Y(n_6156)
);

INVx2_ASAP7_75t_L g6157 ( 
.A(n_6141),
.Y(n_6157)
);

BUFx3_ASAP7_75t_L g6158 ( 
.A(n_6099),
.Y(n_6158)
);

NAND2xp5_ASAP7_75t_L g6159 ( 
.A(n_6121),
.B(n_5974),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_6102),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_6141),
.Y(n_6161)
);

BUFx2_ASAP7_75t_L g6162 ( 
.A(n_6100),
.Y(n_6162)
);

INVxp67_ASAP7_75t_L g6163 ( 
.A(n_6080),
.Y(n_6163)
);

INVxp67_ASAP7_75t_SL g6164 ( 
.A(n_6128),
.Y(n_6164)
);

AND2x4_ASAP7_75t_L g6165 ( 
.A(n_6141),
.B(n_6000),
.Y(n_6165)
);

INVx2_ASAP7_75t_SL g6166 ( 
.A(n_6062),
.Y(n_6166)
);

AND2x2_ASAP7_75t_L g6167 ( 
.A(n_6056),
.B(n_6076),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_6109),
.Y(n_6168)
);

HB1xp67_ASAP7_75t_L g6169 ( 
.A(n_6144),
.Y(n_6169)
);

BUFx2_ASAP7_75t_L g6170 ( 
.A(n_6113),
.Y(n_6170)
);

NAND2xp5_ASAP7_75t_L g6171 ( 
.A(n_6127),
.B(n_6058),
.Y(n_6171)
);

INVxp67_ASAP7_75t_L g6172 ( 
.A(n_6104),
.Y(n_6172)
);

NAND2xp5_ASAP7_75t_L g6173 ( 
.A(n_6127),
.B(n_6016),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_6081),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_6088),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_6050),
.Y(n_6176)
);

INVxp67_ASAP7_75t_L g6177 ( 
.A(n_6110),
.Y(n_6177)
);

AOI21xp5_ASAP7_75t_L g6178 ( 
.A1(n_6060),
.A2(n_6000),
.B(n_6039),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_6089),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_6052),
.Y(n_6180)
);

AND2x2_ASAP7_75t_L g6181 ( 
.A(n_6051),
.B(n_6005),
.Y(n_6181)
);

AND2x4_ASAP7_75t_L g6182 ( 
.A(n_6116),
.B(n_5929),
.Y(n_6182)
);

AOI22xp33_ASAP7_75t_L g6183 ( 
.A1(n_6060),
.A2(n_6091),
.B1(n_6146),
.B2(n_6066),
.Y(n_6183)
);

INVx2_ASAP7_75t_SL g6184 ( 
.A(n_6063),
.Y(n_6184)
);

INVx8_ASAP7_75t_L g6185 ( 
.A(n_6098),
.Y(n_6185)
);

HB1xp67_ASAP7_75t_L g6186 ( 
.A(n_6070),
.Y(n_6186)
);

BUFx3_ASAP7_75t_L g6187 ( 
.A(n_6110),
.Y(n_6187)
);

AND2x2_ASAP7_75t_L g6188 ( 
.A(n_6065),
.B(n_6009),
.Y(n_6188)
);

OR2x2_ASAP7_75t_L g6189 ( 
.A(n_6090),
.B(n_5986),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_6057),
.Y(n_6190)
);

AND2x4_ASAP7_75t_L g6191 ( 
.A(n_6116),
.B(n_6039),
.Y(n_6191)
);

AND2x2_ASAP7_75t_L g6192 ( 
.A(n_6053),
.B(n_5971),
.Y(n_6192)
);

NAND2xp5_ASAP7_75t_L g6193 ( 
.A(n_6091),
.B(n_5980),
.Y(n_6193)
);

HB1xp67_ASAP7_75t_L g6194 ( 
.A(n_6117),
.Y(n_6194)
);

NAND2x1_ASAP7_75t_L g6195 ( 
.A(n_6110),
.B(n_5948),
.Y(n_6195)
);

AND2x2_ASAP7_75t_L g6196 ( 
.A(n_6069),
.B(n_5962),
.Y(n_6196)
);

BUFx3_ASAP7_75t_L g6197 ( 
.A(n_6063),
.Y(n_6197)
);

AND2x4_ASAP7_75t_L g6198 ( 
.A(n_6105),
.B(n_5984),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_6122),
.Y(n_6199)
);

INVx3_ASAP7_75t_L g6200 ( 
.A(n_6101),
.Y(n_6200)
);

INVx2_ASAP7_75t_L g6201 ( 
.A(n_6107),
.Y(n_6201)
);

NAND2x1_ASAP7_75t_L g6202 ( 
.A(n_6122),
.B(n_5965),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_6054),
.B(n_6020),
.Y(n_6203)
);

HB1xp67_ASAP7_75t_L g6204 ( 
.A(n_6112),
.Y(n_6204)
);

BUFx6f_ASAP7_75t_L g6205 ( 
.A(n_6122),
.Y(n_6205)
);

INVxp67_ASAP7_75t_SL g6206 ( 
.A(n_6103),
.Y(n_6206)
);

AND2x2_ASAP7_75t_L g6207 ( 
.A(n_6067),
.B(n_5945),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_6085),
.Y(n_6208)
);

HB1xp67_ASAP7_75t_L g6209 ( 
.A(n_6124),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_6133),
.Y(n_6210)
);

AND2x2_ASAP7_75t_L g6211 ( 
.A(n_6108),
.B(n_5945),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_6074),
.Y(n_6212)
);

NAND2xp5_ASAP7_75t_L g6213 ( 
.A(n_6068),
.B(n_6010),
.Y(n_6213)
);

OAI22xp33_ASAP7_75t_L g6214 ( 
.A1(n_6068),
.A2(n_6124),
.B1(n_5947),
.B2(n_6125),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_6084),
.Y(n_6215)
);

OR2x2_ASAP7_75t_L g6216 ( 
.A(n_6125),
.B(n_6073),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_6061),
.B(n_6015),
.Y(n_6217)
);

AND2x2_ASAP7_75t_L g6218 ( 
.A(n_6087),
.B(n_6119),
.Y(n_6218)
);

INVx1_ASAP7_75t_L g6219 ( 
.A(n_6086),
.Y(n_6219)
);

INVx1_ASAP7_75t_L g6220 ( 
.A(n_6092),
.Y(n_6220)
);

BUFx2_ASAP7_75t_L g6221 ( 
.A(n_6087),
.Y(n_6221)
);

AND2x2_ASAP7_75t_L g6222 ( 
.A(n_6132),
.B(n_6077),
.Y(n_6222)
);

AND2x2_ASAP7_75t_L g6223 ( 
.A(n_6072),
.B(n_6013),
.Y(n_6223)
);

INVx4_ASAP7_75t_L g6224 ( 
.A(n_6129),
.Y(n_6224)
);

INVx1_ASAP7_75t_L g6225 ( 
.A(n_6156),
.Y(n_6225)
);

CKINVDCx5p33_ASAP7_75t_R g6226 ( 
.A(n_6185),
.Y(n_6226)
);

AND2x2_ASAP7_75t_L g6227 ( 
.A(n_6221),
.B(n_6078),
.Y(n_6227)
);

NAND4xp25_ASAP7_75t_L g6228 ( 
.A(n_6183),
.B(n_6111),
.C(n_6096),
.D(n_6134),
.Y(n_6228)
);

AOI221xp5_ASAP7_75t_L g6229 ( 
.A1(n_6214),
.A2(n_6143),
.B1(n_6134),
.B2(n_6083),
.C(n_6075),
.Y(n_6229)
);

BUFx3_ASAP7_75t_L g6230 ( 
.A(n_6185),
.Y(n_6230)
);

AO21x2_ASAP7_75t_L g6231 ( 
.A1(n_6149),
.A2(n_6154),
.B(n_6152),
.Y(n_6231)
);

OR2x6_ASAP7_75t_L g6232 ( 
.A(n_6163),
.B(n_5979),
.Y(n_6232)
);

OAI221xp5_ASAP7_75t_L g6233 ( 
.A1(n_6183),
.A2(n_6024),
.B1(n_5977),
.B2(n_5970),
.C(n_5983),
.Y(n_6233)
);

AOI33xp33_ASAP7_75t_L g6234 ( 
.A1(n_6207),
.A2(n_6024),
.A3(n_6044),
.B1(n_6145),
.B2(n_5983),
.B3(n_5970),
.Y(n_6234)
);

AOI22xp33_ASAP7_75t_L g6235 ( 
.A1(n_6171),
.A2(n_6059),
.B1(n_6120),
.B2(n_6106),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_6169),
.Y(n_6236)
);

INVx2_ASAP7_75t_L g6237 ( 
.A(n_6205),
.Y(n_6237)
);

A2O1A1Ixp33_ASAP7_75t_L g6238 ( 
.A1(n_6206),
.A2(n_6035),
.B(n_6040),
.C(n_6007),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_6169),
.Y(n_6239)
);

OAI22xp33_ASAP7_75t_L g6240 ( 
.A1(n_6213),
.A2(n_5947),
.B1(n_6007),
.B2(n_6035),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_6194),
.Y(n_6241)
);

AOI22xp33_ASAP7_75t_L g6242 ( 
.A1(n_6164),
.A2(n_6095),
.B1(n_6126),
.B2(n_6135),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_6205),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_6194),
.Y(n_6244)
);

INVx2_ASAP7_75t_L g6245 ( 
.A(n_6205),
.Y(n_6245)
);

BUFx3_ASAP7_75t_L g6246 ( 
.A(n_6191),
.Y(n_6246)
);

AOI22xp33_ASAP7_75t_L g6247 ( 
.A1(n_6209),
.A2(n_6142),
.B1(n_6093),
.B2(n_6094),
.Y(n_6247)
);

OAI332xp33_ASAP7_75t_SL g6248 ( 
.A1(n_6209),
.A2(n_6055),
.A3(n_5954),
.B1(n_6115),
.B2(n_6137),
.B3(n_6114),
.C1(n_6131),
.C2(n_6139),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_6186),
.Y(n_6249)
);

INVx3_ASAP7_75t_L g6250 ( 
.A(n_6165),
.Y(n_6250)
);

NAND2xp33_ASAP7_75t_SL g6251 ( 
.A(n_6202),
.B(n_6079),
.Y(n_6251)
);

AOI221xp5_ASAP7_75t_L g6252 ( 
.A1(n_6178),
.A2(n_6140),
.B1(n_6138),
.B2(n_6118),
.C(n_5950),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_6186),
.Y(n_6253)
);

INVx1_ASAP7_75t_L g6254 ( 
.A(n_6204),
.Y(n_6254)
);

AND2x4_ASAP7_75t_L g6255 ( 
.A(n_6158),
.B(n_5979),
.Y(n_6255)
);

CKINVDCx20_ASAP7_75t_R g6256 ( 
.A(n_6197),
.Y(n_6256)
);

AND2x4_ASAP7_75t_L g6257 ( 
.A(n_6158),
.B(n_6136),
.Y(n_6257)
);

NAND5xp2_ASAP7_75t_SL g6258 ( 
.A(n_6167),
.B(n_6037),
.C(n_6017),
.D(n_5898),
.E(n_5961),
.Y(n_6258)
);

OAI211xp5_ASAP7_75t_SL g6259 ( 
.A1(n_6173),
.A2(n_6037),
.B(n_6017),
.C(n_5939),
.Y(n_6259)
);

NOR4xp25_ASAP7_75t_SL g6260 ( 
.A(n_6170),
.B(n_5972),
.C(n_5937),
.D(n_6123),
.Y(n_6260)
);

INVx1_ASAP7_75t_L g6261 ( 
.A(n_6204),
.Y(n_6261)
);

OAI211xp5_ASAP7_75t_L g6262 ( 
.A1(n_6178),
.A2(n_5898),
.B(n_6004),
.C(n_6029),
.Y(n_6262)
);

HB1xp67_ASAP7_75t_L g6263 ( 
.A(n_6162),
.Y(n_6263)
);

AND2x2_ASAP7_75t_L g6264 ( 
.A(n_6218),
.B(n_5956),
.Y(n_6264)
);

INVx2_ASAP7_75t_L g6265 ( 
.A(n_6187),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_6160),
.Y(n_6266)
);

OA21x2_ASAP7_75t_L g6267 ( 
.A1(n_6155),
.A2(n_6147),
.B(n_6148),
.Y(n_6267)
);

NAND4xp25_ASAP7_75t_SL g6268 ( 
.A(n_6148),
.B(n_6025),
.C(n_6042),
.D(n_6045),
.Y(n_6268)
);

AOI22xp33_ASAP7_75t_L g6269 ( 
.A1(n_6153),
.A2(n_5806),
.B1(n_5808),
.B2(n_6049),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_6168),
.Y(n_6270)
);

BUFx4f_ASAP7_75t_L g6271 ( 
.A(n_6184),
.Y(n_6271)
);

OAI22xp5_ASAP7_75t_L g6272 ( 
.A1(n_6189),
.A2(n_5797),
.B1(n_5922),
.B2(n_5899),
.Y(n_6272)
);

OAI221xp5_ASAP7_75t_L g6273 ( 
.A1(n_6216),
.A2(n_5889),
.B1(n_5887),
.B2(n_5812),
.C(n_5924),
.Y(n_6273)
);

INVx4_ASAP7_75t_L g6274 ( 
.A(n_6165),
.Y(n_6274)
);

OR2x6_ASAP7_75t_L g6275 ( 
.A(n_6166),
.B(n_5972),
.Y(n_6275)
);

OAI21x1_ASAP7_75t_L g6276 ( 
.A1(n_6195),
.A2(n_5918),
.B(n_5842),
.Y(n_6276)
);

INVx4_ASAP7_75t_L g6277 ( 
.A(n_6157),
.Y(n_6277)
);

INVx4_ASAP7_75t_L g6278 ( 
.A(n_6161),
.Y(n_6278)
);

OAI31xp33_ASAP7_75t_L g6279 ( 
.A1(n_6193),
.A2(n_5818),
.A3(n_381),
.B(n_380),
.Y(n_6279)
);

INVx3_ASAP7_75t_L g6280 ( 
.A(n_6182),
.Y(n_6280)
);

AOI22xp33_ASAP7_75t_L g6281 ( 
.A1(n_6211),
.A2(n_1340),
.B1(n_1236),
.B2(n_382),
.Y(n_6281)
);

AND2x4_ASAP7_75t_L g6282 ( 
.A(n_6151),
.B(n_384),
.Y(n_6282)
);

HB1xp67_ASAP7_75t_L g6283 ( 
.A(n_6177),
.Y(n_6283)
);

OR2x2_ASAP7_75t_L g6284 ( 
.A(n_6159),
.B(n_386),
.Y(n_6284)
);

INVx3_ASAP7_75t_L g6285 ( 
.A(n_6182),
.Y(n_6285)
);

OR2x6_ASAP7_75t_L g6286 ( 
.A(n_6179),
.B(n_387),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_6174),
.Y(n_6287)
);

AOI33xp33_ASAP7_75t_L g6288 ( 
.A1(n_6175),
.A2(n_389),
.A3(n_390),
.B1(n_391),
.B2(n_394),
.B3(n_395),
.Y(n_6288)
);

HB1xp67_ASAP7_75t_L g6289 ( 
.A(n_6201),
.Y(n_6289)
);

NAND3xp33_ASAP7_75t_L g6290 ( 
.A(n_6172),
.B(n_396),
.C(n_397),
.Y(n_6290)
);

NOR3xp33_ASAP7_75t_SL g6291 ( 
.A(n_6208),
.B(n_396),
.C(n_398),
.Y(n_6291)
);

HB1xp67_ASAP7_75t_L g6292 ( 
.A(n_6201),
.Y(n_6292)
);

AND2x2_ASAP7_75t_L g6293 ( 
.A(n_6227),
.B(n_6217),
.Y(n_6293)
);

HB1xp67_ASAP7_75t_L g6294 ( 
.A(n_6231),
.Y(n_6294)
);

NOR2xp33_ASAP7_75t_L g6295 ( 
.A(n_6274),
.B(n_6224),
.Y(n_6295)
);

INVx2_ASAP7_75t_L g6296 ( 
.A(n_6267),
.Y(n_6296)
);

NAND2xp5_ASAP7_75t_L g6297 ( 
.A(n_6267),
.B(n_6200),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_6230),
.B(n_6203),
.Y(n_6298)
);

INVx2_ASAP7_75t_L g6299 ( 
.A(n_6250),
.Y(n_6299)
);

INVx2_ASAP7_75t_L g6300 ( 
.A(n_6250),
.Y(n_6300)
);

OR2x2_ASAP7_75t_L g6301 ( 
.A(n_6280),
.B(n_6199),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_6263),
.Y(n_6302)
);

INVx2_ASAP7_75t_SL g6303 ( 
.A(n_6246),
.Y(n_6303)
);

OR2x2_ASAP7_75t_L g6304 ( 
.A(n_6285),
.B(n_6150),
.Y(n_6304)
);

AND2x2_ASAP7_75t_L g6305 ( 
.A(n_6257),
.B(n_6223),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6225),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_6236),
.Y(n_6307)
);

AND2x2_ASAP7_75t_L g6308 ( 
.A(n_6264),
.B(n_6222),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_6239),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_6271),
.B(n_6192),
.Y(n_6310)
);

INVx2_ASAP7_75t_L g6311 ( 
.A(n_6286),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_6283),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_6289),
.Y(n_6313)
);

AND2x4_ASAP7_75t_SL g6314 ( 
.A(n_6256),
.B(n_6224),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6292),
.Y(n_6315)
);

INVx3_ASAP7_75t_L g6316 ( 
.A(n_6277),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_6241),
.Y(n_6317)
);

INVx2_ASAP7_75t_L g6318 ( 
.A(n_6244),
.Y(n_6318)
);

NAND2x1_ASAP7_75t_L g6319 ( 
.A(n_6277),
.B(n_6198),
.Y(n_6319)
);

AND2x2_ASAP7_75t_L g6320 ( 
.A(n_6226),
.B(n_6196),
.Y(n_6320)
);

INVx2_ASAP7_75t_L g6321 ( 
.A(n_6249),
.Y(n_6321)
);

INVx2_ASAP7_75t_L g6322 ( 
.A(n_6253),
.Y(n_6322)
);

AND2x2_ASAP7_75t_L g6323 ( 
.A(n_6265),
.B(n_6188),
.Y(n_6323)
);

INVxp67_ASAP7_75t_L g6324 ( 
.A(n_6251),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_6254),
.Y(n_6325)
);

NAND2xp5_ASAP7_75t_L g6326 ( 
.A(n_6261),
.B(n_6198),
.Y(n_6326)
);

NAND3xp33_ASAP7_75t_L g6327 ( 
.A(n_6229),
.B(n_6260),
.C(n_6228),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_6282),
.Y(n_6328)
);

INVx2_ASAP7_75t_L g6329 ( 
.A(n_6278),
.Y(n_6329)
);

AND2x2_ASAP7_75t_L g6330 ( 
.A(n_6238),
.B(n_6181),
.Y(n_6330)
);

INVx2_ASAP7_75t_L g6331 ( 
.A(n_6278),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_6275),
.Y(n_6332)
);

INVx2_ASAP7_75t_L g6333 ( 
.A(n_6255),
.Y(n_6333)
);

INVx2_ASAP7_75t_L g6334 ( 
.A(n_6237),
.Y(n_6334)
);

AND2x2_ASAP7_75t_L g6335 ( 
.A(n_6243),
.B(n_6210),
.Y(n_6335)
);

HB1xp67_ASAP7_75t_L g6336 ( 
.A(n_6232),
.Y(n_6336)
);

AND2x2_ASAP7_75t_L g6337 ( 
.A(n_6245),
.B(n_6176),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_6232),
.Y(n_6338)
);

INVx2_ASAP7_75t_L g6339 ( 
.A(n_6284),
.Y(n_6339)
);

NAND2xp5_ASAP7_75t_L g6340 ( 
.A(n_6240),
.B(n_6180),
.Y(n_6340)
);

AND2x2_ASAP7_75t_L g6341 ( 
.A(n_6293),
.B(n_6308),
.Y(n_6341)
);

HB1xp67_ASAP7_75t_L g6342 ( 
.A(n_6294),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_6294),
.Y(n_6343)
);

AND2x4_ASAP7_75t_L g6344 ( 
.A(n_6314),
.B(n_6266),
.Y(n_6344)
);

INVxp67_ASAP7_75t_L g6345 ( 
.A(n_6297),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_6296),
.B(n_6297),
.Y(n_6346)
);

INVx2_ASAP7_75t_L g6347 ( 
.A(n_6319),
.Y(n_6347)
);

INVx2_ASAP7_75t_L g6348 ( 
.A(n_6316),
.Y(n_6348)
);

AND2x2_ASAP7_75t_L g6349 ( 
.A(n_6305),
.B(n_6242),
.Y(n_6349)
);

OAI21xp5_ASAP7_75t_L g6350 ( 
.A1(n_6327),
.A2(n_6233),
.B(n_6262),
.Y(n_6350)
);

OR2x2_ASAP7_75t_L g6351 ( 
.A(n_6304),
.B(n_6287),
.Y(n_6351)
);

NAND2xp5_ASAP7_75t_L g6352 ( 
.A(n_6299),
.B(n_6234),
.Y(n_6352)
);

OR2x2_ASAP7_75t_L g6353 ( 
.A(n_6301),
.B(n_6326),
.Y(n_6353)
);

NAND2xp5_ASAP7_75t_L g6354 ( 
.A(n_6300),
.B(n_6235),
.Y(n_6354)
);

INVx1_ASAP7_75t_SL g6355 ( 
.A(n_6314),
.Y(n_6355)
);

INVx1_ASAP7_75t_L g6356 ( 
.A(n_6336),
.Y(n_6356)
);

AND2x2_ASAP7_75t_L g6357 ( 
.A(n_6298),
.B(n_6247),
.Y(n_6357)
);

AOI22xp33_ASAP7_75t_L g6358 ( 
.A1(n_6303),
.A2(n_6258),
.B1(n_6259),
.B2(n_6268),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_L g6359 ( 
.A(n_6328),
.B(n_6270),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_6310),
.B(n_6190),
.Y(n_6360)
);

AND2x2_ASAP7_75t_L g6361 ( 
.A(n_6320),
.B(n_6291),
.Y(n_6361)
);

NAND2xp5_ASAP7_75t_L g6362 ( 
.A(n_6329),
.B(n_6252),
.Y(n_6362)
);

AND2x4_ASAP7_75t_L g6363 ( 
.A(n_6333),
.B(n_6212),
.Y(n_6363)
);

AND2x4_ASAP7_75t_L g6364 ( 
.A(n_6329),
.B(n_6215),
.Y(n_6364)
);

AND2x2_ASAP7_75t_L g6365 ( 
.A(n_6323),
.B(n_6330),
.Y(n_6365)
);

NAND2xp5_ASAP7_75t_L g6366 ( 
.A(n_6331),
.B(n_6219),
.Y(n_6366)
);

AND2x4_ASAP7_75t_L g6367 ( 
.A(n_6311),
.B(n_6220),
.Y(n_6367)
);

OR2x2_ASAP7_75t_L g6368 ( 
.A(n_6312),
.B(n_6338),
.Y(n_6368)
);

INVxp67_ASAP7_75t_L g6369 ( 
.A(n_6295),
.Y(n_6369)
);

INVxp67_ASAP7_75t_SL g6370 ( 
.A(n_6342),
.Y(n_6370)
);

NAND4xp75_ASAP7_75t_L g6371 ( 
.A(n_6350),
.B(n_6313),
.C(n_6315),
.D(n_6302),
.Y(n_6371)
);

AND2x2_ASAP7_75t_L g6372 ( 
.A(n_6341),
.B(n_6324),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_6355),
.B(n_6324),
.Y(n_6373)
);

AND2x2_ASAP7_75t_L g6374 ( 
.A(n_6355),
.B(n_6335),
.Y(n_6374)
);

AND2x2_ASAP7_75t_L g6375 ( 
.A(n_6349),
.B(n_6337),
.Y(n_6375)
);

NAND2xp5_ASAP7_75t_L g6376 ( 
.A(n_6344),
.B(n_6318),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_6353),
.Y(n_6377)
);

XNOR2xp5_ASAP7_75t_L g6378 ( 
.A(n_6357),
.B(n_6290),
.Y(n_6378)
);

HB1xp67_ASAP7_75t_L g6379 ( 
.A(n_6343),
.Y(n_6379)
);

AND2x4_ASAP7_75t_L g6380 ( 
.A(n_6347),
.B(n_6318),
.Y(n_6380)
);

CKINVDCx6p67_ASAP7_75t_R g6381 ( 
.A(n_6368),
.Y(n_6381)
);

AND2x2_ASAP7_75t_L g6382 ( 
.A(n_6365),
.B(n_6334),
.Y(n_6382)
);

XOR2xp5_ASAP7_75t_L g6383 ( 
.A(n_6358),
.B(n_6340),
.Y(n_6383)
);

AND2x2_ASAP7_75t_L g6384 ( 
.A(n_6361),
.B(n_6339),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6351),
.Y(n_6385)
);

INVx2_ASAP7_75t_L g6386 ( 
.A(n_6348),
.Y(n_6386)
);

NAND2xp5_ASAP7_75t_L g6387 ( 
.A(n_6345),
.B(n_6321),
.Y(n_6387)
);

INVx2_ASAP7_75t_L g6388 ( 
.A(n_6356),
.Y(n_6388)
);

HB1xp67_ASAP7_75t_L g6389 ( 
.A(n_6346),
.Y(n_6389)
);

INVx2_ASAP7_75t_L g6390 ( 
.A(n_6363),
.Y(n_6390)
);

NOR3xp33_ASAP7_75t_L g6391 ( 
.A(n_6362),
.B(n_6322),
.C(n_6325),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6360),
.Y(n_6392)
);

NAND4xp75_ASAP7_75t_L g6393 ( 
.A(n_6354),
.B(n_6317),
.C(n_6306),
.D(n_6307),
.Y(n_6393)
);

INVx5_ASAP7_75t_L g6394 ( 
.A(n_6364),
.Y(n_6394)
);

NOR2xp33_ASAP7_75t_L g6395 ( 
.A(n_6369),
.B(n_6309),
.Y(n_6395)
);

OAI22xp33_ASAP7_75t_L g6396 ( 
.A1(n_6381),
.A2(n_6362),
.B1(n_6354),
.B2(n_6352),
.Y(n_6396)
);

OR2x6_ASAP7_75t_L g6397 ( 
.A(n_6382),
.B(n_6359),
.Y(n_6397)
);

AOI22xp5_ASAP7_75t_L g6398 ( 
.A1(n_6372),
.A2(n_6367),
.B1(n_6272),
.B2(n_6269),
.Y(n_6398)
);

AOI22xp5_ASAP7_75t_L g6399 ( 
.A1(n_6373),
.A2(n_6332),
.B1(n_6273),
.B2(n_6366),
.Y(n_6399)
);

AO221x2_ASAP7_75t_L g6400 ( 
.A1(n_6383),
.A2(n_6366),
.B1(n_6332),
.B2(n_6248),
.C(n_6288),
.Y(n_6400)
);

OAI22xp33_ASAP7_75t_L g6401 ( 
.A1(n_6394),
.A2(n_6279),
.B1(n_6276),
.B2(n_6281),
.Y(n_6401)
);

AND2x2_ASAP7_75t_L g6402 ( 
.A(n_6374),
.B(n_399),
.Y(n_6402)
);

INVx1_ASAP7_75t_L g6403 ( 
.A(n_6394),
.Y(n_6403)
);

NAND2xp5_ASAP7_75t_L g6404 ( 
.A(n_6380),
.B(n_400),
.Y(n_6404)
);

OAI221xp5_ASAP7_75t_L g6405 ( 
.A1(n_6391),
.A2(n_405),
.B1(n_402),
.B2(n_404),
.C(n_406),
.Y(n_6405)
);

NOR2x1p5_ASAP7_75t_L g6406 ( 
.A(n_6371),
.B(n_404),
.Y(n_6406)
);

OR2x2_ASAP7_75t_L g6407 ( 
.A(n_6376),
.B(n_406),
.Y(n_6407)
);

NOR2xp67_ASAP7_75t_L g6408 ( 
.A(n_6390),
.B(n_411),
.Y(n_6408)
);

OAI22xp33_ASAP7_75t_L g6409 ( 
.A1(n_6389),
.A2(n_414),
.B1(n_411),
.B2(n_412),
.Y(n_6409)
);

AO221x2_ASAP7_75t_L g6410 ( 
.A1(n_6392),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.C(n_420),
.Y(n_6410)
);

NAND2xp5_ASAP7_75t_L g6411 ( 
.A(n_6375),
.B(n_416),
.Y(n_6411)
);

NAND2xp5_ASAP7_75t_L g6412 ( 
.A(n_6384),
.B(n_422),
.Y(n_6412)
);

AOI22xp5_ASAP7_75t_L g6413 ( 
.A1(n_6377),
.A2(n_428),
.B1(n_424),
.B2(n_427),
.Y(n_6413)
);

NAND2xp5_ASAP7_75t_L g6414 ( 
.A(n_6388),
.B(n_424),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_6385),
.B(n_6391),
.Y(n_6415)
);

O2A1O1Ixp33_ASAP7_75t_L g6416 ( 
.A1(n_6396),
.A2(n_6370),
.B(n_6387),
.C(n_6379),
.Y(n_6416)
);

AND2x2_ASAP7_75t_L g6417 ( 
.A(n_6402),
.B(n_6386),
.Y(n_6417)
);

INVx2_ASAP7_75t_L g6418 ( 
.A(n_6403),
.Y(n_6418)
);

INVx1_ASAP7_75t_SL g6419 ( 
.A(n_6397),
.Y(n_6419)
);

INVx2_ASAP7_75t_L g6420 ( 
.A(n_6397),
.Y(n_6420)
);

AND2x2_ASAP7_75t_L g6421 ( 
.A(n_6406),
.B(n_6378),
.Y(n_6421)
);

OAI21xp33_ASAP7_75t_L g6422 ( 
.A1(n_6415),
.A2(n_6395),
.B(n_6393),
.Y(n_6422)
);

AND2x4_ASAP7_75t_L g6423 ( 
.A(n_6408),
.B(n_429),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6410),
.Y(n_6424)
);

NAND2xp5_ASAP7_75t_L g6425 ( 
.A(n_6400),
.B(n_430),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6410),
.Y(n_6426)
);

NAND2xp5_ASAP7_75t_L g6427 ( 
.A(n_6400),
.B(n_431),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6423),
.Y(n_6428)
);

INVx1_ASAP7_75t_L g6429 ( 
.A(n_6423),
.Y(n_6429)
);

INVx1_ASAP7_75t_SL g6430 ( 
.A(n_6419),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6416),
.Y(n_6431)
);

INVx3_ASAP7_75t_L g6432 ( 
.A(n_6420),
.Y(n_6432)
);

HB1xp67_ASAP7_75t_L g6433 ( 
.A(n_6424),
.Y(n_6433)
);

OR2x2_ASAP7_75t_L g6434 ( 
.A(n_6426),
.B(n_6411),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6417),
.Y(n_6435)
);

OAI22xp5_ASAP7_75t_L g6436 ( 
.A1(n_6425),
.A2(n_6398),
.B1(n_6399),
.B2(n_6412),
.Y(n_6436)
);

INVx2_ASAP7_75t_L g6437 ( 
.A(n_6418),
.Y(n_6437)
);

OR2x2_ASAP7_75t_L g6438 ( 
.A(n_6427),
.B(n_6407),
.Y(n_6438)
);

AO21x2_ASAP7_75t_L g6439 ( 
.A1(n_6422),
.A2(n_6404),
.B(n_6414),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6421),
.Y(n_6440)
);

INVxp67_ASAP7_75t_L g6441 ( 
.A(n_6428),
.Y(n_6441)
);

OAI22xp5_ASAP7_75t_L g6442 ( 
.A1(n_6431),
.A2(n_6401),
.B1(n_6405),
.B2(n_6413),
.Y(n_6442)
);

NAND2xp5_ASAP7_75t_L g6443 ( 
.A(n_6429),
.B(n_6409),
.Y(n_6443)
);

INVx1_ASAP7_75t_SL g6444 ( 
.A(n_6434),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6432),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6435),
.Y(n_6446)
);

BUFx8_ASAP7_75t_SL g6447 ( 
.A(n_6437),
.Y(n_6447)
);

OAI21xp5_ASAP7_75t_SL g6448 ( 
.A1(n_6440),
.A2(n_434),
.B(n_436),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_6438),
.Y(n_6449)
);

NAND3xp33_ASAP7_75t_L g6450 ( 
.A(n_6436),
.B(n_438),
.C(n_442),
.Y(n_6450)
);

OR2x2_ASAP7_75t_L g6451 ( 
.A(n_6439),
.B(n_446),
.Y(n_6451)
);

AND2x2_ASAP7_75t_L g6452 ( 
.A(n_6430),
.B(n_449),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_6433),
.Y(n_6453)
);

NAND2xp5_ASAP7_75t_L g6454 ( 
.A(n_6452),
.B(n_450),
.Y(n_6454)
);

NAND2xp5_ASAP7_75t_L g6455 ( 
.A(n_6445),
.B(n_451),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6451),
.Y(n_6456)
);

INVx3_ASAP7_75t_L g6457 ( 
.A(n_6447),
.Y(n_6457)
);

NOR2xp33_ASAP7_75t_L g6458 ( 
.A(n_6441),
.B(n_456),
.Y(n_6458)
);

NAND2x1p5_ASAP7_75t_L g6459 ( 
.A(n_6444),
.B(n_457),
.Y(n_6459)
);

AOI22xp5_ASAP7_75t_L g6460 ( 
.A1(n_6453),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_6460)
);

INVx1_ASAP7_75t_L g6461 ( 
.A(n_6443),
.Y(n_6461)
);

NAND2xp5_ASAP7_75t_L g6462 ( 
.A(n_6448),
.B(n_465),
.Y(n_6462)
);

OAI22xp5_ASAP7_75t_L g6463 ( 
.A1(n_6446),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_6463)
);

NAND2xp5_ASAP7_75t_L g6464 ( 
.A(n_6449),
.B(n_468),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_6450),
.Y(n_6465)
);

OAI221xp5_ASAP7_75t_L g6466 ( 
.A1(n_6442),
.A2(n_471),
.B1(n_472),
.B2(n_473),
.C(n_474),
.Y(n_6466)
);

OR2x2_ASAP7_75t_L g6467 ( 
.A(n_6459),
.B(n_479),
.Y(n_6467)
);

NAND2xp5_ASAP7_75t_L g6468 ( 
.A(n_6457),
.B(n_481),
.Y(n_6468)
);

NAND2x1_ASAP7_75t_SL g6469 ( 
.A(n_6456),
.B(n_482),
.Y(n_6469)
);

OR2x2_ASAP7_75t_L g6470 ( 
.A(n_6464),
.B(n_483),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_6454),
.Y(n_6471)
);

AOI22xp33_ASAP7_75t_L g6472 ( 
.A1(n_6461),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_6472)
);

NOR2xp33_ASAP7_75t_L g6473 ( 
.A(n_6466),
.B(n_485),
.Y(n_6473)
);

NAND2xp5_ASAP7_75t_L g6474 ( 
.A(n_6458),
.B(n_486),
.Y(n_6474)
);

AOI22xp33_ASAP7_75t_L g6475 ( 
.A1(n_6465),
.A2(n_490),
.B1(n_487),
.B2(n_488),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_6455),
.Y(n_6476)
);

INVx2_ASAP7_75t_L g6477 ( 
.A(n_6462),
.Y(n_6477)
);

INVx1_ASAP7_75t_SL g6478 ( 
.A(n_6460),
.Y(n_6478)
);

NAND2xp5_ASAP7_75t_L g6479 ( 
.A(n_6469),
.B(n_6463),
.Y(n_6479)
);

HB1xp67_ASAP7_75t_L g6480 ( 
.A(n_6467),
.Y(n_6480)
);

NOR2x1_ASAP7_75t_L g6481 ( 
.A(n_6468),
.B(n_499),
.Y(n_6481)
);

INVx1_ASAP7_75t_SL g6482 ( 
.A(n_6470),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_6474),
.Y(n_6483)
);

AND2x2_ASAP7_75t_L g6484 ( 
.A(n_6478),
.B(n_506),
.Y(n_6484)
);

INVx1_ASAP7_75t_SL g6485 ( 
.A(n_6471),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_6481),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6484),
.Y(n_6487)
);

INVx2_ASAP7_75t_SL g6488 ( 
.A(n_6479),
.Y(n_6488)
);

INVx1_ASAP7_75t_L g6489 ( 
.A(n_6480),
.Y(n_6489)
);

INVxp33_ASAP7_75t_SL g6490 ( 
.A(n_6485),
.Y(n_6490)
);

OAI22xp5_ASAP7_75t_L g6491 ( 
.A1(n_6490),
.A2(n_6473),
.B1(n_6482),
.B2(n_6477),
.Y(n_6491)
);

AOI221xp5_ASAP7_75t_L g6492 ( 
.A1(n_6489),
.A2(n_6476),
.B1(n_6483),
.B2(n_6472),
.C(n_6475),
.Y(n_6492)
);

OAI22xp5_ASAP7_75t_L g6493 ( 
.A1(n_6488),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.Y(n_6493)
);

AO22x2_ASAP7_75t_L g6494 ( 
.A1(n_6487),
.A2(n_515),
.B1(n_516),
.B2(n_518),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_6486),
.Y(n_6495)
);

NAND4xp25_ASAP7_75t_SL g6496 ( 
.A(n_6492),
.B(n_533),
.C(n_534),
.D(n_535),
.Y(n_6496)
);

AOI222xp33_ASAP7_75t_L g6497 ( 
.A1(n_6495),
.A2(n_538),
.B1(n_541),
.B2(n_542),
.C1(n_543),
.C2(n_544),
.Y(n_6497)
);

AOI211xp5_ASAP7_75t_L g6498 ( 
.A1(n_6491),
.A2(n_542),
.B(n_543),
.C(n_544),
.Y(n_6498)
);

AOI22xp33_ASAP7_75t_L g6499 ( 
.A1(n_6493),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_6499)
);

NAND2xp33_ASAP7_75t_R g6500 ( 
.A(n_6494),
.B(n_552),
.Y(n_6500)
);

HB1xp67_ASAP7_75t_L g6501 ( 
.A(n_6500),
.Y(n_6501)
);

OR2x2_ASAP7_75t_L g6502 ( 
.A(n_6496),
.B(n_558),
.Y(n_6502)
);

NAND3xp33_ASAP7_75t_L g6503 ( 
.A(n_6498),
.B(n_563),
.C(n_564),
.Y(n_6503)
);

NAND3xp33_ASAP7_75t_L g6504 ( 
.A(n_6499),
.B(n_570),
.C(n_573),
.Y(n_6504)
);

AND2x2_ASAP7_75t_L g6505 ( 
.A(n_6501),
.B(n_6497),
.Y(n_6505)
);

AOI22xp5_ASAP7_75t_L g6506 ( 
.A1(n_6505),
.A2(n_6504),
.B1(n_6503),
.B2(n_6502),
.Y(n_6506)
);

INVx1_ASAP7_75t_L g6507 ( 
.A(n_6506),
.Y(n_6507)
);

HB1xp67_ASAP7_75t_L g6508 ( 
.A(n_6507),
.Y(n_6508)
);

HB1xp67_ASAP7_75t_L g6509 ( 
.A(n_6508),
.Y(n_6509)
);

CKINVDCx5p33_ASAP7_75t_R g6510 ( 
.A(n_6509),
.Y(n_6510)
);

HB1xp67_ASAP7_75t_L g6511 ( 
.A(n_6510),
.Y(n_6511)
);

NAND3xp33_ASAP7_75t_L g6512 ( 
.A(n_6511),
.B(n_596),
.C(n_597),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_6512),
.Y(n_6513)
);

OAI22xp5_ASAP7_75t_L g6514 ( 
.A1(n_6513),
.A2(n_616),
.B1(n_617),
.B2(n_618),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_6514),
.Y(n_6515)
);

OAI21x1_ASAP7_75t_L g6516 ( 
.A1(n_6515),
.A2(n_1908),
.B(n_1977),
.Y(n_6516)
);

AOI22xp5_ASAP7_75t_L g6517 ( 
.A1(n_6516),
.A2(n_1953),
.B1(n_1977),
.B2(n_2601),
.Y(n_6517)
);

AO22x1_ASAP7_75t_L g6518 ( 
.A1(n_6517),
.A2(n_2001),
.B1(n_1973),
.B2(n_1980),
.Y(n_6518)
);

INVx2_ASAP7_75t_L g6519 ( 
.A(n_6518),
.Y(n_6519)
);

INVx1_ASAP7_75t_SL g6520 ( 
.A(n_6519),
.Y(n_6520)
);

AOI21xp33_ASAP7_75t_L g6521 ( 
.A1(n_6520),
.A2(n_2007),
.B(n_1980),
.Y(n_6521)
);

OA22x2_ASAP7_75t_L g6522 ( 
.A1(n_6520),
.A2(n_1950),
.B1(n_2021),
.B2(n_2043),
.Y(n_6522)
);

AOI221xp5_ASAP7_75t_SL g6523 ( 
.A1(n_6521),
.A2(n_1980),
.B1(n_2001),
.B2(n_1968),
.C(n_1950),
.Y(n_6523)
);

AOI21xp33_ASAP7_75t_L g6524 ( 
.A1(n_6523),
.A2(n_6522),
.B(n_2001),
.Y(n_6524)
);

AOI211xp5_ASAP7_75t_L g6525 ( 
.A1(n_6524),
.A2(n_1968),
.B(n_2579),
.C(n_2955),
.Y(n_6525)
);


endmodule