module real_jpeg_4298_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_1),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_1),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_1),
.Y(n_141)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_1),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_1),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_1),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_2),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_117),
.B1(n_147),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_2),
.A2(n_147),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_2),
.A2(n_147),
.B1(n_174),
.B2(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_3),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_3),
.A2(n_260),
.B1(n_290),
.B2(n_294),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_307),
.C(n_311),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_3),
.B(n_98),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_3),
.B(n_44),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_3),
.B(n_84),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_3),
.B(n_382),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_6),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_6),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_6),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_7),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_7),
.A2(n_39),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_58),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_8),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_8),
.A2(n_81),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_8),
.A2(n_81),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_9),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_9),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_64),
.B1(n_109),
.B2(n_158),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_9),
.A2(n_109),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_9),
.A2(n_109),
.B1(n_388),
.B2(n_392),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_10),
.A2(n_46),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_12),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_12),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_57),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_13),
.A2(n_57),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_14),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_14),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_14),
.A2(n_142),
.B1(n_208),
.B2(n_277),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_14),
.A2(n_142),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_14),
.A2(n_142),
.B1(n_290),
.B2(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_15),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_15),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_15),
.A2(n_58),
.B1(n_187),
.B2(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_15),
.A2(n_187),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_15),
.A2(n_187),
.B1(n_249),
.B2(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_234),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_233),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_198),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_20),
.B(n_198),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_152),
.C(n_165),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_21),
.B(n_152),
.CI(n_165),
.CON(n_279),
.SN(n_279)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_85),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_22),
.B(n_86),
.C(n_119),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_23),
.B(n_51),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_33),
.B1(n_42),
.B2(n_45),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_24),
.A2(n_45),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_24),
.A2(n_43),
.B1(n_266),
.B2(n_273),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_24),
.A2(n_317),
.B(n_324),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_24),
.A2(n_260),
.B(n_324),
.Y(n_345)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_25),
.A2(n_173),
.B1(n_179),
.B2(n_180),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_25),
.B(n_327),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_25),
.A2(n_325),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_25),
.A2(n_267),
.B1(n_387),
.B2(n_422),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_28),
.Y(n_181)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_28),
.Y(n_423)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_32),
.Y(n_268)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_33),
.Y(n_179)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_37),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_40),
.Y(n_349)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_50),
.Y(n_323)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_50),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_80),
.B2(n_84),
.Y(n_51)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_52),
.Y(n_171)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_56),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_56),
.Y(n_399)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_60),
.Y(n_160)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_60),
.Y(n_218)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_60),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_61),
.A2(n_80),
.B1(n_84),
.B2(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_61),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_61),
.A2(n_84),
.B1(n_155),
.B2(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_61),
.B(n_297),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_67),
.B2(n_69),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_66),
.Y(n_310)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_71),
.A2(n_332),
.B(n_335),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_76),
.Y(n_314)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_76),
.Y(n_391)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_99),
.B1(n_102),
.B2(n_105),
.Y(n_98)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_84),
.B(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_119),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_87),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_87),
.A2(n_112),
.B1(n_276),
.B2(n_416),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_90),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_93),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_93),
.Y(n_379)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_94),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_94),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_94),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_94),
.Y(n_383)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_95),
.Y(n_405)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22x1_ASAP7_75t_L g192 ( 
.A1(n_98),
.A2(n_193),
.B1(n_194),
.B2(n_197),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_98),
.A2(n_193),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_104),
.Y(n_373)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_112),
.B(n_195),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_112),
.A2(n_416),
.B(n_418),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g398 ( 
.A1(n_116),
.A2(n_381),
.A3(n_399),
.B1(n_400),
.B2(n_403),
.Y(n_398)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_139),
.B(n_145),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_133),
.B1(n_139),
.B2(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_121),
.B(n_146),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_121),
.A2(n_438),
.B(n_439),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_133),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_126),
.B1(n_129),
.B2(n_131),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_132),
.Y(n_255)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_133),
.B(n_260),
.Y(n_420)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g196 ( 
.A(n_136),
.Y(n_196)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_145),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_151),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_161),
.B2(n_164),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_161),
.Y(n_222)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_160),
.Y(n_295)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_161),
.A2(n_164),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_182),
.C(n_192),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_166),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_167),
.B(n_172),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_168),
.A2(n_289),
.B(n_296),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_168),
.A2(n_170),
.B1(n_332),
.B2(n_370),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_168),
.A2(n_296),
.B(n_370),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_169),
.A2(n_170),
.B(n_335),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_178),
.Y(n_343)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_182),
.A2(n_183),
.B1(n_192),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_184),
.A2(n_232),
.B(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_193),
.A2(n_275),
.B(n_278),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_193),
.A2(n_278),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_193),
.B(n_194),
.Y(n_418)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_196),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_220),
.B2(n_221),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_212),
.B(n_219),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_213),
.Y(n_219)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_218),
.Y(n_305)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g438 ( 
.A1(n_228),
.A2(n_259),
.B(n_260),
.Y(n_438)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_280),
.B(n_467),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_279),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_237),
.B(n_279),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_242),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_243),
.B(n_457),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.C(n_274),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_244),
.A2(n_245),
.B1(n_274),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_247),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_264),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_248),
.A2(n_264),
.B1(n_265),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_248),
.Y(n_431)
);

OAI32xp33_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.A3(n_252),
.B1(n_254),
.B2(n_259),
.Y(n_248)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_SL g376 ( 
.A1(n_260),
.A2(n_377),
.B(n_380),
.Y(n_376)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_274),
.Y(n_452)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_279),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_445),
.B(n_464),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_426),
.B(n_444),
.Y(n_282)
);

AO21x1_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_407),
.B(n_425),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_364),
.B(n_406),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_338),
.B(n_363),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_315),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_287),
.B(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_301),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_288),
.A2(n_301),
.B1(n_302),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

INVx5_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_329),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_330),
.C(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_336),
.B2(n_337),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_SL g403 ( 
.A(n_333),
.B(n_404),
.Y(n_403)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_356),
.B(n_362),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_346),
.B(n_355),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_354),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_352),
.B(n_353),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_348),
.Y(n_358)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_386),
.B(n_395),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_360),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_366),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_384),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_374),
.B2(n_375),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_374),
.C(n_384),
.Y(n_408)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_398),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_398),
.Y(n_413)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_408),
.B(n_409),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B1(n_414),
.B2(n_424),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_413),
.C(n_424),
.Y(n_427)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_414),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_419),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_420),
.C(n_421),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_427),
.B(n_428),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_435),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_432),
.B1(n_433),
.B2(n_434),
.Y(n_429)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_432),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_433),
.C(n_435),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_440),
.B2(n_443),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_441),
.C(n_442),
.Y(n_455)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_440),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_459),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_465),
.B(n_466),
.Y(n_464)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_456),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_456),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_453),
.C(n_455),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_462),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_453),
.A2(n_454),
.B1(n_455),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_455),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_461),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);


endmodule