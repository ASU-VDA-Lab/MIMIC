module real_aes_7835_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g497 ( .A(n_1), .Y(n_497) );
INVx1_ASAP7_75t_L g203 ( .A(n_2), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_3), .A2(n_38), .B1(n_164), .B2(n_527), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g171 ( .A1(n_4), .A2(n_145), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_5), .B(n_138), .Y(n_510) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_7), .A2(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_8), .B(n_39), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_8), .B(n_39), .Y(n_462) );
INVx1_ASAP7_75t_L g178 ( .A(n_9), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_10), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g143 ( .A(n_11), .Y(n_143) );
INVx1_ASAP7_75t_L g491 ( .A(n_12), .Y(n_491) );
INVx1_ASAP7_75t_L g259 ( .A(n_13), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_14), .B(n_186), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_15), .B(n_139), .Y(n_568) );
AO32x2_ASAP7_75t_L g540 ( .A1(n_16), .A2(n_138), .A3(n_183), .B1(n_519), .B2(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_17), .A2(n_63), .B1(n_127), .B2(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_17), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_18), .B(n_164), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_19), .B(n_159), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_20), .B(n_139), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_21), .A2(n_51), .B1(n_164), .B2(n_527), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_22), .B(n_145), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_23), .A2(n_80), .B1(n_164), .B2(n_186), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_24), .B(n_164), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_25), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_26), .A2(n_257), .B(n_258), .C(n_260), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_27), .A2(n_105), .B1(n_113), .B2(n_776), .Y(n_104) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_29), .B(n_180), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_30), .B(n_176), .Y(n_205) );
INVx1_ASAP7_75t_L g192 ( .A(n_31), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_32), .A2(n_33), .B1(n_121), .B2(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_32), .Y(n_122) );
INVxp67_ASAP7_75t_L g121 ( .A(n_33), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_33), .B(n_180), .Y(n_557) );
INVx2_ASAP7_75t_L g148 ( .A(n_34), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_35), .B(n_164), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_36), .B(n_180), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_37), .A2(n_150), .B(n_154), .C(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g190 ( .A(n_40), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_41), .A2(n_470), .B1(n_473), .B2(n_474), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_41), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_42), .B(n_176), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_43), .B(n_164), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_44), .A2(n_90), .B1(n_222), .B2(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_45), .B(n_164), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_46), .B(n_164), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_47), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_48), .A2(n_70), .B1(n_471), .B2(n_472), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_48), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_49), .B(n_496), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_50), .B(n_145), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_52), .A2(n_61), .B1(n_164), .B2(n_186), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_53), .A2(n_154), .B1(n_186), .B2(n_188), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_54), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_55), .B(n_164), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_56), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_57), .B(n_164), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_58), .A2(n_163), .B(n_175), .C(n_177), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_59), .Y(n_235) );
INVx1_ASAP7_75t_L g173 ( .A(n_60), .Y(n_173) );
INVx1_ASAP7_75t_L g151 ( .A(n_62), .Y(n_151) );
INVx1_ASAP7_75t_L g127 ( .A(n_63), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_64), .B(n_164), .Y(n_498) );
INVx1_ASAP7_75t_L g142 ( .A(n_65), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
AO32x2_ASAP7_75t_L g524 ( .A1(n_67), .A2(n_138), .A3(n_239), .B1(n_519), .B2(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g517 ( .A(n_68), .Y(n_517) );
INVx1_ASAP7_75t_L g552 ( .A(n_69), .Y(n_552) );
INVx1_ASAP7_75t_L g471 ( .A(n_70), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_SL g158 ( .A1(n_71), .A2(n_159), .B(n_160), .C(n_163), .Y(n_158) );
INVxp67_ASAP7_75t_L g161 ( .A(n_72), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_73), .B(n_186), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_74), .A2(n_468), .B1(n_469), .B2(n_475), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_74), .Y(n_468) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_76), .B(n_458), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_77), .A2(n_460), .B1(n_466), .B2(n_771), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_78), .Y(n_196) );
INVx1_ASAP7_75t_L g228 ( .A(n_79), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_81), .A2(n_150), .B(n_154), .C(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_82), .B(n_527), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_83), .B(n_186), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_84), .B(n_204), .Y(n_218) );
INVx2_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_86), .B(n_159), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_87), .B(n_186), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_88), .A2(n_150), .B(n_154), .C(n_202), .Y(n_201) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_89), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g459 ( .A(n_89), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g477 ( .A(n_89), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_91), .A2(n_103), .B1(n_186), .B2(n_187), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_92), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_93), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_94), .A2(n_150), .B(n_154), .C(n_242), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_95), .Y(n_249) );
INVx1_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_97), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_98), .B(n_204), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_99), .B(n_186), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_100), .B(n_138), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_101), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_102), .A2(n_145), .B(n_152), .Y(n_144) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g776 ( .A(n_106), .Y(n_776) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g461 ( .A(n_109), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_464), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g775 ( .A(n_117), .Y(n_775) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_456), .B(n_463), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B1(n_124), .B2(n_455), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_120), .Y(n_455) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_454), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g454 ( .A(n_129), .Y(n_454) );
AOI22xp5_ASAP7_75t_SL g476 ( .A1(n_129), .A2(n_477), .B1(n_478), .B2(n_770), .Y(n_476) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND4x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_372), .C(n_419), .D(n_439), .Y(n_130) );
NOR3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_302), .C(n_327), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_210), .B(n_262), .C(n_292), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_181), .Y(n_134) );
INVx3_ASAP7_75t_SL g344 ( .A(n_135), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_135), .B(n_275), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_135), .B(n_197), .Y(n_425) );
AND2x2_ASAP7_75t_L g448 ( .A(n_135), .B(n_314), .Y(n_448) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_169), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g266 ( .A(n_137), .B(n_170), .Y(n_266) );
INVx3_ASAP7_75t_L g279 ( .A(n_137), .Y(n_279) );
AND2x2_ASAP7_75t_L g284 ( .A(n_137), .B(n_169), .Y(n_284) );
OR2x2_ASAP7_75t_L g335 ( .A(n_137), .B(n_276), .Y(n_335) );
BUFx2_ASAP7_75t_L g355 ( .A(n_137), .Y(n_355) );
AND2x2_ASAP7_75t_L g365 ( .A(n_137), .B(n_276), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_137), .B(n_182), .Y(n_371) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_166), .Y(n_137) );
INVx4_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_138), .A2(n_503), .B(n_510), .Y(n_502) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_140), .B(n_141), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx2_ASAP7_75t_L g253 ( .A(n_145), .Y(n_253) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_146), .B(n_150), .Y(n_194) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g496 ( .A(n_147), .Y(n_496) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g155 ( .A(n_148), .Y(n_155) );
INVx1_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
INVx4_ASAP7_75t_SL g165 ( .A(n_150), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_150), .A2(n_490), .B(n_494), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_150), .A2(n_504), .B(n_507), .Y(n_503) );
BUFx3_ASAP7_75t_L g519 ( .A(n_150), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_150), .A2(n_532), .B(n_536), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_150), .A2(n_551), .B(n_554), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B(n_158), .C(n_165), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_165), .B(n_173), .C(n_174), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_153), .A2(n_165), .B(n_255), .C(n_256), .Y(n_254) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_155), .Y(n_164) );
BUFx3_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
INVx1_ASAP7_75t_L g527 ( .A(n_155), .Y(n_527) );
INVx1_ASAP7_75t_L g535 ( .A(n_159), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_162), .B(n_178), .Y(n_177) );
INVx5_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
OAI22xp5_ASAP7_75t_SL g525 ( .A1(n_162), .A2(n_176), .B1(n_526), .B2(n_528), .Y(n_525) );
O2A1O1Ixp5_ASAP7_75t_SL g551 ( .A1(n_163), .A2(n_204), .B(n_552), .C(n_553), .Y(n_551) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_164), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_165), .A2(n_185), .B1(n_193), .B2(n_194), .Y(n_184) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_167), .A2(n_171), .B(n_179), .Y(n_170) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_168), .B(n_225), .Y(n_224) );
AO21x1_ASAP7_75t_L g563 ( .A1(n_168), .A2(n_564), .B(n_567), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g582 ( .A(n_168), .B(n_519), .C(n_564), .Y(n_582) );
INVx1_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_170), .B(n_276), .Y(n_290) );
INVx2_ASAP7_75t_L g300 ( .A(n_170), .Y(n_300) );
AND2x2_ASAP7_75t_L g313 ( .A(n_170), .B(n_279), .Y(n_313) );
OR2x2_ASAP7_75t_L g324 ( .A(n_170), .B(n_276), .Y(n_324) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_170), .B(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g382 ( .A(n_170), .Y(n_382) );
AND2x2_ASAP7_75t_L g428 ( .A(n_170), .B(n_182), .Y(n_428) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_175), .A2(n_495), .B(n_517), .C(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_175), .A2(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g245 ( .A(n_176), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_176), .A2(n_499), .B1(n_542), .B2(n_543), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_176), .A2(n_499), .B1(n_565), .B2(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
INVx2_ASAP7_75t_L g239 ( .A(n_180), .Y(n_239) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_180), .A2(n_252), .B(n_261), .Y(n_251) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_180), .A2(n_531), .B(n_539), .Y(n_530) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_180), .A2(n_550), .B(n_557), .Y(n_549) );
INVx3_ASAP7_75t_SL g301 ( .A(n_181), .Y(n_301) );
OR2x2_ASAP7_75t_L g354 ( .A(n_181), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_197), .Y(n_181) );
INVx3_ASAP7_75t_L g276 ( .A(n_182), .Y(n_276) );
AND2x2_ASAP7_75t_L g343 ( .A(n_182), .B(n_198), .Y(n_343) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_182), .Y(n_411) );
AOI33xp33_ASAP7_75t_L g415 ( .A1(n_182), .A2(n_344), .A3(n_351), .B1(n_360), .B2(n_416), .B3(n_417), .Y(n_415) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_195), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_183), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_183), .A2(n_199), .B(n_207), .Y(n_198) );
INVx2_ASAP7_75t_L g223 ( .A(n_183), .Y(n_223) );
INVx2_ASAP7_75t_L g206 ( .A(n_186), .Y(n_206) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_189), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_188) );
INVx2_ASAP7_75t_L g191 ( .A(n_189), .Y(n_191) );
INVx4_ASAP7_75t_L g257 ( .A(n_189), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_194), .A2(n_200), .B(n_201), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_194), .A2(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g264 ( .A(n_197), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
NOR3xp33_ASAP7_75t_L g338 ( .A(n_197), .B(n_339), .C(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g364 ( .A(n_197), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_197), .B(n_371), .Y(n_374) );
AND2x2_ASAP7_75t_L g427 ( .A(n_197), .B(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g283 ( .A(n_198), .Y(n_283) );
OR2x2_ASAP7_75t_L g377 ( .A(n_198), .B(n_276), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .C(n_206), .Y(n_202) );
INVx2_ASAP7_75t_L g499 ( .A(n_204), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_204), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_204), .A2(n_514), .B(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_206), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_209), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_209), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_236), .Y(n_210) );
AOI32xp33_ASAP7_75t_L g328 ( .A1(n_211), .A2(n_329), .A3(n_331), .B1(n_333), .B2(n_336), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_211), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g431 ( .A(n_211), .Y(n_431) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g363 ( .A(n_212), .B(n_347), .Y(n_363) );
AND2x2_ASAP7_75t_L g383 ( .A(n_212), .B(n_309), .Y(n_383) );
AND2x2_ASAP7_75t_L g451 ( .A(n_212), .B(n_369), .Y(n_451) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
INVx3_ASAP7_75t_L g272 ( .A(n_213), .Y(n_272) );
AND2x2_ASAP7_75t_L g286 ( .A(n_213), .B(n_270), .Y(n_286) );
OR2x2_ASAP7_75t_L g291 ( .A(n_213), .B(n_269), .Y(n_291) );
INVx1_ASAP7_75t_L g298 ( .A(n_213), .Y(n_298) );
AND2x2_ASAP7_75t_L g306 ( .A(n_213), .B(n_280), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_213), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_213), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g361 ( .A(n_213), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_213), .B(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_216), .B(n_223), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_220), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g260 ( .A(n_222), .Y(n_260) );
INVx1_ASAP7_75t_L g233 ( .A(n_223), .Y(n_233) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_223), .A2(n_489), .B(n_500), .Y(n_488) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_223), .A2(n_512), .B(n_520), .Y(n_511) );
INVx2_ASAP7_75t_L g270 ( .A(n_226), .Y(n_270) );
AND2x2_ASAP7_75t_L g316 ( .A(n_226), .B(n_237), .Y(n_316) );
AND2x2_ASAP7_75t_L g326 ( .A(n_226), .B(n_251), .Y(n_326) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_233), .B(n_234), .Y(n_226) );
INVx2_ASAP7_75t_L g446 ( .A(n_236), .Y(n_446) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_250), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_237), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
AND2x2_ASAP7_75t_L g331 ( .A(n_237), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g347 ( .A(n_237), .B(n_310), .Y(n_347) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g295 ( .A(n_238), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_238), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g360 ( .A(n_238), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_238), .B(n_270), .Y(n_392) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_248), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_246), .Y(n_242) );
AND2x2_ASAP7_75t_L g271 ( .A(n_250), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g332 ( .A(n_250), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_250), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g369 ( .A(n_250), .Y(n_369) );
INVx1_ASAP7_75t_L g402 ( .A(n_250), .Y(n_402) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g280 ( .A(n_251), .B(n_270), .Y(n_280) );
INVx1_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_257), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g493 ( .A(n_257), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_257), .A2(n_555), .B(n_556), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B1(n_273), .B2(n_280), .C(n_281), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_264), .B(n_284), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_264), .B(n_347), .Y(n_424) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_266), .B(n_314), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_266), .B(n_275), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_266), .B(n_289), .Y(n_418) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g340 ( .A(n_270), .Y(n_340) );
AND2x2_ASAP7_75t_L g315 ( .A(n_271), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g393 ( .A(n_271), .Y(n_393) );
AND2x2_ASAP7_75t_L g325 ( .A(n_272), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_272), .B(n_295), .Y(n_341) );
AND2x2_ASAP7_75t_L g405 ( .A(n_272), .B(n_331), .Y(n_405) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g314 ( .A(n_276), .B(n_283), .Y(n_314) );
AND2x2_ASAP7_75t_L g410 ( .A(n_277), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_279), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_280), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_280), .B(n_287), .Y(n_375) );
AND2x2_ASAP7_75t_L g395 ( .A(n_280), .B(n_295), .Y(n_395) );
AND2x2_ASAP7_75t_L g416 ( .A(n_280), .B(n_360), .Y(n_416) );
OAI32xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .A3(n_287), .B1(n_288), .B2(n_291), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_SL g289 ( .A(n_283), .Y(n_289) );
NAND2x1_ASAP7_75t_L g330 ( .A(n_283), .B(n_313), .Y(n_330) );
OR2x2_ASAP7_75t_L g334 ( .A(n_283), .B(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_283), .B(n_382), .Y(n_435) );
INVx1_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_285), .A2(n_376), .B1(n_422), .B2(n_425), .C(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_286), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g336 ( .A(n_286), .B(n_309), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_286), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g414 ( .A(n_286), .B(n_347), .Y(n_414) );
INVxp67_ASAP7_75t_L g350 ( .A(n_287), .Y(n_350) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g420 ( .A(n_289), .B(n_407), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_289), .B(n_370), .Y(n_443) );
INVx1_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_291), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g436 ( .A(n_291), .B(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_296), .B(n_299), .Y(n_292) );
AND2x2_ASAP7_75t_L g305 ( .A(n_294), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g389 ( .A(n_298), .B(n_309), .Y(n_389) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g407 ( .A(n_300), .B(n_365), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_300), .B(n_364), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_301), .B(n_313), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_307), .C(n_317), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_303), .A2(n_338), .B1(n_342), .B2(n_345), .C(n_348), .Y(n_337) );
AOI31xp33_ASAP7_75t_L g432 ( .A1(n_303), .A2(n_433), .A3(n_434), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_313), .B2(n_315), .Y(n_307) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g433 ( .A(n_313), .Y(n_433) );
INVx1_ASAP7_75t_L g396 ( .A(n_314), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_316), .A2(n_440), .B(n_442), .C(n_444), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_321), .B2(n_325), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_322), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_324), .A2(n_358), .B1(n_377), .B2(n_413), .C(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g408 ( .A(n_325), .Y(n_408) );
INVx1_ASAP7_75t_L g362 ( .A(n_326), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g327 ( .A(n_328), .B(n_337), .C(n_352), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g378 ( .A1(n_329), .A2(n_379), .B(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_331), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g438 ( .A(n_332), .Y(n_438) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g376 ( .A(n_339), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g351 ( .A(n_340), .Y(n_351) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g349 ( .A(n_343), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_343), .B(n_381), .Y(n_380) );
NOR4xp25_ASAP7_75t_L g348 ( .A(n_344), .B(n_349), .C(n_350), .D(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_357), .B1(n_363), .B2(n_364), .C1(n_366), .C2(n_370), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g450 ( .A(n_354), .Y(n_450) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_366), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_371), .A2(n_427), .B(n_429), .Y(n_426) );
NOR4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_384), .C(n_397), .D(n_412), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_377), .C(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g453 ( .A(n_374), .Y(n_453) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_381), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B1(n_390), .B2(n_391), .C1(n_394), .C2(n_396), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_389), .A2(n_420), .B(n_421), .C(n_432), .Y(n_419) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OAI222xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_403), .B1(n_404), .B2(n_406), .C1(n_408), .C2(n_409), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_414), .A2(n_417), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI211xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_447), .B(n_449), .C(n_452), .Y(n_444) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR2x2_ASAP7_75t_L g773 ( .A(n_460), .B(n_477), .Y(n_773) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_463), .A2(n_465), .B(n_774), .Y(n_464) );
XNOR2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
INVx1_ASAP7_75t_L g475 ( .A(n_469), .Y(n_475) );
INVx1_ASAP7_75t_L g473 ( .A(n_470), .Y(n_473) );
INVx2_ASAP7_75t_L g770 ( .A(n_477), .Y(n_770) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_480), .B(n_736), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_640), .C(n_724), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_583), .C(n_605), .D(n_621), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_521), .B1(n_544), .B2(n_562), .C(n_569), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_501), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_485), .B(n_562), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_485), .B(n_623), .C(n_636), .D(n_638), .Y(n_635) );
INVxp67_ASAP7_75t_L g752 ( .A(n_485), .Y(n_752) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g634 ( .A(n_486), .B(n_572), .Y(n_634) );
AND2x2_ASAP7_75t_L g658 ( .A(n_486), .B(n_501), .Y(n_658) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g625 ( .A(n_487), .B(n_561), .Y(n_625) );
AND2x2_ASAP7_75t_L g665 ( .A(n_487), .B(n_646), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_487), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_487), .B(n_502), .Y(n_706) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g560 ( .A(n_488), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g577 ( .A(n_488), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g589 ( .A(n_488), .B(n_502), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_488), .B(n_511), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_497), .B(n_498), .C(n_499), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_499), .A2(n_508), .B(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_L g592 ( .A(n_501), .B(n_593), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_501), .A2(n_642), .B1(n_645), .B2(n_647), .C(n_651), .Y(n_641) );
AND2x2_ASAP7_75t_L g700 ( .A(n_501), .B(n_665), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_501), .B(n_682), .Y(n_734) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
INVx3_ASAP7_75t_L g561 ( .A(n_502), .Y(n_561) );
AND2x2_ASAP7_75t_L g609 ( .A(n_502), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g663 ( .A(n_502), .B(n_578), .Y(n_663) );
AND2x2_ASAP7_75t_L g721 ( .A(n_502), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g562 ( .A(n_511), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g578 ( .A(n_511), .Y(n_578) );
INVx1_ASAP7_75t_L g633 ( .A(n_511), .Y(n_633) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_511), .Y(n_639) );
AND2x2_ASAP7_75t_L g684 ( .A(n_511), .B(n_561), .Y(n_684) );
OR2x2_ASAP7_75t_L g723 ( .A(n_511), .B(n_563), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_516), .B(n_519), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_521), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_529), .Y(n_521) );
AND2x2_ASAP7_75t_L g719 ( .A(n_522), .B(n_716), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_522), .B(n_701), .Y(n_751) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g650 ( .A(n_523), .B(n_574), .Y(n_650) );
AND2x2_ASAP7_75t_L g699 ( .A(n_523), .B(n_547), .Y(n_699) );
INVx1_ASAP7_75t_L g745 ( .A(n_523), .Y(n_745) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_524), .Y(n_559) );
AND2x2_ASAP7_75t_L g600 ( .A(n_524), .B(n_574), .Y(n_600) );
INVx1_ASAP7_75t_L g617 ( .A(n_524), .Y(n_617) );
AND2x2_ASAP7_75t_L g623 ( .A(n_524), .B(n_540), .Y(n_623) );
AND2x2_ASAP7_75t_L g691 ( .A(n_529), .B(n_599), .Y(n_691) );
INVx2_ASAP7_75t_L g756 ( .A(n_529), .Y(n_756) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_540), .Y(n_529) );
AND2x2_ASAP7_75t_L g573 ( .A(n_530), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g586 ( .A(n_530), .B(n_548), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_530), .B(n_547), .Y(n_614) );
INVx1_ASAP7_75t_L g620 ( .A(n_530), .Y(n_620) );
INVx1_ASAP7_75t_L g637 ( .A(n_530), .Y(n_637) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_530), .Y(n_649) );
INVx2_ASAP7_75t_L g717 ( .A(n_530), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
INVx2_ASAP7_75t_L g574 ( .A(n_540), .Y(n_574) );
BUFx2_ASAP7_75t_L g671 ( .A(n_540), .Y(n_671) );
AND2x2_ASAP7_75t_L g716 ( .A(n_540), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_546), .B(n_653), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_546), .A2(n_715), .B(n_729), .Y(n_739) );
AND2x2_ASAP7_75t_L g764 ( .A(n_546), .B(n_650), .Y(n_764) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g686 ( .A(n_548), .Y(n_686) );
AND2x2_ASAP7_75t_L g715 ( .A(n_548), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_549), .Y(n_599) );
INVx2_ASAP7_75t_L g618 ( .A(n_549), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_549), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
OR2x2_ASAP7_75t_L g585 ( .A(n_559), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g653 ( .A(n_559), .B(n_649), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_559), .B(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g754 ( .A(n_559), .B(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_559), .B(n_691), .Y(n_766) );
AND2x2_ASAP7_75t_L g645 ( .A(n_560), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g668 ( .A(n_560), .B(n_562), .Y(n_668) );
INVx2_ASAP7_75t_L g580 ( .A(n_561), .Y(n_580) );
AND2x2_ASAP7_75t_L g608 ( .A(n_561), .B(n_581), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_561), .B(n_633), .Y(n_689) );
AND2x2_ASAP7_75t_L g603 ( .A(n_562), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g750 ( .A(n_562), .Y(n_750) );
AND2x2_ASAP7_75t_L g762 ( .A(n_562), .B(n_625), .Y(n_762) );
AND2x2_ASAP7_75t_L g588 ( .A(n_563), .B(n_578), .Y(n_588) );
INVx1_ASAP7_75t_L g683 ( .A(n_563), .Y(n_683) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g581 ( .A(n_568), .B(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_572), .B(n_619), .Y(n_628) );
OR2x2_ASAP7_75t_L g760 ( .A(n_572), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g677 ( .A(n_573), .B(n_618), .Y(n_677) );
AND2x2_ASAP7_75t_L g685 ( .A(n_573), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g744 ( .A(n_573), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g768 ( .A(n_573), .B(n_615), .Y(n_768) );
NOR2xp67_ASAP7_75t_L g726 ( .A(n_574), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g755 ( .A(n_574), .B(n_618), .Y(n_755) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
AND2x2_ASAP7_75t_L g607 ( .A(n_577), .B(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g769 ( .A(n_577), .Y(n_769) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g604 ( .A(n_580), .Y(n_604) );
AND2x2_ASAP7_75t_L g655 ( .A(n_580), .B(n_588), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_580), .B(n_723), .Y(n_749) );
INVx2_ASAP7_75t_L g594 ( .A(n_581), .Y(n_594) );
INVx3_ASAP7_75t_L g646 ( .A(n_581), .Y(n_646) );
OR2x2_ASAP7_75t_L g674 ( .A(n_581), .B(n_675), .Y(n_674) );
AOI311xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .A3(n_589), .B(n_590), .C(n_601), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_584), .A2(n_622), .B(n_624), .C(n_626), .Y(n_621) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_SL g606 ( .A(n_586), .Y(n_606) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g624 ( .A(n_588), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_588), .B(n_604), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_588), .B(n_589), .Y(n_757) );
AND2x2_ASAP7_75t_L g679 ( .A(n_589), .B(n_593), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_595), .B(n_596), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g737 ( .A(n_593), .B(n_625), .Y(n_737) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_594), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g631 ( .A(n_594), .Y(n_631) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_L g622 ( .A(n_598), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g667 ( .A(n_600), .Y(n_667) );
AND2x4_ASAP7_75t_L g729 ( .A(n_600), .B(n_698), .Y(n_729) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_603), .A2(n_669), .B1(n_681), .B2(n_685), .C1(n_687), .C2(n_691), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B(n_609), .C(n_612), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_606), .B(n_650), .Y(n_673) );
INVx1_ASAP7_75t_L g695 ( .A(n_608), .Y(n_695) );
INVx1_ASAP7_75t_L g629 ( .A(n_610), .Y(n_629) );
OR2x2_ASAP7_75t_L g694 ( .A(n_611), .B(n_695), .Y(n_694) );
OAI21xp33_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_615), .B(n_619), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_613), .B(n_631), .C(n_632), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_613), .A2(n_650), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_617), .Y(n_670) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_618), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g727 ( .A(n_618), .Y(n_727) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_618), .Y(n_743) );
INVx2_ASAP7_75t_L g701 ( .A(n_619), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_623), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g675 ( .A(n_625), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_630), .B2(n_634), .C(n_635), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_629), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g763 ( .A(n_629), .Y(n_763) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g644 ( .A(n_636), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_636), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g702 ( .A(n_636), .B(n_650), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_636), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g735 ( .A(n_636), .B(n_670), .Y(n_735) );
BUFx3_ASAP7_75t_L g698 ( .A(n_637), .Y(n_698) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND5xp2_ASAP7_75t_L g640 ( .A(n_641), .B(n_659), .C(n_680), .D(n_692), .E(n_707), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI32xp33_ASAP7_75t_L g732 ( .A1(n_644), .A2(n_671), .A3(n_687), .B1(n_733), .B2(n_735), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_646), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g656 ( .A(n_650), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_666), .B1(n_668), .B2(n_669), .C(n_672), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g731 ( .A(n_663), .B(n_682), .Y(n_731) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_668), .A2(n_729), .B1(n_747), .B2(n_752), .C(n_753), .Y(n_746) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_L g712 ( .A(n_671), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_676), .B2(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g690 ( .A(n_682), .Y(n_690) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_696), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_703), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_701), .A2(n_748), .B1(n_750), .B2(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_713), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_718), .B(n_720), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g761 ( .A(n_716), .Y(n_761) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B(n_730), .C(n_732), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI211xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B(n_740), .C(n_765), .Y(n_736) );
CKINVDCx16_ASAP7_75t_R g741 ( .A(n_737), .Y(n_741) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B(n_746), .C(n_758), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .B(n_757), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI21xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B(n_769), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
endmodule