module fake_jpeg_7092_n_39 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_39);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_7),
.B1(n_10),
.B2(n_14),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_17),
.B1(n_5),
.B2(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_19),
.A2(n_15),
.B1(n_8),
.B2(n_12),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_2),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_23),
.B1(n_35),
.B2(n_28),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_35),
.A3(n_23),
.B1(n_31),
.B2(n_22),
.C1(n_20),
.C2(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_27),
.Y(n_39)
);


endmodule