module fake_netlist_6_4231_n_1671 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1671);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1671;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_29),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_27),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_72),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_48),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_33),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_52),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_17),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_130),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_6),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_24),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_80),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_8),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_43),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_30),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_50),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_17),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_14),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_75),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_104),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_66),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_121),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_51),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_4),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_56),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_45),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_101),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_57),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_48),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_5),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_13),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_40),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_63),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_49),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_30),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_132),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_41),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_38),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_124),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_144),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_24),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_71),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_103),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_23),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_96),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_69),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_29),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_53),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_108),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_134),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_126),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_95),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_82),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_109),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_102),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_20),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_15),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_31),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_89),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_28),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_70),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_81),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_100),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_49),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_15),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_51),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_64),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_99),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_61),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_25),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_123),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_58),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_46),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_44),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_106),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_6),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_13),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_68),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_1),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_44),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_92),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_34),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_54),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_65),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_36),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_45),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_9),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_59),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_67),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_84),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_87),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_47),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_37),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_62),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_19),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_18),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_25),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_27),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_20),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_18),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_77),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_83),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_22),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_285),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_188),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_190),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_189),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_200),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_184),
.B(n_1),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_206),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_206),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_206),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_249),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_R g308 ( 
.A(n_205),
.B(n_210),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_222),
.B(n_3),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_214),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_206),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_217),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_218),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_221),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_224),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_191),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_226),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_227),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_229),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_231),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_259),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_259),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_259),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_254),
.B(n_7),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_237),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_194),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_240),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_194),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_243),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_245),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_246),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_247),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_209),
.B(n_8),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_253),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_255),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_259),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_238),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g343 ( 
.A(n_250),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_186),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_148),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_173),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_196),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_148),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_201),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_173),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_201),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_198),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_208),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_209),
.B(n_10),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_208),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_154),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_213),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_238),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_213),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_234),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_261),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_261),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_149),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_154),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_202),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_149),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_147),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_203),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_147),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_298),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_151),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_299),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_156),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_301),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_310),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_304),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_304),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_360),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_297),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_318),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_305),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_317),
.B(n_274),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_317),
.B(n_274),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_201),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_305),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_313),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_306),
.B(n_156),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_314),
.Y(n_396)
);

AND3x2_ASAP7_75t_L g397 ( 
.A(n_302),
.B(n_174),
.C(n_212),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_306),
.B(n_158),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_350),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_352),
.B(n_212),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_315),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_150),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_322),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_324),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_353),
.B(n_157),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_338),
.A2(n_160),
.B(n_146),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_325),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_346),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_311),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_312),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_330),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_357),
.B(n_273),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_312),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_323),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_316),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_335),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_233),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_333),
.B(n_155),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_319),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_332),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_321),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_321),
.B(n_161),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_334),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_309),
.B(n_201),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_337),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_326),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_327),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_320),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_327),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_328),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

CKINVDCx11_ASAP7_75t_R g442 ( 
.A(n_385),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_409),
.Y(n_443)
);

INVx4_ASAP7_75t_SL g444 ( 
.A(n_430),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_390),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_309),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_422),
.A2(n_355),
.B1(n_343),
.B2(n_155),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_201),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_383),
.B(n_408),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_339),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_383),
.B(n_303),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_418),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_303),
.Y(n_461)
);

NAND2x1p5_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_383),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_386),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_406),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_430),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_376),
.B(n_308),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_328),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_391),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_376),
.B(n_341),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_423),
.B(n_365),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_391),
.B(n_400),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_369),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_430),
.B(n_395),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_437),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_398),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_400),
.B(n_233),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_398),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_430),
.B(n_341),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_392),
.B(n_257),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_410),
.A2(n_271),
.B1(n_371),
.B2(n_197),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_412),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_373),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_424),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_397),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_400),
.B(n_257),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_424),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_379),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_379),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_410),
.B(n_368),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_387),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_411),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_400),
.B(n_344),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_392),
.B(n_257),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_381),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_410),
.B(n_368),
.Y(n_509)
);

INVx4_ASAP7_75t_SL g510 ( 
.A(n_392),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_380),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_377),
.B(n_336),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_387),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_378),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_372),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_400),
.B(n_257),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_381),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_428),
.B(n_257),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_394),
.B(n_340),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_387),
.Y(n_522)
);

BUFx8_ASAP7_75t_SL g523 ( 
.A(n_416),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_412),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_392),
.Y(n_526)
);

NOR2x1p5_ASAP7_75t_L g527 ( 
.A(n_396),
.B(n_271),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_428),
.B(n_165),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_401),
.B(n_349),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_410),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_382),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_405),
.A2(n_366),
.B1(n_358),
.B2(n_307),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_402),
.B(n_347),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_419),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_389),
.B(n_347),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_392),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_426),
.B(n_161),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_429),
.B(n_265),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_434),
.A2(n_171),
.B1(n_179),
.B2(n_295),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_421),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_372),
.B(n_275),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_393),
.B(n_168),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_393),
.B(n_170),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_432),
.B(n_265),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_397),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_399),
.B(n_265),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_403),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_433),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_440),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_387),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_413),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_433),
.B(n_162),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_413),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_415),
.Y(n_559)
);

BUFx4f_ASAP7_75t_L g560 ( 
.A(n_392),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_392),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_440),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_402),
.B(n_164),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_420),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_435),
.B(n_351),
.Y(n_567)
);

OR2x2_ASAP7_75t_SL g568 ( 
.A(n_435),
.B(n_185),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_388),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_427),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_427),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_440),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_407),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_436),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_455),
.B(n_436),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_441),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_449),
.A2(n_260),
.B1(n_187),
.B2(n_219),
.Y(n_578)
);

AND2x2_ASAP7_75t_SL g579 ( 
.A(n_454),
.B(n_265),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_477),
.B(n_162),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_449),
.A2(n_166),
.B1(n_295),
.B2(n_293),
.Y(n_581)
);

BUFx5_ASAP7_75t_L g582 ( 
.A(n_530),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_456),
.B(n_436),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_469),
.B(n_466),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_450),
.B(n_166),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_458),
.B(n_167),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_449),
.A2(n_239),
.B1(n_235),
.B2(n_242),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_458),
.B(n_167),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_462),
.B(n_265),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_461),
.B(n_169),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_460),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_460),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_471),
.B(n_351),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_470),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_470),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_475),
.B(n_169),
.Y(n_596)
);

BUFx6f_ASAP7_75t_SL g597 ( 
.A(n_504),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_449),
.B(n_404),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_446),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_462),
.A2(n_192),
.B1(n_195),
.B2(n_193),
.Y(n_600)
);

NOR2xp67_ASAP7_75t_L g601 ( 
.A(n_537),
.B(n_171),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_449),
.B(n_574),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_449),
.A2(n_176),
.B1(n_293),
.B2(n_177),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_447),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_459),
.B(n_207),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_559),
.B(n_404),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_481),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_481),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_492),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_559),
.B(n_407),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_482),
.B(n_443),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_473),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_471),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_448),
.Y(n_615)
);

AND2x6_ASAP7_75t_SL g616 ( 
.A(n_529),
.B(n_248),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_453),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_528),
.B(n_407),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_542),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_452),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_473),
.B(n_354),
.Y(n_621)
);

INVxp33_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_552),
.B(n_288),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_473),
.B(n_414),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_459),
.B(n_207),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_501),
.B(n_414),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_493),
.B(n_354),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_501),
.B(n_414),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_493),
.B(n_356),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_509),
.B(n_180),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_445),
.B(n_177),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_445),
.B(n_178),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_509),
.B(n_183),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_495),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_457),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_547),
.B(n_557),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_511),
.B(n_152),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_547),
.B(n_178),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_468),
.B(n_228),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_549),
.A2(n_181),
.B1(n_179),
.B2(n_182),
.Y(n_640)
);

AND2x2_ASAP7_75t_SL g641 ( 
.A(n_454),
.B(n_230),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_472),
.B(n_467),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_526),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_495),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_544),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_467),
.B(n_232),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_497),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_467),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_539),
.B(n_181),
.Y(n_649)
);

INVxp33_ASAP7_75t_L g650 ( 
.A(n_464),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_497),
.Y(n_651)
);

AO22x1_ASAP7_75t_L g652 ( 
.A1(n_530),
.A2(n_175),
.B1(n_296),
.B2(n_294),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_499),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_544),
.B(n_288),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_479),
.A2(n_244),
.B(n_258),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_499),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_527),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_489),
.A2(n_519),
.B1(n_451),
.B2(n_485),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_483),
.A2(n_182),
.B1(n_268),
.B2(n_262),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_506),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_539),
.B(n_262),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_506),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_535),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_535),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_540),
.B(n_268),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_519),
.A2(n_289),
.B1(n_277),
.B2(n_287),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_563),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_508),
.B(n_282),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_518),
.B(n_225),
.C(n_236),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_459),
.B(n_207),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_505),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_490),
.B(n_288),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_567),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_563),
.A2(n_276),
.B1(n_204),
.B2(n_263),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_531),
.B(n_207),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_543),
.B(n_207),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_567),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_569),
.A2(n_364),
.B(n_363),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_465),
.B(n_207),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_551),
.B(n_211),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_553),
.B(n_207),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_556),
.B(n_564),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_568),
.A2(n_215),
.B1(n_216),
.B2(n_220),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_505),
.Y(n_686)
);

BUFx6f_ASAP7_75t_SL g687 ( 
.A(n_504),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_565),
.B(n_207),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_465),
.B(n_223),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_558),
.B(n_241),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_566),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_571),
.B(n_251),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_525),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_563),
.A2(n_484),
.B1(n_558),
.B2(n_465),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_484),
.A2(n_267),
.B1(n_290),
.B2(n_256),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_558),
.B(n_152),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_572),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_496),
.B(n_153),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_491),
.B(n_153),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_575),
.B(n_159),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_569),
.A2(n_364),
.B(n_363),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_512),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_502),
.B(n_361),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_545),
.B(n_159),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_533),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_504),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_521),
.B(n_361),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_491),
.B(n_515),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_533),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_502),
.B(n_359),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_496),
.B(n_296),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_515),
.B(n_294),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_546),
.B(n_292),
.C(n_291),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_513),
.B(n_291),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_533),
.A2(n_286),
.B1(n_284),
.B2(n_283),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_569),
.A2(n_286),
.B1(n_284),
.B2(n_283),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_520),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_526),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_513),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_570),
.B(n_278),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_444),
.B(n_79),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_570),
.B(n_278),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_534),
.B(n_272),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_496),
.B(n_272),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_522),
.B(n_555),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_463),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_541),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_658),
.A2(n_560),
.B1(n_486),
.B2(n_526),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_708),
.B(n_693),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_626),
.A2(n_560),
.B(n_514),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_614),
.B(n_444),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_584),
.B(n_570),
.Y(n_733)
);

CKINVDCx6p67_ASAP7_75t_R g734 ( 
.A(n_597),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_628),
.A2(n_536),
.B(n_514),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_602),
.A2(n_536),
.B(n_561),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_598),
.A2(n_536),
.B(n_561),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_636),
.B(n_532),
.Y(n_738)
);

AOI21x1_ASAP7_75t_L g739 ( 
.A1(n_605),
.A2(n_494),
.B(n_517),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_619),
.B(n_444),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_624),
.A2(n_500),
.B(n_498),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_580),
.B(n_478),
.Y(n_742)
);

OAI21xp5_ASAP7_75t_L g743 ( 
.A1(n_630),
.A2(n_488),
.B(n_480),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_637),
.B(n_494),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_643),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_699),
.A2(n_487),
.B(n_507),
.C(n_554),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_621),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_633),
.A2(n_488),
.B(n_480),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_699),
.A2(n_487),
.B(n_507),
.C(n_554),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_580),
.B(n_522),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_606),
.A2(n_500),
.B(n_474),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_703),
.B(n_522),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_613),
.A2(n_555),
.B1(n_522),
.B2(n_488),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_621),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_613),
.A2(n_555),
.B1(n_480),
.B2(n_478),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_583),
.B(n_478),
.Y(n_756)
);

AOI21x1_ASAP7_75t_L g757 ( 
.A1(n_605),
.A2(n_573),
.B(n_562),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_658),
.A2(n_573),
.B(n_562),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_620),
.B(n_442),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_684),
.B(n_555),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_684),
.B(n_538),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_674),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_667),
.B(n_163),
.C(n_172),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_611),
.B(n_163),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_599),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_618),
.A2(n_476),
.B(n_498),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_663),
.Y(n_767)
);

OAI21xp33_ASAP7_75t_L g768 ( 
.A1(n_596),
.A2(n_172),
.B(n_175),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_610),
.A2(n_500),
.B(n_476),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_707),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_623),
.B(n_463),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_576),
.A2(n_548),
.B(n_550),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_705),
.B(n_510),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_625),
.A2(n_550),
.B(n_270),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_611),
.B(n_631),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_705),
.B(n_510),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_586),
.A2(n_264),
.B(n_269),
.C(n_270),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_586),
.A2(n_264),
.B(n_269),
.C(n_503),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_665),
.B(n_510),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_666),
.B(n_550),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_601),
.B(n_503),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_631),
.B(n_442),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_582),
.B(n_464),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_632),
.B(n_10),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_660),
.A2(n_550),
.B1(n_113),
.B2(n_141),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_712),
.A2(n_725),
.B(n_679),
.C(n_675),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_643),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_625),
.A2(n_138),
.B(n_137),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_578),
.B(n_587),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_604),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_642),
.A2(n_133),
.B(n_120),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_672),
.A2(n_118),
.B(n_116),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_726),
.A2(n_114),
.B(n_107),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_587),
.B(n_11),
.Y(n_795)
);

OAI21xp33_ASAP7_75t_L g796 ( 
.A1(n_596),
.A2(n_523),
.B(n_16),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_681),
.A2(n_105),
.B(n_97),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_694),
.A2(n_93),
.B1(n_86),
.B2(n_74),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_691),
.B(n_12),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_689),
.A2(n_19),
.B(n_21),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_689),
.A2(n_21),
.B(n_22),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_577),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_643),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_645),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_615),
.B(n_26),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_660),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_617),
.B(n_28),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_635),
.B(n_31),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_667),
.B(n_523),
.C(n_33),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_597),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_664),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_577),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_654),
.B(n_32),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_638),
.B(n_32),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_709),
.B(n_34),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_638),
.B(n_649),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_712),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_662),
.A2(n_39),
.B(n_40),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_643),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_632),
.B(n_39),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_662),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_648),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_649),
.B(n_42),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_661),
.B(n_706),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_SL g825 ( 
.A1(n_600),
.A2(n_688),
.B(n_678),
.C(n_677),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_701),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_655),
.A2(n_607),
.B(n_647),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_661),
.B(n_710),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_588),
.B(n_627),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_700),
.B(n_713),
.C(n_724),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_585),
.B(n_588),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_704),
.A2(n_711),
.B(n_639),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_646),
.A2(n_719),
.B(n_721),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_622),
.B(n_585),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_627),
.B(n_629),
.Y(n_835)
);

AO21x1_ASAP7_75t_L g836 ( 
.A1(n_581),
.A2(n_603),
.B(n_683),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_582),
.B(n_723),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_629),
.B(n_593),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_719),
.A2(n_720),
.B(n_595),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_590),
.B(n_696),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_594),
.A2(n_697),
.B(n_715),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_692),
.A2(n_722),
.B(n_644),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_722),
.Y(n_843)
);

OR2x6_ASAP7_75t_SL g844 ( 
.A(n_717),
.B(n_714),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_593),
.B(n_582),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_591),
.A2(n_651),
.B(n_718),
.Y(n_846)
);

OR2x4_ASAP7_75t_L g847 ( 
.A(n_682),
.B(n_701),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_582),
.B(n_682),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_582),
.B(n_695),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_591),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_582),
.B(n_695),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_592),
.A2(n_644),
.B(n_608),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_670),
.B(n_647),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_609),
.A2(n_686),
.B(n_612),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_612),
.A2(n_656),
.B(n_718),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_634),
.A2(n_673),
.B(n_656),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_651),
.A2(n_653),
.B(n_702),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_653),
.B(n_652),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_690),
.A2(n_685),
.B(n_668),
.C(n_657),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_641),
.A2(n_680),
.B(n_579),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_641),
.A2(n_579),
.B(n_671),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_659),
.B(n_669),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_668),
.B(n_716),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_640),
.B(n_676),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_698),
.B(n_728),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_616),
.A2(n_650),
.B(n_687),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_727),
.A2(n_658),
.B1(n_636),
.B2(n_578),
.Y(n_867)
);

AND2x6_ASAP7_75t_SL g868 ( 
.A(n_687),
.B(n_529),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_621),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_584),
.B(n_455),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_626),
.A2(n_569),
.B(n_628),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_643),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_636),
.B(n_584),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_626),
.A2(n_569),
.B(n_628),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_584),
.B(n_455),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_584),
.B(n_455),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_584),
.B(n_455),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_626),
.A2(n_569),
.B(n_628),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_584),
.B(n_455),
.Y(n_879)
);

NAND3xp33_ASAP7_75t_L g880 ( 
.A(n_580),
.B(n_636),
.C(n_667),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_658),
.A2(n_636),
.B1(n_578),
.B2(n_587),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_584),
.B(n_455),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_584),
.B(n_455),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_584),
.B(n_455),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_655),
.A2(n_576),
.B(n_589),
.C(n_584),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_597),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_589),
.A2(n_462),
.B(n_626),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_584),
.B(n_455),
.Y(n_888)
);

AO32x1_ASAP7_75t_L g889 ( 
.A1(n_600),
.A2(n_697),
.A3(n_599),
.B1(n_617),
.B2(n_615),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_584),
.B(n_455),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_584),
.A2(n_455),
.B(n_636),
.C(n_422),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_693),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_621),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_708),
.B(n_693),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_584),
.A2(n_455),
.B(n_636),
.C(n_422),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_626),
.A2(n_569),
.B(n_628),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_643),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_880),
.A2(n_816),
.B1(n_877),
.B2(n_882),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_848),
.A2(n_874),
.B(n_871),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_878),
.A2(n_896),
.B(n_733),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_SL g901 ( 
.A(n_886),
.B(n_810),
.Y(n_901)
);

BUFx10_ASAP7_75t_L g902 ( 
.A(n_868),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_802),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_831),
.B(n_775),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_767),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_812),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_887),
.A2(n_876),
.B(n_870),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_745),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_875),
.B(n_877),
.Y(n_909)
);

AO21x1_ASAP7_75t_L g910 ( 
.A1(n_881),
.A2(n_820),
.B(n_785),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_775),
.B(n_738),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_879),
.B(n_883),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_884),
.B(n_888),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_765),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_885),
.A2(n_882),
.B(n_875),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_788),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_791),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_890),
.B(n_873),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_843),
.B(n_788),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_891),
.B(n_895),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_SL g921 ( 
.A1(n_864),
.A2(n_809),
.B(n_764),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_885),
.A2(n_842),
.B(n_748),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_730),
.B(n_894),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_785),
.A2(n_820),
.B(n_790),
.C(n_787),
.Y(n_924)
);

AOI21x1_ASAP7_75t_SL g925 ( 
.A1(n_823),
.A2(n_814),
.B(n_858),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_743),
.A2(n_760),
.B(n_825),
.Y(n_926)
);

BUFx2_ASAP7_75t_SL g927 ( 
.A(n_767),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_829),
.A2(n_859),
.B(n_840),
.C(n_862),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_867),
.B(n_826),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_834),
.B(n_764),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_834),
.B(n_762),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_826),
.B(n_761),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_830),
.A2(n_840),
.B1(n_762),
.B2(n_843),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_846),
.A2(n_856),
.B(n_741),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_745),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_849),
.A2(n_851),
.B(n_729),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_759),
.B(n_770),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_860),
.A2(n_861),
.B(n_758),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_759),
.B(n_804),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_800),
.A2(n_863),
.B1(n_795),
.B2(n_763),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_847),
.B(n_892),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_833),
.A2(n_731),
.B(n_750),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_824),
.B(n_828),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_766),
.A2(n_751),
.B(n_852),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_750),
.B(n_845),
.Y(n_945)
);

NAND3x1_ASAP7_75t_L g946 ( 
.A(n_783),
.B(n_830),
.C(n_821),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_747),
.B(n_754),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_771),
.Y(n_948)
);

OAI21xp33_ASAP7_75t_L g949 ( 
.A1(n_768),
.A2(n_815),
.B(n_796),
.Y(n_949)
);

OAI21x1_ASAP7_75t_SL g950 ( 
.A1(n_789),
.A2(n_797),
.B(n_793),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_854),
.A2(n_855),
.B(n_769),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_739),
.A2(n_841),
.B(n_832),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_745),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_892),
.B(n_813),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_778),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_742),
.A2(n_756),
.B(n_772),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_837),
.A2(n_746),
.B(n_749),
.Y(n_957)
);

AOI221x1_ASAP7_75t_L g958 ( 
.A1(n_801),
.A2(n_779),
.B1(n_798),
.B2(n_777),
.C(n_818),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_839),
.A2(n_736),
.B(n_737),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_752),
.B(n_853),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_752),
.B(n_806),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_806),
.B(n_835),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_732),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_735),
.A2(n_773),
.B(n_776),
.Y(n_964)
);

NAND2x1_ASAP7_75t_L g965 ( 
.A(n_745),
.B(n_872),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_838),
.B(n_744),
.Y(n_966)
);

AOI21xp33_ASAP7_75t_L g967 ( 
.A1(n_865),
.A2(n_893),
.B(n_869),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_778),
.B(n_783),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_811),
.Y(n_969)
);

OAI21xp33_ASAP7_75t_L g970 ( 
.A1(n_799),
.A2(n_807),
.B(n_805),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_847),
.B(n_822),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_759),
.B(n_784),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_803),
.A2(n_897),
.B(n_819),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_850),
.B(n_872),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_781),
.A2(n_780),
.B(n_774),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_734),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_836),
.A2(n_889),
.B(n_808),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_755),
.A2(n_753),
.B(n_732),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_782),
.B(n_844),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_872),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_850),
.B(n_872),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_792),
.B(n_740),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_850),
.A2(n_786),
.B1(n_817),
.B2(n_794),
.Y(n_983)
);

AO21x2_ASAP7_75t_L g984 ( 
.A1(n_889),
.A2(n_850),
.B(n_866),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_767),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_848),
.A2(n_896),
.B(n_874),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_775),
.B(n_703),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_848),
.A2(n_896),
.B(n_874),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_757),
.A2(n_857),
.B(n_827),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_880),
.A2(n_877),
.B(n_882),
.C(n_875),
.Y(n_990)
);

OA22x2_ASAP7_75t_L g991 ( 
.A1(n_796),
.A2(n_676),
.B1(n_738),
.B2(n_864),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_730),
.B(n_727),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_767),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_875),
.B(n_877),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_757),
.A2(n_857),
.B(n_827),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_843),
.B(n_788),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_880),
.A2(n_885),
.B(n_816),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_757),
.A2(n_857),
.B(n_827),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_757),
.A2(n_857),
.B(n_827),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_730),
.B(n_894),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_875),
.B(n_877),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_875),
.B(n_877),
.Y(n_1002)
);

CKINVDCx6p67_ASAP7_75t_R g1003 ( 
.A(n_759),
.Y(n_1003)
);

AOI21xp33_ASAP7_75t_L g1004 ( 
.A1(n_880),
.A2(n_775),
.B(n_816),
.Y(n_1004)
);

AO31x2_ASAP7_75t_L g1005 ( 
.A1(n_881),
.A2(n_836),
.A3(n_600),
.B(n_860),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_767),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_875),
.B(n_877),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_802),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_875),
.B(n_877),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_802),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_875),
.B(n_877),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_816),
.A2(n_880),
.B(n_823),
.C(n_636),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_875),
.B(n_877),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_880),
.A2(n_816),
.B1(n_877),
.B2(n_875),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_880),
.A2(n_877),
.B(n_882),
.C(n_875),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_730),
.B(n_894),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_875),
.B(n_877),
.Y(n_1017)
);

INVxp67_ASAP7_75t_SL g1018 ( 
.A(n_845),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_730),
.B(n_727),
.Y(n_1019)
);

NOR2xp67_ASAP7_75t_L g1020 ( 
.A(n_762),
.B(n_693),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_767),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_880),
.A2(n_885),
.B(n_816),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_745),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_880),
.A2(n_877),
.B1(n_882),
.B2(n_875),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_875),
.B(n_877),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_L g1026 ( 
.A(n_880),
.B(n_544),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_880),
.A2(n_816),
.B1(n_877),
.B2(n_875),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_765),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_930),
.B(n_1000),
.Y(n_1029)
);

INVx3_ASAP7_75t_SL g1030 ( 
.A(n_976),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_921),
.A2(n_990),
.B(n_1015),
.C(n_1004),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1016),
.B(n_931),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_908),
.B(n_916),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_911),
.A2(n_1024),
.B(n_1017),
.C(n_1013),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_991),
.A2(n_910),
.B1(n_949),
.B2(n_987),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_905),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_985),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_947),
.B(n_955),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_909),
.A2(n_1002),
.B(n_1017),
.C(n_1007),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_909),
.A2(n_1011),
.B1(n_1002),
.B2(n_1001),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_923),
.B(n_954),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_991),
.A2(n_898),
.B1(n_1027),
.B2(n_1014),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_935),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_979),
.A2(n_940),
.B1(n_904),
.B2(n_941),
.Y(n_1044)
);

NAND2x1p5_ASAP7_75t_L g1045 ( 
.A(n_908),
.B(n_916),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_948),
.A2(n_1007),
.B1(n_1009),
.B2(n_1025),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_1006),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_935),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_968),
.B(n_992),
.Y(n_1049)
);

CKINVDCx8_ASAP7_75t_R g1050 ( 
.A(n_927),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_993),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_963),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_947),
.B(n_963),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_935),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_994),
.B(n_1001),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1019),
.B(n_1026),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_1020),
.B(n_994),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1009),
.B(n_1011),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1013),
.B(n_1025),
.Y(n_1059)
);

OAI321xp33_ASAP7_75t_L g1060 ( 
.A1(n_924),
.A2(n_915),
.A3(n_920),
.B1(n_929),
.B2(n_928),
.C(n_1022),
.Y(n_1060)
);

CKINVDCx6p67_ASAP7_75t_R g1061 ( 
.A(n_937),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_918),
.B(n_929),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_917),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_939),
.Y(n_1064)
);

BUFx4_ASAP7_75t_SL g1065 ( 
.A(n_937),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1012),
.A2(n_913),
.B1(n_912),
.B2(n_920),
.C(n_971),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_918),
.B(n_932),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_932),
.B(n_971),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1028),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_933),
.B(n_969),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_953),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_943),
.B(n_960),
.Y(n_1072)
);

CKINVDCx6p67_ASAP7_75t_R g1073 ( 
.A(n_937),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_943),
.B(n_960),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_1021),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_903),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_966),
.B(n_962),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_906),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_939),
.B(n_972),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_907),
.A2(n_922),
.B(n_900),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_953),
.Y(n_1081)
);

BUFx2_ASAP7_75t_R g1082 ( 
.A(n_984),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1008),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_939),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_962),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_967),
.B(n_972),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_945),
.B(n_961),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_972),
.B(n_1010),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_1023),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_1023),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_946),
.A2(n_945),
.B1(n_961),
.B2(n_978),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_974),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_997),
.B(n_1018),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_900),
.A2(n_942),
.B(n_926),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_901),
.B(n_970),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_936),
.B(n_974),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_908),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_981),
.B(n_956),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_981),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_902),
.Y(n_1100)
);

BUFx12f_ASAP7_75t_SL g1101 ( 
.A(n_1003),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_902),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_980),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1005),
.B(n_938),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_942),
.A2(n_926),
.B(n_988),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_980),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_984),
.B(n_996),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_965),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1005),
.B(n_958),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_950),
.A2(n_983),
.B1(n_957),
.B2(n_975),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_919),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_982),
.A2(n_996),
.B1(n_919),
.B2(n_977),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_973),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_952),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_899),
.A2(n_988),
.B(n_986),
.C(n_964),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1005),
.B(n_899),
.Y(n_1116)
);

INVx3_ASAP7_75t_SL g1117 ( 
.A(n_925),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_986),
.A2(n_964),
.B(n_959),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_934),
.A2(n_944),
.B1(n_951),
.B2(n_989),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_995),
.A2(n_738),
.B(n_921),
.C(n_775),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_998),
.B(n_999),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_947),
.B(n_778),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_909),
.A2(n_1001),
.B1(n_1002),
.B2(n_994),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_905),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_993),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_905),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_905),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_930),
.B(n_1000),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_909),
.B(n_994),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_909),
.A2(n_1001),
.B1(n_1002),
.B2(n_994),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_923),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_905),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_908),
.B(n_843),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_914),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_909),
.B(n_994),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_930),
.B(n_1000),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_993),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_914),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_911),
.A2(n_880),
.B1(n_991),
.B2(n_738),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_905),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_911),
.B(n_552),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_935),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_909),
.B(n_994),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_909),
.B(n_994),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_935),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_909),
.B(n_994),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_927),
.B(n_843),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_909),
.B(n_994),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_914),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_SL g1150 ( 
.A1(n_928),
.A2(n_881),
.B(n_990),
.Y(n_1150)
);

AND2x6_ASAP7_75t_L g1151 ( 
.A(n_963),
.B(n_916),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_947),
.B(n_778),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_935),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_911),
.A2(n_880),
.B(n_1024),
.C(n_775),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_935),
.Y(n_1155)
);

AO32x2_ASAP7_75t_L g1156 ( 
.A1(n_898),
.A2(n_1027),
.A3(n_1014),
.B1(n_881),
.B2(n_867),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_911),
.B(n_552),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_930),
.B(n_1000),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_909),
.B(n_994),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_990),
.A2(n_1015),
.B(n_924),
.C(n_928),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_909),
.B(n_994),
.Y(n_1161)
);

OR2x2_ASAP7_75t_SL g1162 ( 
.A(n_923),
.B(n_809),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_911),
.B(n_552),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_930),
.B(n_1000),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_914),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_909),
.A2(n_1001),
.B1(n_1002),
.B2(n_994),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1047),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1063),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1070),
.Y(n_1169)
);

CKINVDCx11_ASAP7_75t_R g1170 ( 
.A(n_1030),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1069),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1165),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1044),
.A2(n_1046),
.B1(n_1139),
.B2(n_1074),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1134),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_1125),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1138),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1149),
.Y(n_1177)
);

CKINVDCx11_ASAP7_75t_R g1178 ( 
.A(n_1100),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1076),
.Y(n_1179)
);

CKINVDCx9p33_ASAP7_75t_R g1180 ( 
.A(n_1037),
.Y(n_1180)
);

AO21x1_ASAP7_75t_SL g1181 ( 
.A1(n_1042),
.A2(n_1110),
.B(n_1109),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1070),
.B(n_1112),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1086),
.A2(n_1091),
.B1(n_1056),
.B2(n_1088),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1095),
.A2(n_1035),
.B1(n_1157),
.B2(n_1163),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1118),
.A2(n_1094),
.B(n_1080),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1043),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_1096),
.B(n_1104),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1053),
.B(n_1052),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_1047),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1078),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1051),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1083),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1092),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1151),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1085),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1068),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1077),
.Y(n_1197)
);

INVx6_ASAP7_75t_L g1198 ( 
.A(n_1043),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1154),
.B(n_1034),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_1097),
.B(n_1043),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1131),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1067),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1062),
.B(n_1072),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1141),
.A2(n_1144),
.B1(n_1161),
.B2(n_1159),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1092),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1029),
.B(n_1128),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1081),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1121),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1136),
.B(n_1158),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1091),
.A2(n_1164),
.B1(n_1057),
.B2(n_1079),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1099),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1099),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1032),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1031),
.A2(n_1120),
.B(n_1150),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1151),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1055),
.B(n_1058),
.Y(n_1216)
);

AO21x1_ASAP7_75t_L g1217 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1116),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1055),
.B(n_1058),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1079),
.A2(n_1049),
.B1(n_1131),
.B2(n_1166),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1084),
.A2(n_1064),
.B1(n_1135),
.B2(n_1143),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1041),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1098),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1098),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1079),
.A2(n_1166),
.B1(n_1130),
.B2(n_1123),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1096),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1093),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1108),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1072),
.B(n_1074),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1104),
.B(n_1087),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1103),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1065),
.Y(n_1231)
);

CKINVDCx11_ASAP7_75t_R g1232 ( 
.A(n_1102),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1081),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1127),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1116),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1059),
.B(n_1129),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1081),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1156),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1087),
.A2(n_1113),
.B(n_1123),
.Y(n_1239)
);

AND2x6_ASAP7_75t_L g1240 ( 
.A(n_1107),
.B(n_1135),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1040),
.A2(n_1130),
.B1(n_1129),
.B2(n_1146),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1089),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1097),
.B(n_1155),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1059),
.A2(n_1148),
.B1(n_1143),
.B2(n_1146),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1132),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1145),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1052),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1039),
.B(n_1159),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1122),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1075),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1060),
.A2(n_1119),
.B(n_1114),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1122),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1152),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1050),
.Y(n_1254)
);

INVx8_ASAP7_75t_L g1255 ( 
.A(n_1145),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1152),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1151),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1145),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1115),
.A2(n_1066),
.B(n_1040),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1048),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1144),
.B(n_1148),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1117),
.A2(n_1161),
.B1(n_1053),
.B2(n_1038),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1033),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1082),
.B(n_1038),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1048),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1101),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1155),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1061),
.A2(n_1073),
.B1(n_1036),
.B2(n_1124),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1162),
.A2(n_1137),
.B1(n_1147),
.B2(n_1140),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1126),
.A2(n_1147),
.B1(n_1111),
.B2(n_1106),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1054),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1147),
.A2(n_1133),
.B1(n_1045),
.B2(n_1033),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1155),
.Y(n_1273)
);

AO21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1160),
.A2(n_1133),
.B(n_1045),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1071),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1090),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1142),
.B(n_1153),
.Y(n_1277)
);

BUFx2_ASAP7_75t_R g1278 ( 
.A(n_1030),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1063),
.Y(n_1279)
);

INVx11_ASAP7_75t_L g1280 ( 
.A(n_1100),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1118),
.A2(n_1094),
.B(n_1105),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1047),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1063),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1199),
.A2(n_1214),
.B1(n_1173),
.B2(n_1183),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1235),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1281),
.A2(n_1259),
.B(n_1217),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1238),
.B(n_1261),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1193),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1178),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1255),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1169),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1206),
.B(n_1209),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1238),
.B(n_1261),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1217),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1170),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1228),
.B(n_1187),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1193),
.Y(n_1297)
);

INVx8_ASAP7_75t_L g1298 ( 
.A(n_1255),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1205),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1228),
.B(n_1203),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1255),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1205),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1199),
.A2(n_1184),
.B1(n_1210),
.B2(n_1169),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1239),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1187),
.B(n_1229),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1229),
.B(n_1203),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1212),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1189),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1207),
.A2(n_1258),
.B(n_1267),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1224),
.B(n_1226),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1216),
.B(n_1218),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1212),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1250),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1208),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1182),
.B(n_1248),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1201),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1185),
.A2(n_1204),
.B(n_1244),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1248),
.B(n_1181),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1182),
.B(n_1272),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1219),
.A2(n_1269),
.B1(n_1262),
.B2(n_1241),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1181),
.B(n_1240),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1251),
.A2(n_1182),
.B(n_1215),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1274),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1197),
.B(n_1195),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1240),
.B(n_1177),
.Y(n_1325)
);

INVx8_ASAP7_75t_L g1326 ( 
.A(n_1277),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1236),
.B(n_1196),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1202),
.B(n_1221),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1251),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1240),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1240),
.B(n_1222),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1174),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1167),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1223),
.B(n_1225),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1220),
.A2(n_1270),
.B1(n_1213),
.B2(n_1268),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1211),
.B(n_1282),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1176),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1249),
.A2(n_1252),
.B1(n_1253),
.B2(n_1256),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1194),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1168),
.B(n_1283),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1207),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1227),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1247),
.A2(n_1263),
.B(n_1171),
.Y(n_1343)
);

XOR2xp5_ASAP7_75t_L g1344 ( 
.A(n_1231),
.B(n_1278),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1175),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1245),
.B(n_1191),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1172),
.B(n_1279),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1215),
.B(n_1257),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1264),
.B(n_1190),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1179),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1192),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1264),
.B(n_1188),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1188),
.B(n_1230),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1200),
.A2(n_1243),
.B(n_1242),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1275),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1188),
.A2(n_1170),
.B1(n_1254),
.B2(n_1234),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1200),
.A2(n_1243),
.B(n_1271),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1287),
.B(n_1274),
.Y(n_1358)
);

INVx4_ASAP7_75t_L g1359 ( 
.A(n_1326),
.Y(n_1359)
);

AOI322xp5_ASAP7_75t_L g1360 ( 
.A1(n_1284),
.A2(n_1231),
.A3(n_1254),
.B1(n_1266),
.B2(n_1246),
.C1(n_1186),
.C2(n_1180),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1287),
.B(n_1260),
.Y(n_1361)
);

AOI21xp33_ASAP7_75t_L g1362 ( 
.A1(n_1317),
.A2(n_1246),
.B(n_1186),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1320),
.A2(n_1303),
.B1(n_1335),
.B2(n_1349),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1320),
.A2(n_1198),
.B1(n_1258),
.B2(n_1207),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1343),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1318),
.B(n_1267),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1330),
.Y(n_1367)
);

AND2x4_ASAP7_75t_SL g1368 ( 
.A(n_1319),
.B(n_1267),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1322),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1315),
.B(n_1265),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1293),
.B(n_1277),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1304),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1318),
.A2(n_1198),
.B1(n_1273),
.B2(n_1207),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1305),
.B(n_1258),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_1232),
.B2(n_1234),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1294),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1291),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1305),
.B(n_1258),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1329),
.B(n_1258),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1325),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1325),
.B(n_1331),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1331),
.B(n_1237),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1296),
.B(n_1237),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1289),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1317),
.A2(n_1233),
.B(n_1237),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1306),
.B(n_1267),
.Y(n_1386)
);

AOI221xp5_ASAP7_75t_L g1387 ( 
.A1(n_1292),
.A2(n_1266),
.B1(n_1267),
.B2(n_1273),
.C(n_1232),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1306),
.B(n_1285),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1388),
.B(n_1288),
.Y(n_1389)
);

OAI221xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1363),
.A2(n_1356),
.B1(n_1315),
.B2(n_1319),
.C(n_1310),
.Y(n_1390)
);

NAND3xp33_ASAP7_75t_L g1391 ( 
.A(n_1363),
.B(n_1338),
.C(n_1311),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1388),
.B(n_1302),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1370),
.B(n_1307),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1370),
.B(n_1316),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1374),
.B(n_1312),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1381),
.B(n_1321),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1374),
.B(n_1312),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1378),
.B(n_1300),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1381),
.B(n_1321),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1381),
.B(n_1319),
.Y(n_1400)
);

NAND3xp33_ASAP7_75t_L g1401 ( 
.A(n_1360),
.B(n_1333),
.C(n_1345),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1387),
.A2(n_1354),
.B1(n_1353),
.B2(n_1346),
.C(n_1313),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1360),
.B(n_1310),
.C(n_1327),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1378),
.B(n_1297),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1387),
.A2(n_1319),
.B1(n_1308),
.B2(n_1328),
.C(n_1336),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1364),
.A2(n_1352),
.B1(n_1289),
.B2(n_1348),
.Y(n_1406)
);

AOI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1362),
.A2(n_1355),
.B1(n_1332),
.B2(n_1337),
.C(n_1317),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1375),
.A2(n_1336),
.B1(n_1344),
.B2(n_1348),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1380),
.B(n_1322),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1375),
.A2(n_1344),
.B1(n_1348),
.B2(n_1295),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1364),
.A2(n_1352),
.B1(n_1348),
.B2(n_1291),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1359),
.B(n_1290),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1361),
.B(n_1299),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1361),
.B(n_1299),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1361),
.B(n_1299),
.Y(n_1415)
);

AND2x2_ASAP7_75t_SL g1416 ( 
.A(n_1368),
.B(n_1359),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1384),
.B(n_1324),
.Y(n_1417)
);

OAI21xp33_ASAP7_75t_L g1418 ( 
.A1(n_1373),
.A2(n_1324),
.B(n_1334),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1362),
.B(n_1350),
.C(n_1347),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1359),
.B(n_1290),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_L g1421 ( 
.A(n_1385),
.B(n_1314),
.C(n_1342),
.Y(n_1421)
);

AOI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_1376),
.A2(n_1337),
.B1(n_1332),
.B2(n_1350),
.C(n_1334),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1371),
.B(n_1286),
.Y(n_1423)
);

AND2x2_ASAP7_75t_SL g1424 ( 
.A(n_1368),
.B(n_1323),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1386),
.B(n_1347),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1368),
.A2(n_1326),
.B1(n_1323),
.B2(n_1339),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1385),
.B(n_1351),
.C(n_1340),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1358),
.B(n_1304),
.Y(n_1428)
);

NOR3xp33_ASAP7_75t_L g1429 ( 
.A(n_1373),
.B(n_1341),
.C(n_1357),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1359),
.B(n_1301),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1409),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1401),
.B(n_1366),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1409),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1425),
.B(n_1376),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1423),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1423),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1427),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1419),
.B(n_1365),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1427),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1396),
.B(n_1369),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1396),
.B(n_1369),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1428),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1389),
.B(n_1372),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1416),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1419),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1428),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1392),
.B(n_1365),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1399),
.B(n_1367),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1398),
.B(n_1422),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1400),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1416),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1421),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1401),
.B(n_1424),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1416),
.B(n_1379),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1424),
.B(n_1369),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1407),
.B(n_1372),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1395),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1393),
.B(n_1394),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1397),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1442),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1440),
.B(n_1424),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1442),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1449),
.B(n_1383),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1448),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1449),
.B(n_1383),
.Y(n_1465)
);

NOR4xp75_ASAP7_75t_L g1466 ( 
.A(n_1453),
.B(n_1410),
.C(n_1408),
.D(n_1405),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1442),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1442),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1446),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1446),
.Y(n_1470)
);

NAND2xp67_ASAP7_75t_L g1471 ( 
.A(n_1456),
.B(n_1280),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1446),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1437),
.B(n_1413),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1446),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_1434),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1447),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1444),
.B(n_1451),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1458),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1451),
.B(n_1444),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1437),
.B(n_1414),
.Y(n_1481)
);

OAI21xp33_ASAP7_75t_L g1482 ( 
.A1(n_1453),
.A2(n_1418),
.B(n_1390),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1452),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1452),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1457),
.B(n_1383),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1440),
.B(n_1382),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1451),
.B(n_1429),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1452),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1457),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1436),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1437),
.B(n_1415),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1404),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1447),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1439),
.B(n_1377),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1477),
.B(n_1439),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1473),
.B(n_1434),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1482),
.A2(n_1432),
.B1(n_1391),
.B2(n_1444),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1479),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1494),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1483),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1484),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1476),
.A2(n_1432),
.B1(n_1391),
.B2(n_1444),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1463),
.B(n_1445),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1492),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1474),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1488),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1465),
.B(n_1445),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1445),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1493),
.B(n_1447),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1489),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1493),
.B(n_1456),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1474),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1438),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1494),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1461),
.B(n_1433),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1481),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1480),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1481),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1490),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1491),
.B(n_1459),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1480),
.B(n_1451),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1490),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1478),
.Y(n_1524)
);

INVxp67_ASAP7_75t_SL g1525 ( 
.A(n_1478),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1459),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1461),
.B(n_1433),
.Y(n_1527)
);

NAND2xp33_ASAP7_75t_L g1528 ( 
.A(n_1466),
.B(n_1403),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1433),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1487),
.A2(n_1444),
.B1(n_1451),
.B2(n_1403),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1485),
.Y(n_1531)
);

NOR2x1p5_ASAP7_75t_SL g1532 ( 
.A(n_1460),
.B(n_1438),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1486),
.B(n_1459),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1486),
.B(n_1458),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1487),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1462),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1460),
.B(n_1438),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1500),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1497),
.B(n_1280),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1501),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1516),
.B(n_1487),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1502),
.A2(n_1467),
.B(n_1462),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1506),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1524),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1498),
.B(n_1450),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1510),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1518),
.B(n_1451),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1499),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1527),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1495),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1518),
.Y(n_1551)
);

CKINVDCx16_ASAP7_75t_R g1552 ( 
.A(n_1530),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1495),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_L g1555 ( 
.A(n_1528),
.B(n_1417),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1504),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1524),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1450),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1508),
.B(n_1309),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1517),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1511),
.B(n_1475),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1503),
.B(n_1471),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1527),
.B(n_1478),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1535),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1507),
.A2(n_1402),
.B(n_1443),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1522),
.B(n_1464),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1519),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1509),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1522),
.B(n_1529),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1522),
.B(n_1464),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1505),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1515),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1550),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1565),
.B(n_1534),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1565),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1550),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1570),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1558),
.Y(n_1580)
);

NAND2x1_ASAP7_75t_L g1581 ( 
.A(n_1560),
.B(n_1529),
.Y(n_1581)
);

OAI21xp33_ASAP7_75t_L g1582 ( 
.A1(n_1555),
.A2(n_1557),
.B(n_1568),
.Y(n_1582)
);

NOR3xp33_ASAP7_75t_SL g1583 ( 
.A(n_1552),
.B(n_1525),
.C(n_1521),
.Y(n_1583)
);

AOI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1555),
.A2(n_1511),
.B(n_1513),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1553),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1552),
.A2(n_1444),
.B1(n_1526),
.B2(n_1514),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1554),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1554),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1538),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1538),
.Y(n_1590)
);

NAND2x1_ASAP7_75t_L g1591 ( 
.A(n_1560),
.B(n_1505),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1566),
.A2(n_1513),
.B1(n_1444),
.B2(n_1512),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1570),
.Y(n_1593)
);

NOR3xp33_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1561),
.C(n_1539),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1563),
.A2(n_1444),
.B1(n_1512),
.B2(n_1531),
.Y(n_1595)
);

AOI21xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1559),
.A2(n_1509),
.B(n_1533),
.Y(n_1596)
);

AOI21xp33_ASAP7_75t_SL g1597 ( 
.A1(n_1561),
.A2(n_1537),
.B(n_1455),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1548),
.B(n_1532),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1549),
.A2(n_1444),
.B1(n_1455),
.B2(n_1454),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1576),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1576),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1574),
.B(n_1573),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1575),
.B(n_1569),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1589),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1580),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1590),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1579),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1585),
.B(n_1587),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1582),
.B(n_1549),
.Y(n_1610)
);

AOI222xp33_ASAP7_75t_L g1611 ( 
.A1(n_1592),
.A2(n_1569),
.B1(n_1540),
.B2(n_1543),
.C1(n_1546),
.C2(n_1564),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1578),
.B(n_1541),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1593),
.B(n_1551),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1598),
.B(n_1545),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1588),
.B(n_1540),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1584),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1618),
.A2(n_1583),
.B1(n_1592),
.B2(n_1594),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1610),
.A2(n_1584),
.B1(n_1586),
.B2(n_1595),
.Y(n_1620)
);

AOI211x1_ASAP7_75t_L g1621 ( 
.A1(n_1600),
.A2(n_1564),
.B(n_1541),
.C(n_1571),
.Y(n_1621)
);

OAI21xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1611),
.A2(n_1558),
.B(n_1567),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1612),
.B(n_1558),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1601),
.B(n_1615),
.Y(n_1624)
);

NOR4xp25_ASAP7_75t_L g1625 ( 
.A(n_1609),
.B(n_1546),
.C(n_1543),
.D(n_1544),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1602),
.A2(n_1597),
.B1(n_1596),
.B2(n_1542),
.C(n_1581),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1615),
.B(n_1599),
.Y(n_1627)
);

OAI222xp33_ASAP7_75t_L g1628 ( 
.A1(n_1617),
.A2(n_1544),
.B1(n_1547),
.B2(n_1572),
.C1(n_1571),
.C2(n_1567),
.Y(n_1628)
);

NAND4xp25_ASAP7_75t_L g1629 ( 
.A(n_1613),
.B(n_1544),
.C(n_1572),
.D(n_1547),
.Y(n_1629)
);

OAI211xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1603),
.A2(n_1562),
.B(n_1556),
.C(n_1542),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1624),
.B(n_1605),
.C(n_1602),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1629),
.B(n_1614),
.Y(n_1632)
);

NAND4xp75_ASAP7_75t_L g1633 ( 
.A(n_1622),
.B(n_1608),
.C(n_1607),
.D(n_1609),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1621),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1623),
.Y(n_1635)
);

NOR2x1_ASAP7_75t_L g1636 ( 
.A(n_1630),
.B(n_1604),
.Y(n_1636)
);

NOR3xp33_ASAP7_75t_L g1637 ( 
.A(n_1619),
.B(n_1606),
.C(n_1616),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1627),
.Y(n_1638)
);

NOR3xp33_ASAP7_75t_L g1639 ( 
.A(n_1626),
.B(n_1616),
.C(n_1547),
.Y(n_1639)
);

NOR3xp33_ASAP7_75t_L g1640 ( 
.A(n_1628),
.B(n_1547),
.C(n_1562),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1635),
.B(n_1620),
.Y(n_1641)
);

NOR3x1_ASAP7_75t_L g1642 ( 
.A(n_1633),
.B(n_1625),
.C(n_1556),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1537),
.C(n_1276),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1632),
.A2(n_1542),
.B(n_1276),
.C(n_1536),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1636),
.B(n_1523),
.C(n_1520),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1642),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1645),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1641),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1643),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1644),
.A2(n_1638),
.B1(n_1637),
.B2(n_1639),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1641),
.A2(n_1634),
.B1(n_1640),
.B2(n_1455),
.Y(n_1651)
);

NAND4xp25_ASAP7_75t_L g1652 ( 
.A(n_1650),
.B(n_1406),
.C(n_1426),
.D(n_1411),
.Y(n_1652)
);

NOR3xp33_ASAP7_75t_L g1653 ( 
.A(n_1646),
.B(n_1523),
.C(n_1520),
.Y(n_1653)
);

CKINVDCx16_ASAP7_75t_R g1654 ( 
.A(n_1648),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1647),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1649),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1654),
.B(n_1651),
.Y(n_1657)
);

AO211x2_ASAP7_75t_L g1658 ( 
.A1(n_1653),
.A2(n_1471),
.B(n_1467),
.C(n_1472),
.Y(n_1658)
);

NOR2xp67_ASAP7_75t_L g1659 ( 
.A(n_1655),
.B(n_1273),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1657),
.Y(n_1660)
);

NAND4xp25_ASAP7_75t_L g1661 ( 
.A(n_1660),
.B(n_1656),
.C(n_1659),
.D(n_1652),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1661),
.A2(n_1658),
.B1(n_1472),
.B2(n_1470),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1661),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1663),
.B(n_1468),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1662),
.A2(n_1273),
.B(n_1290),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1664),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1665),
.A2(n_1309),
.B(n_1468),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1666),
.A2(n_1470),
.B(n_1469),
.Y(n_1668)
);

AOI322xp5_ASAP7_75t_L g1669 ( 
.A1(n_1668),
.A2(n_1667),
.A3(n_1431),
.B1(n_1455),
.B2(n_1469),
.C1(n_1435),
.C2(n_1441),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_R g1670 ( 
.A1(n_1669),
.A2(n_1298),
.B1(n_1326),
.B2(n_1431),
.C(n_1198),
.Y(n_1670)
);

AOI211xp5_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1430),
.B(n_1420),
.C(n_1412),
.Y(n_1671)
);


endmodule