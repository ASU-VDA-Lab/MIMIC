module fake_jpeg_8032_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_12),
.B(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_8),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_30),
.B1(n_16),
.B2(n_18),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_30),
.B1(n_22),
.B2(n_23),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_57),
.B1(n_26),
.B2(n_21),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_30),
.B1(n_22),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_30),
.B1(n_22),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_22),
.B1(n_16),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_17),
.B(n_19),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_15),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_16),
.B1(n_29),
.B2(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_32),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_15),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_65),
.C(n_53),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_37),
.B1(n_34),
.B2(n_32),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_56),
.B1(n_54),
.B2(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_28),
.B1(n_27),
.B2(n_2),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_28),
.C(n_34),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_20),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_27),
.Y(n_100)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_25),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_74),
.B1(n_79),
.B2(n_56),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_48),
.B(n_41),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_9),
.C(n_1),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_43),
.B1(n_56),
.B2(n_54),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_100),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_43),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_94),
.C(n_103),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_25),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_59),
.B1(n_37),
.B2(n_34),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_104),
.B1(n_62),
.B2(n_67),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_27),
.B(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_101),
.B1(n_68),
.B2(n_28),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_28),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_28),
.B1(n_27),
.B2(n_2),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_113),
.B1(n_115),
.B2(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_116),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_74),
.B1(n_60),
.B2(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_116),
.B1(n_119),
.B2(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_95),
.B1(n_98),
.B2(n_103),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_123),
.B(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_137),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_133),
.B1(n_142),
.B2(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_90),
.B1(n_97),
.B2(n_89),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_81),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_139),
.C(n_140),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_89),
.B(n_1),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_146),
.B(n_9),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_93),
.C(n_96),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_93),
.C(n_79),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_88),
.B1(n_76),
.B2(n_73),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_118),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_27),
.B(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_158),
.Y(n_175)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_153),
.B1(n_155),
.B2(n_145),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_0),
.C(n_4),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_114),
.B1(n_120),
.B2(n_117),
.Y(n_153)
);

NOR4xp25_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_108),
.C(n_125),
.D(n_145),
.Y(n_154)
);

OA21x2_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_135),
.B(n_3),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_114),
.B1(n_126),
.B2(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_0),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_78),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_164),
.B(n_165),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_88),
.B1(n_3),
.B2(n_4),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_133),
.B1(n_128),
.B2(n_4),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_143),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

BUFx12f_ASAP7_75t_SL g185 ( 
.A(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_140),
.B1(n_139),
.B2(n_144),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_180),
.B1(n_161),
.B2(n_164),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_149),
.B1(n_158),
.B2(n_151),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_153),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_176),
.C(n_166),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_6),
.C(n_7),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_188),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_152),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_189),
.C(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_148),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_162),
.C(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_191),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_178),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_185),
.B(n_168),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_196),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_172),
.B(n_175),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_177),
.B(n_192),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_202),
.C(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_179),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_167),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_186),
.B1(n_193),
.B2(n_172),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_206),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_177),
.B1(n_182),
.B2(n_179),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_196),
.C(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_202),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_174),
.B1(n_180),
.B2(n_156),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_200),
.Y(n_211)
);

OAI21x1_ASAP7_75t_SL g217 ( 
.A1(n_211),
.A2(n_207),
.B(n_206),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_214),
.B(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_174),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_195),
.C(n_10),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_218),
.A3(n_213),
.B1(n_212),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_210),
.CI(n_213),
.CON(n_218),
.SN(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_11),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_222),
.C(n_223),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_8),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_219),
.B(n_220),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

OAI21x1_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_224),
.B(n_11),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_12),
.Y(n_228)
);


endmodule