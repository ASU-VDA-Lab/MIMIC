module real_aes_7707_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g181 ( .A1(n_0), .A2(n_182), .B(n_183), .C(n_187), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_1), .B(n_177), .Y(n_188) );
INVx1_ASAP7_75t_L g440 ( .A(n_2), .Y(n_440) );
NAND3xp33_ASAP7_75t_SL g756 ( .A(n_2), .B(n_454), .C(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_3), .B(n_142), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_4), .A2(n_123), .B(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_5), .A2(n_128), .B(n_133), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_6), .A2(n_123), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_7), .B(n_177), .Y(n_483) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_8), .A2(n_156), .B(n_206), .Y(n_205) );
AND2x6_ASAP7_75t_L g128 ( .A(n_9), .B(n_129), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_10), .A2(n_128), .B(n_133), .C(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g538 ( .A(n_11), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_12), .B(n_42), .Y(n_441) );
INVx1_ASAP7_75t_L g754 ( .A(n_12), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_13), .B(n_186), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g103 ( .A1(n_14), .A2(n_104), .B1(n_749), .B2(n_760), .Y(n_103) );
INVx1_ASAP7_75t_L g152 ( .A(n_15), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_16), .B(n_142), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_17), .A2(n_143), .B(n_523), .C(n_525), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_18), .B(n_177), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_19), .B(n_170), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_20), .A2(n_133), .B(n_164), .C(n_169), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_21), .A2(n_185), .B(n_200), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_22), .B(n_186), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_23), .A2(n_78), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_23), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_24), .B(n_186), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_25), .Y(n_464) );
INVx1_ASAP7_75t_L g489 ( .A(n_26), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_27), .A2(n_133), .B(n_169), .C(n_209), .Y(n_208) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_28), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_29), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_30), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_30), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_31), .Y(n_746) );
INVx1_ASAP7_75t_L g565 ( .A(n_32), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_33), .A2(n_123), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g126 ( .A(n_34), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g130 ( .A1(n_35), .A2(n_131), .B(n_136), .C(n_146), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_36), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_37), .A2(n_185), .B(n_480), .C(n_482), .Y(n_479) );
INVxp67_ASAP7_75t_L g566 ( .A(n_38), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_39), .B(n_211), .Y(n_210) );
CKINVDCx14_ASAP7_75t_R g478 ( .A(n_40), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_41), .A2(n_133), .B(n_169), .C(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_42), .B(n_754), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_43), .A2(n_187), .B(n_536), .C(n_537), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_44), .B(n_162), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_45), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_46), .B(n_142), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_47), .B(n_123), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_48), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_49), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_50), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_51), .A2(n_131), .B(n_146), .C(n_220), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g112 ( .A1(n_52), .A2(n_88), .B1(n_113), .B2(n_114), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_52), .Y(n_114) );
INVx1_ASAP7_75t_L g184 ( .A(n_53), .Y(n_184) );
INVx1_ASAP7_75t_L g221 ( .A(n_54), .Y(n_221) );
INVx1_ASAP7_75t_L g501 ( .A(n_55), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_56), .B(n_123), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_57), .Y(n_173) );
CKINVDCx14_ASAP7_75t_R g534 ( .A(n_58), .Y(n_534) );
INVx1_ASAP7_75t_L g129 ( .A(n_59), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_60), .B(n_123), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_61), .B(n_177), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_62), .A2(n_168), .B(n_231), .C(n_233), .Y(n_230) );
INVx1_ASAP7_75t_L g151 ( .A(n_63), .Y(n_151) );
INVx1_ASAP7_75t_SL g481 ( .A(n_64), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_65), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_66), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_67), .B(n_177), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_68), .B(n_143), .Y(n_197) );
INVx1_ASAP7_75t_L g467 ( .A(n_69), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_70), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_71), .B(n_139), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_72), .A2(n_133), .B(n_146), .C(n_257), .Y(n_256) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_73), .Y(n_229) );
INVx1_ASAP7_75t_L g759 ( .A(n_74), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_75), .A2(n_123), .B(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_76), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_77), .A2(n_123), .B(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_78), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_79), .A2(n_162), .B(n_561), .Y(n_560) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_80), .Y(n_486) );
INVx1_ASAP7_75t_L g521 ( .A(n_81), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_82), .B(n_138), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_83), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_84), .A2(n_123), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g524 ( .A(n_85), .Y(n_524) );
INVx2_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
INVx1_ASAP7_75t_L g514 ( .A(n_87), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_88), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_89), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_90), .B(n_186), .Y(n_198) );
OR2x2_ASAP7_75t_L g437 ( .A(n_91), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g450 ( .A(n_91), .B(n_439), .Y(n_450) );
INVx2_ASAP7_75t_L g454 ( .A(n_91), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_92), .A2(n_133), .B(n_146), .C(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_93), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g137 ( .A(n_94), .Y(n_137) );
INVxp67_ASAP7_75t_L g234 ( .A(n_95), .Y(n_234) );
OAI22xp33_ASAP7_75t_SL g110 ( .A1(n_96), .A2(n_111), .B1(n_433), .B2(n_434), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_96), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_97), .B(n_156), .Y(n_539) );
INVx1_ASAP7_75t_L g193 ( .A(n_98), .Y(n_193) );
INVx1_ASAP7_75t_L g258 ( .A(n_99), .Y(n_258) );
INVx2_ASAP7_75t_L g504 ( .A(n_100), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_101), .B(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g223 ( .A(n_102), .B(n_148), .Y(n_223) );
OAI21x1_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_109), .B(n_446), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g748 ( .A(n_107), .Y(n_748) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_435), .B(n_442), .Y(n_109) );
INVx1_ASAP7_75t_L g434 ( .A(n_111), .Y(n_434) );
XOR2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_115), .Y(n_111) );
INVx2_ASAP7_75t_L g451 ( .A(n_115), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_115), .A2(n_738), .B1(n_741), .B2(n_742), .Y(n_737) );
OR3x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_347), .C(n_390), .Y(n_115) );
NAND5xp2_ASAP7_75t_L g116 ( .A(n_117), .B(n_274), .C(n_304), .D(n_321), .E(n_336), .Y(n_116) );
AOI221xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_189), .B1(n_236), .B2(n_242), .C(n_246), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_158), .Y(n_118) );
OR2x2_ASAP7_75t_L g251 ( .A(n_119), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g291 ( .A(n_119), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_119), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_119), .B(n_244), .Y(n_326) );
OR2x2_ASAP7_75t_L g338 ( .A(n_119), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_119), .B(n_297), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_119), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_119), .B(n_275), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_119), .B(n_283), .Y(n_389) );
AND2x2_ASAP7_75t_L g421 ( .A(n_119), .B(n_175), .Y(n_421) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_119), .Y(n_429) );
INVx5_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_120), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g248 ( .A(n_120), .B(n_224), .Y(n_248) );
BUFx2_ASAP7_75t_L g271 ( .A(n_120), .Y(n_271) );
AND2x2_ASAP7_75t_L g300 ( .A(n_120), .B(n_159), .Y(n_300) );
AND2x2_ASAP7_75t_L g355 ( .A(n_120), .B(n_252), .Y(n_355) );
OR2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_153), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_130), .B(n_148), .Y(n_121) );
BUFx2_ASAP7_75t_L g162 ( .A(n_123), .Y(n_162) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_128), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_124), .B(n_128), .Y(n_194) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
INVx1_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
INVx1_ASAP7_75t_L g201 ( .A(n_126), .Y(n_201) );
INVx1_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
INVx3_ASAP7_75t_L g143 ( .A(n_127), .Y(n_143) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_127), .Y(n_186) );
INVx1_ASAP7_75t_L g211 ( .A(n_127), .Y(n_211) );
INVx4_ASAP7_75t_SL g147 ( .A(n_128), .Y(n_147) );
BUFx3_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_SL g179 ( .A1(n_132), .A2(n_147), .B(n_180), .C(n_181), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_132), .A2(n_147), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_132), .A2(n_147), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_132), .A2(n_147), .B(n_501), .C(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_SL g520 ( .A1(n_132), .A2(n_147), .B(n_521), .C(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_132), .A2(n_147), .B(n_534), .C(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_SL g561 ( .A1(n_132), .A2(n_147), .B(n_562), .C(n_563), .Y(n_561) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx3_ASAP7_75t_L g145 ( .A(n_134), .Y(n_145) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_134), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_141), .C(n_144), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_138), .A2(n_144), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_138), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_138), .A2(n_469), .B(n_514), .C(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx4_ASAP7_75t_L g232 ( .A(n_140), .Y(n_232) );
INVx2_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_142), .B(n_234), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_142), .A2(n_167), .B(n_489), .C(n_490), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g564 ( .A1(n_142), .A2(n_232), .B1(n_565), .B2(n_566), .Y(n_564) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_143), .B(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx1_ASAP7_75t_L g525 ( .A(n_145), .Y(n_525) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx1_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_148), .A2(n_218), .B(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_148), .A2(n_194), .B(n_486), .C(n_487), .Y(n_485) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_148), .A2(n_532), .B(n_539), .Y(n_531) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_L g157 ( .A(n_149), .B(n_150), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx3_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_192), .B(n_202), .Y(n_191) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_155), .A2(n_255), .B(n_263), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_155), .B(n_264), .Y(n_263) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_155), .A2(n_463), .B(n_470), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_155), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_155), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_156), .A2(n_207), .B(n_208), .Y(n_206) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_156), .Y(n_226) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_158), .B(n_309), .Y(n_318) );
OAI32xp33_ASAP7_75t_L g332 ( .A1(n_158), .A2(n_268), .A3(n_333), .B1(n_334), .B2(n_335), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_158), .B(n_334), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_158), .B(n_251), .Y(n_375) );
INVx1_ASAP7_75t_SL g404 ( .A(n_158), .Y(n_404) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_158), .B(n_191), .C(n_355), .D(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_175), .Y(n_158) );
INVx5_ASAP7_75t_L g245 ( .A(n_159), .Y(n_245) );
AND2x2_ASAP7_75t_L g275 ( .A(n_159), .B(n_176), .Y(n_275) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_159), .Y(n_354) );
AND2x2_ASAP7_75t_L g424 ( .A(n_159), .B(n_371), .Y(n_424) );
OR2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_172), .Y(n_159) );
AOI21xp5_ASAP7_75t_SL g160 ( .A1(n_161), .A2(n_163), .B(n_170), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .Y(n_164) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_168), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_171), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_174), .A2(n_510), .B(n_516), .Y(n_509) );
AND2x4_ASAP7_75t_L g297 ( .A(n_175), .B(n_245), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_175), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g331 ( .A(n_175), .B(n_252), .Y(n_331) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g244 ( .A(n_176), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g283 ( .A(n_176), .B(n_254), .Y(n_283) );
AND2x2_ASAP7_75t_L g292 ( .A(n_176), .B(n_253), .Y(n_292) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_188), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_185), .B(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g536 ( .A(n_186), .Y(n_536) );
INVx2_ASAP7_75t_L g469 ( .A(n_187), .Y(n_469) );
AOI222xp33_ASAP7_75t_L g360 ( .A1(n_189), .A2(n_361), .B1(n_363), .B2(n_365), .C1(n_368), .C2(n_369), .Y(n_360) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_213), .Y(n_189) );
AND2x2_ASAP7_75t_L g293 ( .A(n_190), .B(n_294), .Y(n_293) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_190), .B(n_271), .C(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_205), .Y(n_190) );
INVx5_ASAP7_75t_SL g241 ( .A(n_191), .Y(n_241) );
OAI322xp33_ASAP7_75t_L g246 ( .A1(n_191), .A2(n_247), .A3(n_249), .B1(n_250), .B2(n_265), .C1(n_268), .C2(n_270), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_191), .B(n_239), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_191), .B(n_225), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_194), .A2(n_464), .B(n_465), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_194), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_199), .A2(n_210), .B(n_212), .Y(n_209) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx2_ASAP7_75t_L g559 ( .A(n_204), .Y(n_559) );
INVx2_ASAP7_75t_L g239 ( .A(n_205), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_205), .B(n_215), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_213), .B(n_278), .Y(n_333) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g312 ( .A(n_214), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
OR2x2_ASAP7_75t_L g240 ( .A(n_215), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_215), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g280 ( .A(n_215), .B(n_225), .Y(n_280) );
AND2x2_ASAP7_75t_L g303 ( .A(n_215), .B(n_239), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_215), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_215), .B(n_278), .Y(n_319) );
AND2x2_ASAP7_75t_L g327 ( .A(n_215), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_215), .B(n_287), .Y(n_377) );
INVx5_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g267 ( .A(n_216), .B(n_241), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_216), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g294 ( .A(n_216), .B(n_225), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_216), .B(n_341), .Y(n_382) );
OR2x2_ASAP7_75t_L g398 ( .A(n_216), .B(n_342), .Y(n_398) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_216), .B(n_359), .Y(n_405) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_216), .Y(n_412) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
AND2x2_ASAP7_75t_L g266 ( .A(n_224), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g316 ( .A(n_224), .B(n_239), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_224), .B(n_241), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_224), .B(n_278), .Y(n_400) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_225), .B(n_241), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_225), .B(n_239), .Y(n_288) );
OR2x2_ASAP7_75t_L g342 ( .A(n_225), .B(n_239), .Y(n_342) );
AND2x2_ASAP7_75t_L g359 ( .A(n_225), .B(n_238), .Y(n_359) );
INVxp67_ASAP7_75t_L g381 ( .A(n_225), .Y(n_381) );
AND2x2_ASAP7_75t_L g408 ( .A(n_225), .B(n_278), .Y(n_408) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_225), .Y(n_415) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_226), .A2(n_476), .B(n_483), .Y(n_475) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_226), .A2(n_499), .B(n_505), .Y(n_498) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_226), .A2(n_519), .B(n_526), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_231), .A2(n_258), .B(n_259), .C(n_260), .Y(n_257) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_232), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_232), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_238), .B(n_289), .Y(n_362) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g278 ( .A(n_239), .B(n_241), .Y(n_278) );
OR2x2_ASAP7_75t_L g345 ( .A(n_239), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
OR2x2_ASAP7_75t_L g350 ( .A(n_240), .B(n_342), .Y(n_350) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g249 ( .A(n_244), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_244), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g250 ( .A(n_245), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_245), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_245), .B(n_252), .Y(n_285) );
INVx2_ASAP7_75t_L g330 ( .A(n_245), .Y(n_330) );
AND2x2_ASAP7_75t_L g343 ( .A(n_245), .B(n_283), .Y(n_343) );
AND2x2_ASAP7_75t_L g368 ( .A(n_245), .B(n_292), .Y(n_368) );
INVx1_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
INVx2_ASAP7_75t_SL g307 ( .A(n_251), .Y(n_307) );
INVx1_ASAP7_75t_L g310 ( .A(n_252), .Y(n_310) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_253), .Y(n_273) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
BUFx2_ASAP7_75t_L g371 ( .A(n_254), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_262), .Y(n_255) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g482 ( .A(n_261), .Y(n_482) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g340 ( .A(n_267), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g346 ( .A(n_267), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_267), .A2(n_349), .B1(n_351), .B2(n_356), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_267), .B(n_359), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_268), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g302 ( .A(n_269), .Y(n_302) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
OR2x2_ASAP7_75t_L g284 ( .A(n_271), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_271), .B(n_275), .Y(n_335) );
AND2x2_ASAP7_75t_L g358 ( .A(n_271), .B(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g334 ( .A(n_273), .Y(n_334) );
AOI211xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_281), .C(n_295), .Y(n_274) );
INVx1_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_275), .A2(n_407), .B1(n_409), .B2(n_410), .C(n_413), .Y(n_406) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g425 ( .A(n_278), .Y(n_425) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g374 ( .A(n_280), .B(n_313), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B(n_286), .C(n_290), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OAI32xp33_ASAP7_75t_L g399 ( .A1(n_288), .A2(n_289), .A3(n_352), .B1(n_389), .B2(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
AND2x2_ASAP7_75t_L g431 ( .A(n_291), .B(n_330), .Y(n_431) );
AND2x2_ASAP7_75t_L g378 ( .A(n_292), .B(n_330), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_292), .B(n_300), .Y(n_396) );
AOI31xp33_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_298), .A3(n_299), .B(n_301), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_297), .B(n_309), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_297), .B(n_307), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_297), .A2(n_327), .B1(n_417), .B2(n_420), .C(n_422), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g322 ( .A(n_302), .B(n_323), .Y(n_322) );
AOI222xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_311), .B1(n_314), .B2(n_317), .C1(n_319), .C2(n_320), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g387 ( .A(n_306), .Y(n_387) );
INVx1_ASAP7_75t_L g409 ( .A(n_309), .Y(n_409) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_312), .A2(n_423), .B1(n_425), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g328 ( .A(n_313), .Y(n_328) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B1(n_327), .B2(n_329), .C(n_332), .Y(n_321) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g366 ( .A(n_324), .B(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g418 ( .A(n_324), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g393 ( .A(n_329), .Y(n_393) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
INVx1_ASAP7_75t_L g339 ( .A(n_331), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_334), .B(n_421), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B1(n_343), .B2(n_344), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g430 ( .A(n_343), .Y(n_430) );
INVxp33_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_345), .B(n_389), .Y(n_388) );
OAI32xp33_ASAP7_75t_L g379 ( .A1(n_346), .A2(n_380), .A3(n_381), .B1(n_382), .B2(n_383), .Y(n_379) );
NAND4xp25_ASAP7_75t_L g347 ( .A(n_348), .B(n_360), .C(n_372), .D(n_384), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NAND2xp33_ASAP7_75t_SL g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_355), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_369), .A2(n_385), .B1(n_402), .B2(n_405), .C(n_406), .Y(n_401) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g420 ( .A(n_371), .B(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B1(n_376), .B2(n_378), .C(n_379), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_381), .B(n_412), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_391), .B(n_401), .C(n_416), .D(n_427), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B(n_397), .C(n_399), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g432 ( .A(n_419), .Y(n_432) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_431), .B(n_432), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g445 ( .A(n_437), .Y(n_445) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_438), .B(n_454), .Y(n_745) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g453 ( .A(n_439), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_442), .A2(n_447), .B(n_747), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI222xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_731), .B1(n_737), .B2(n_743), .C1(n_744), .C2(n_746), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_451), .B1(n_452), .B2(n_455), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g740 ( .A(n_450), .Y(n_740) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx6_ASAP7_75t_L g741 ( .A(n_453), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_455), .Y(n_742) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_456), .B(n_686), .Y(n_455) );
NOR4xp25_ASAP7_75t_L g456 ( .A(n_457), .B(n_623), .C(n_657), .D(n_673), .Y(n_456) );
NAND4xp25_ASAP7_75t_SL g457 ( .A(n_458), .B(n_552), .C(n_587), .D(n_603), .Y(n_457) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_493), .B1(n_527), .B2(n_540), .C1(n_545), .C2(n_551), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI31xp33_ASAP7_75t_L g719 ( .A1(n_460), .A2(n_720), .A3(n_721), .B(n_723), .Y(n_719) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
AND2x2_ASAP7_75t_L g694 ( .A(n_461), .B(n_474), .Y(n_694) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g544 ( .A(n_462), .Y(n_544) );
AND2x2_ASAP7_75t_L g551 ( .A(n_462), .B(n_484), .Y(n_551) );
AND2x2_ASAP7_75t_L g608 ( .A(n_462), .B(n_475), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_472), .B(n_638), .Y(n_637) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_473), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_473), .B(n_555), .Y(n_598) );
AND2x2_ASAP7_75t_L g691 ( .A(n_473), .B(n_631), .Y(n_691) );
OAI321xp33_ASAP7_75t_L g725 ( .A1(n_473), .A2(n_544), .A3(n_698), .B1(n_726), .B2(n_728), .C(n_729), .Y(n_725) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_473), .B(n_530), .C(n_638), .D(n_730), .Y(n_729) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
AND2x2_ASAP7_75t_L g593 ( .A(n_474), .B(n_542), .Y(n_593) );
AND2x2_ASAP7_75t_L g612 ( .A(n_474), .B(n_544), .Y(n_612) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g543 ( .A(n_475), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g568 ( .A(n_475), .B(n_484), .Y(n_568) );
AND2x2_ASAP7_75t_L g654 ( .A(n_475), .B(n_542), .Y(n_654) );
INVx3_ASAP7_75t_SL g542 ( .A(n_484), .Y(n_542) );
AND2x2_ASAP7_75t_L g586 ( .A(n_484), .B(n_573), .Y(n_586) );
OR2x2_ASAP7_75t_L g619 ( .A(n_484), .B(n_544), .Y(n_619) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_484), .Y(n_626) );
AND2x2_ASAP7_75t_L g655 ( .A(n_484), .B(n_543), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_484), .B(n_628), .Y(n_670) );
AND2x2_ASAP7_75t_L g702 ( .A(n_484), .B(n_694), .Y(n_702) );
AND2x2_ASAP7_75t_L g711 ( .A(n_484), .B(n_556), .Y(n_711) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
INVx1_ASAP7_75t_SL g679 ( .A(n_495), .Y(n_679) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g547 ( .A(n_496), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g529 ( .A(n_497), .B(n_508), .Y(n_529) );
AND2x2_ASAP7_75t_L g615 ( .A(n_497), .B(n_531), .Y(n_615) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g585 ( .A(n_498), .B(n_518), .Y(n_585) );
OR2x2_ASAP7_75t_L g596 ( .A(n_498), .B(n_531), .Y(n_596) );
AND2x2_ASAP7_75t_L g622 ( .A(n_498), .B(n_531), .Y(n_622) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_498), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_506), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_506), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g595 ( .A(n_507), .B(n_596), .Y(n_595) );
AOI322xp5_ASAP7_75t_L g681 ( .A1(n_507), .A2(n_585), .A3(n_591), .B1(n_622), .B2(n_672), .C1(n_682), .C2(n_684), .Y(n_681) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_508), .B(n_530), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_508), .B(n_531), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_508), .B(n_548), .Y(n_602) );
AND2x2_ASAP7_75t_L g656 ( .A(n_508), .B(n_622), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_508), .Y(n_660) );
AND2x2_ASAP7_75t_L g672 ( .A(n_508), .B(n_518), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_508), .B(n_547), .Y(n_704) );
INVx4_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g569 ( .A(n_509), .B(n_518), .Y(n_569) );
BUFx3_ASAP7_75t_L g583 ( .A(n_509), .Y(n_583) );
AND3x2_ASAP7_75t_L g665 ( .A(n_509), .B(n_645), .C(n_666), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g528 ( .A(n_518), .B(n_529), .C(n_530), .Y(n_528) );
INVx1_ASAP7_75t_SL g548 ( .A(n_518), .Y(n_548) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_518), .Y(n_650) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g644 ( .A(n_529), .B(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_L g651 ( .A(n_529), .Y(n_651) );
AND2x2_ASAP7_75t_L g689 ( .A(n_530), .B(n_667), .Y(n_689) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g570 ( .A(n_531), .Y(n_570) );
AND2x2_ASAP7_75t_L g645 ( .A(n_531), .B(n_548), .Y(n_645) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
OR2x2_ASAP7_75t_L g589 ( .A(n_542), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g708 ( .A(n_542), .B(n_608), .Y(n_708) );
AND2x2_ASAP7_75t_L g722 ( .A(n_542), .B(n_544), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_543), .B(n_556), .Y(n_663) );
AND2x2_ASAP7_75t_L g710 ( .A(n_543), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g573 ( .A(n_544), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g590 ( .A(n_544), .B(n_556), .Y(n_590) );
INVx1_ASAP7_75t_L g600 ( .A(n_544), .Y(n_600) );
AND2x2_ASAP7_75t_L g631 ( .A(n_544), .B(n_556), .Y(n_631) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_546), .A2(n_674), .B1(n_678), .B2(n_680), .C(n_681), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_L g577 ( .A(n_547), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_550), .B(n_584), .Y(n_727) );
AOI322xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_569), .A3(n_570), .B1(n_571), .B2(n_577), .C1(n_579), .C2(n_586), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_568), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_555), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_555), .B(n_618), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_555), .A2(n_568), .B(n_642), .C(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_555), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_555), .B(n_612), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_555), .B(n_694), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_555), .B(n_722), .Y(n_721) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_556), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_556), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g683 ( .A(n_556), .B(n_570), .Y(n_683) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B(n_567), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_558), .A2(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g575 ( .A(n_560), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_567), .Y(n_576) );
INVx1_ASAP7_75t_L g658 ( .A(n_568), .Y(n_658) );
OAI31xp33_ASAP7_75t_L g668 ( .A1(n_568), .A2(n_593), .A3(n_669), .B(n_671), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_568), .B(n_574), .Y(n_720) );
INVx1_ASAP7_75t_SL g581 ( .A(n_569), .Y(n_581) );
AND2x2_ASAP7_75t_L g614 ( .A(n_569), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g695 ( .A(n_569), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g580 ( .A(n_570), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g605 ( .A(n_570), .Y(n_605) );
AND2x2_ASAP7_75t_L g632 ( .A(n_570), .B(n_585), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_570), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g724 ( .A(n_570), .B(n_672), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_572), .B(n_642), .Y(n_715) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g611 ( .A(n_574), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g629 ( .A(n_574), .Y(n_629) );
NAND2xp33_ASAP7_75t_SL g579 ( .A(n_580), .B(n_582), .Y(n_579) );
OAI211xp5_ASAP7_75t_SL g623 ( .A1(n_581), .A2(n_624), .B(n_630), .C(n_646), .Y(n_623) );
OR2x2_ASAP7_75t_L g698 ( .A(n_581), .B(n_679), .Y(n_698) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
CKINVDCx16_ASAP7_75t_R g635 ( .A(n_583), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_583), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g604 ( .A(n_585), .B(n_605), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .B(n_594), .C(n_597), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g638 ( .A(n_590), .Y(n_638) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_593), .B(n_631), .Y(n_636) );
INVx1_ASAP7_75t_L g642 ( .A(n_593), .Y(n_642) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g601 ( .A(n_596), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g634 ( .A(n_596), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g696 ( .A(n_596), .Y(n_696) );
AOI21xp33_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_599), .B(n_601), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_599), .A2(n_610), .B(n_613), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B(n_609), .C(n_616), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_604), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_607), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_SL g620 ( .A(n_608), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_610), .A2(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_615), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g640 ( .A(n_615), .Y(n_640) );
AOI21xp33_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_620), .B(n_621), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g671 ( .A(n_622), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_628), .B(n_654), .Y(n_680) );
AND2x2_ASAP7_75t_L g693 ( .A(n_628), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g707 ( .A(n_628), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g717 ( .A(n_628), .B(n_655), .Y(n_717) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B(n_633), .C(n_641), .Y(n_630) );
INVx1_ASAP7_75t_L g677 ( .A(n_631), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B1(n_637), .B2(n_639), .Y(n_633) );
OR2x2_ASAP7_75t_L g639 ( .A(n_635), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_635), .B(n_696), .Y(n_718) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g712 ( .A(n_645), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_652), .B1(n_655), .B2(n_656), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g730 ( .A(n_650), .Y(n_730) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g676 ( .A(n_654), .Y(n_676) );
OAI211xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B(n_661), .C(n_668), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_676), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR5xp2_ASAP7_75t_L g686 ( .A(n_687), .B(n_705), .C(n_713), .D(n_719), .E(n_725), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_690), .B(n_692), .C(n_699), .Y(n_687) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B(n_697), .Y(n_692) );
OAI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_702), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_712), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g728 ( .A(n_708), .Y(n_728) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g743 ( .A(n_731), .Y(n_743) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx3_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_SL g760 ( .A(n_751), .Y(n_760) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule