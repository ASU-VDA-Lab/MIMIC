module real_jpeg_18237_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AND2x2_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_0),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_0),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_0),
.B(n_414),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_1),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_1),
.B(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_1),
.B(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_1),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_1),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_1),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_1),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_1),
.B(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_2),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_2),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_3),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_34),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_69),
.Y(n_68)
);

NAND2x1_ASAP7_75t_SL g103 ( 
.A(n_4),
.B(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_105),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_4),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_4),
.B(n_390),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_6),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_6),
.Y(n_261)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_6),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_7),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_7),
.B(n_128),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_7),
.B(n_36),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_7),
.B(n_404),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_32),
.Y(n_31)
);

AOI22x1_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_12),
.B1(n_40),
.B2(n_43),
.Y(n_39)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_8),
.B(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_8),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_9),
.B(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_9),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_9),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_34),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_9),
.B(n_117),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_10),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_10),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_10),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_10),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_10),
.B(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_10),
.Y(n_335)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_11),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_12),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_12),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_12),
.B(n_191),
.Y(n_190)
);

AOI31xp33_ASAP7_75t_L g223 ( 
.A1(n_12),
.A2(n_39),
.A3(n_224),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_12),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_12),
.B(n_83),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_12),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_12),
.B(n_117),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g145 ( 
.A(n_14),
.Y(n_145)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_14),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_15),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_15),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_16),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_376),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_206),
.B(n_375),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_162),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_20),
.B(n_162),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_21),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.C(n_72),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_23),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.C(n_46),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_24),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_26),
.B(n_94),
.Y(n_420)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_27),
.B(n_31),
.C(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_34),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_38),
.A2(n_39),
.B1(n_46),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_41),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_41),
.Y(n_230)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_46),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_52),
.C(n_56),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_47),
.A2(n_48),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_47),
.A2(n_48),
.B1(n_56),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_48),
.B(n_116),
.C(n_142),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_51),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_52),
.B(n_176),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_55),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_56),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_58),
.A2(n_73),
.B1(n_74),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_58),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.C(n_71),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_59),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.C(n_65),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_60),
.A2(n_65),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_60),
.Y(n_221)
);

XNOR2x2_ASAP7_75t_SL g276 ( 
.A(n_60),
.B(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_63),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_65),
.Y(n_222)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_68),
.B(n_71),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_70),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_82),
.C(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_77),
.B(n_232),
.C(n_235),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_77),
.A2(n_90),
.B1(n_235),
.B2(n_236),
.Y(n_361)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_80),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_81),
.Y(n_257)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_138),
.B1(n_160),
.B2(n_161),
.Y(n_86)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_109),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_89),
.B(n_109),
.C(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_91),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_93),
.B(n_98),
.C(n_99),
.Y(n_424)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_95),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.C(n_104),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_104),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2x1_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_122),
.C(n_136),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_110),
.B(n_122),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_116),
.C(n_120),
.Y(n_148)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_121),
.B1(n_142),
.B2(n_146),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_118),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_132),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_123),
.A2(n_132),
.B1(n_133),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_132),
.B(n_254),
.C(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_132),
.A2(n_133),
.B1(n_254),
.B2(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_138),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_147),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_139),
.B(n_148),
.C(n_149),
.Y(n_417)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_142),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_142),
.A2(n_146),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_143),
.B(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_145),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_150),
.B(n_155),
.C(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_154),
.Y(n_401)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_159),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_160),
.B(n_380),
.C(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.C(n_171),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_165),
.B1(n_169),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_201),
.C(n_203),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_173),
.B(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_188),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_SL g264 ( 
.A(n_175),
.B(n_265),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_178),
.B(n_189),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_179),
.B(n_185),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_197),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_190),
.A2(n_193),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_193),
.A2(n_251),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_193),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

XOR2x2_ASAP7_75t_SL g248 ( 
.A(n_197),
.B(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_268),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.C(n_242),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_215),
.Y(n_270)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_239),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_239),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.C(n_231),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_223),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_221),
.B(n_278),
.C(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_232),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_SL g308 ( 
.A(n_233),
.B(n_234),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_233),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_233),
.A2(n_329),
.B1(n_330),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_266),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.C(n_264),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_244),
.B(n_373),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_247),
.B(n_264),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.C(n_262),
.Y(n_247)
);

XOR2x1_ASAP7_75t_L g365 ( 
.A(n_248),
.B(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_253),
.B(n_263),
.Y(n_366)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_369),
.B(n_374),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_355),
.B(n_368),
.Y(n_272)
);

OAI21x1_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_314),
.B(n_354),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_299),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_275),
.B(n_299),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_284),
.C(n_292),
.Y(n_275)
);

XOR2x1_ASAP7_75t_L g348 ( 
.A(n_276),
.B(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_284),
.A2(n_285),
.B1(n_292),
.B2(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_286),
.B(n_289),
.Y(n_319)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

AO22x1_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_293),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_301),
.B(n_302),
.C(n_305),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_306),
.B(n_308),
.C(n_309),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI21x1_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_347),
.B(n_353),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_331),
.B(n_346),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_328),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_328),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_322),
.C(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_338),
.B(n_345),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_336),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_335),
.B(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_SL g353 ( 
.A(n_348),
.B(n_351),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_367),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_367),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_364),
.B2(n_365),
.Y(n_356)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_362),
.B2(n_363),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_359),
.Y(n_371)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_364),
.C(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_372),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_425),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_382),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_416),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_399),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_408),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_413),
.Y(n_408)
);

INVx8_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2x1_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_424),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_419)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_420),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_421),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);


endmodule