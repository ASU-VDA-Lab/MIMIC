module real_jpeg_2593_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_202;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_4),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_43),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_43),
.B1(n_56),
.B2(n_59),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_5),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_7),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_41),
.B1(n_56),
.B2(n_59),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_7),
.B(n_50),
.C(n_56),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_7),
.B(n_33),
.C(n_68),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_7),
.B(n_24),
.C(n_36),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_7),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_7),
.B(n_21),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_7),
.B(n_38),
.Y(n_186)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_104),
.B1(n_224),
.B2(n_225),
.Y(n_12)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_102),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_89),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_15),
.B(n_89),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_63),
.C(n_77),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_16),
.A2(n_63),
.B1(n_64),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_45),
.B2(n_62),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_17),
.A2(n_46),
.B(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_29),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_19),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_19),
.A2(n_29),
.B1(n_61),
.B2(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_24),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_24),
.B(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_27),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_29),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_30),
.A2(n_44),
.B(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_31),
.A2(n_38),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_31),
.A2(n_38),
.B(n_40),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

OA22x2_ASAP7_75t_SL g70 ( 
.A1(n_33),
.A2(n_37),
.B1(n_68),
.B2(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_33),
.B(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_47),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_46),
.A2(n_47),
.B1(n_65),
.B2(n_86),
.Y(n_112)
);

AOI211xp5_ASAP7_75t_SL g126 ( 
.A1(n_46),
.A2(n_84),
.B(n_88),
.C(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_46),
.A2(n_47),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_65),
.Y(n_88)
);

AO21x2_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_55),
.B(n_60),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_116),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_56),
.B(n_162),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_72),
.B(n_76),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_72),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_123),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_65),
.A2(n_84),
.B1(n_86),
.B2(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_118),
.C(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_65),
.A2(n_86),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

AO21x2_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_70),
.B(n_71),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_68),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_70),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_91),
.B1(n_92),
.B2(n_100),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_77),
.A2(n_78),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_87),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_79),
.A2(n_111),
.B1(n_112),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_84),
.B1(n_123),
.B2(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_80),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_119),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_84),
.A2(n_123),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_84),
.A2(n_123),
.B1(n_171),
.B2(n_172),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_84),
.A2(n_86),
.B(n_127),
.C(n_194),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_84),
.A2(n_123),
.B1(n_159),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_87),
.B(n_113),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_85),
.A2(n_87),
.B(n_132),
.Y(n_206)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_104),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_217),
.B(n_223),
.Y(n_104)
);

AOI21x1_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_203),
.B(n_216),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_150),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_136),
.B(n_149),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_151),
.C(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_128),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_128),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_121),
.C(n_125),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_120),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_112),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_118),
.B1(n_147),
.B2(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_117),
.A2(n_118),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_117),
.A2(n_118),
.B1(n_160),
.B2(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_118),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_118),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_123),
.C(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_155),
.C(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_129),
.B(n_131),
.C(n_134),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_146),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_142),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_143),
.A2(n_144),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_166),
.B(n_202),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_163),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_196),
.B(n_201),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_190),
.B(n_195),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_180),
.B(n_189),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_205),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_215),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);


endmodule