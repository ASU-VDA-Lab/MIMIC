module fake_netlist_5_775_n_1616 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1616);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1616;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_21),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_111),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_51),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_93),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_29),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_38),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_57),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_28),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_19),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_96),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_106),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_25),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_18),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_24),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_87),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_54),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_45),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_44),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_48),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_98),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_31),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_1),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_68),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_40),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_22),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_33),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_39),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_118),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_24),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_43),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_92),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_39),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_73),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_56),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_152),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_36),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_123),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_36),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_17),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_62),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_14),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_28),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_53),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_5),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_117),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_29),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_134),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_20),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_64),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_88),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_31),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_22),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_32),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_18),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_78),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_35),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_135),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_46),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_138),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_3),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_105),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_144),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_129),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_40),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_10),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_97),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_27),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_42),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_142),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_4),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_119),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_16),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_69),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_23),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_133),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_14),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_38),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_52),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_45),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_139),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_63),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_80),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_121),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_151),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_15),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_42),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_75),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_141),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_65),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_60),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_131),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_89),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_104),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_109),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_132),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_33),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_26),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_74),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_79),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_113),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_37),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_43),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_13),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_50),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_70),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_95),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_47),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_124),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_91),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_154),
.Y(n_299)
);

BUFx2_ASAP7_75t_SL g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_26),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_7),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_72),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_0),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_0),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_30),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_125),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_76),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_169),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_172),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_169),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_199),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_238),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_296),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_159),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_178),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_191),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_246),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_176),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_176),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_258),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_251),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_193),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_278),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_259),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_297),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_163),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_179),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_187),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_155),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_189),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_194),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_196),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_204),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_206),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_181),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_197),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_155),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_207),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_200),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_218),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_164),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_223),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_253),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_233),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_234),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_170),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_179),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_211),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_258),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_236),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_190),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_242),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_243),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_164),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_254),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_257),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_262),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_216),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_258),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_219),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_199),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_190),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_168),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_265),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_168),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_283),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_289),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_291),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_313),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g383 ( 
.A1(n_372),
.A2(n_212),
.B(n_185),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_337),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_205),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_320),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_313),
.B(n_212),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_293),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_315),
.A2(n_284),
.B1(n_306),
.B2(n_305),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_339),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_293),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_338),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_328),
.A2(n_175),
.B1(n_306),
.B2(n_305),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_316),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_326),
.B(n_205),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_314),
.B(n_213),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_317),
.A2(n_302),
.B1(n_208),
.B2(n_173),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_331),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_213),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_319),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_329),
.B(n_170),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_341),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_360),
.B(n_212),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_199),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_330),
.B(n_170),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_342),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_346),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_370),
.B(n_174),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_309),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_309),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_318),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_349),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_333),
.B(n_156),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_333),
.B(n_174),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_334),
.B(n_156),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_379),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_357),
.Y(n_446)
);

INVxp33_ASAP7_75t_SL g447 ( 
.A(n_406),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_387),
.B(n_359),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_409),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_384),
.B(n_245),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_400),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_415),
.B(n_310),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_384),
.B(n_274),
.Y(n_456)
);

BUFx8_ASAP7_75t_SL g457 ( 
.A(n_437),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_225),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

AO22x2_ASAP7_75t_L g462 ( 
.A1(n_412),
.A2(n_300),
.B1(n_201),
.B2(n_255),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_393),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_423),
.B(n_310),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_400),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_432),
.B(n_353),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_422),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_422),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_392),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_396),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_417),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_199),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_435),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_433),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

AND2x2_ASAP7_75t_SL g484 ( 
.A(n_385),
.B(n_185),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_434),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_441),
.B(n_353),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

AO22x2_ASAP7_75t_L g489 ( 
.A1(n_412),
.A2(n_429),
.B1(n_395),
.B2(n_255),
.Y(n_489)
);

INVx8_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_434),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_435),
.Y(n_492)
);

BUFx8_ASAP7_75t_SL g493 ( 
.A(n_442),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_385),
.A2(n_383),
.B(n_396),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_406),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_395),
.B(n_356),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_L g500 ( 
.A1(n_394),
.A2(n_356),
.B1(n_261),
.B2(n_247),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_436),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_419),
.B(n_347),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_442),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_434),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_419),
.B(n_369),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_430),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_429),
.B(n_371),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_380),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_380),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_436),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_374),
.C(n_351),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

AOI21x1_ASAP7_75t_L g514 ( 
.A1(n_391),
.A2(n_263),
.B(n_201),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_334),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_443),
.B(n_352),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_430),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_413),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_444),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_413),
.B(n_227),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_413),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_402),
.B(n_345),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_398),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_394),
.B(n_374),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_382),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_414),
.A2(n_224),
.B1(n_232),
.B2(n_231),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_443),
.B(n_379),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_443),
.A2(n_294),
.B1(n_263),
.B2(n_325),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_401),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_414),
.B(n_410),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_410),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_382),
.B(n_229),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_443),
.B(n_249),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_416),
.B(n_325),
.C(n_192),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_403),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_416),
.B(n_324),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_436),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_403),
.B(n_271),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_404),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_404),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_382),
.Y(n_549)
);

AO21x2_ASAP7_75t_L g550 ( 
.A1(n_383),
.A2(n_167),
.B(n_166),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_381),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_382),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_405),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_405),
.B(n_311),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_407),
.B(n_354),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_407),
.B(n_332),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_408),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_381),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g559 ( 
.A1(n_383),
.A2(n_186),
.B(n_177),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_381),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_408),
.B(n_249),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_389),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_389),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_418),
.B(n_249),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

AOI22x1_ASAP7_75t_SL g566 ( 
.A1(n_421),
.A2(n_175),
.B1(n_173),
.B2(n_290),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_389),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_421),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_386),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_390),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_386),
.B(n_390),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_390),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_425),
.B(n_335),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_386),
.B(n_230),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_425),
.A2(n_267),
.B(n_266),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_386),
.B(n_239),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_427),
.B(n_240),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_427),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_428),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_440),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_428),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_439),
.Y(n_582)
);

BUFx4f_ASAP7_75t_L g583 ( 
.A(n_424),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_440),
.B(n_244),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_424),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_397),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_397),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_397),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_397),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_452),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_452),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_486),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_467),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_222),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_503),
.B(n_292),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_515),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_521),
.B(n_157),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_471),
.B(n_472),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_471),
.A2(n_260),
.B1(n_270),
.B2(n_268),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_461),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_498),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_506),
.B(n_258),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_461),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_472),
.B(n_199),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_538),
.B(n_354),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_465),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_522),
.A2(n_397),
.B(n_241),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_465),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_525),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_467),
.B(n_355),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_486),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_484),
.B(n_424),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_498),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_523),
.B(n_355),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_469),
.Y(n_617)
);

BUFx12f_ASAP7_75t_L g618 ( 
.A(n_482),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_506),
.B(n_157),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_517),
.B(n_235),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_507),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_484),
.B(n_235),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_499),
.B(n_361),
.C(n_378),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_583),
.B(n_475),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_470),
.Y(n_626)
);

OAI221xp5_ASAP7_75t_L g627 ( 
.A1(n_535),
.A2(n_568),
.B1(n_580),
.B2(n_555),
.C(n_458),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_553),
.B(n_424),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_463),
.B(n_361),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_553),
.B(n_424),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_583),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_523),
.B(n_363),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_475),
.B(n_235),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_476),
.B(n_477),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_555),
.A2(n_367),
.B(n_363),
.C(n_364),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_476),
.B(n_235),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_557),
.B(n_424),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_470),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_557),
.B(n_424),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_477),
.B(n_424),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_485),
.B(n_235),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_485),
.B(n_256),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_490),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_453),
.B(n_279),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_457),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_494),
.A2(n_367),
.B(n_364),
.C(n_378),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_515),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_578),
.B(n_158),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_537),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_490),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_512),
.B(n_290),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_473),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_568),
.B(n_366),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_578),
.B(n_158),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_466),
.B(n_280),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_447),
.A2(n_301),
.B1(n_304),
.B2(n_281),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_543),
.B(n_160),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_160),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_457),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_495),
.B(n_288),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_473),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_586),
.B(n_463),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_496),
.B(n_307),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_491),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_491),
.B(n_258),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_462),
.A2(n_258),
.B1(n_388),
.B2(n_308),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_537),
.A2(n_250),
.B1(n_264),
.B2(n_299),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_474),
.Y(n_668)
);

NAND2x1p5_ASAP7_75t_L g669 ( 
.A(n_504),
.B(n_397),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_502),
.B(n_161),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_527),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_474),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_527),
.B(n_426),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_480),
.B(n_481),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_529),
.B(n_426),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_446),
.B(n_161),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_529),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_532),
.Y(n_678)
);

NOR2xp67_ASAP7_75t_L g679 ( 
.A(n_541),
.B(n_162),
.Y(n_679)
);

NOR2x1p5_ASAP7_75t_L g680 ( 
.A(n_497),
.B(n_301),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_445),
.B(n_162),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_505),
.B(n_366),
.C(n_377),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_459),
.B(n_165),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_532),
.B(n_426),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_536),
.B(n_426),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_462),
.A2(n_388),
.B1(n_426),
.B2(n_304),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_445),
.B(n_165),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_542),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_547),
.B(n_171),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_479),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_445),
.B(n_171),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_519),
.B(n_180),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_554),
.A2(n_368),
.B(n_377),
.C(n_375),
.Y(n_693)
);

BUFx8_ASAP7_75t_L g694 ( 
.A(n_459),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_537),
.B(n_180),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_537),
.B(n_368),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_548),
.B(n_182),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_565),
.B(n_182),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_556),
.B(n_273),
.C(n_188),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_584),
.B(n_183),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_479),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_451),
.B(n_184),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_573),
.A2(n_275),
.B1(n_184),
.B2(n_276),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_554),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_SL g705 ( 
.A1(n_450),
.A2(n_226),
.B1(n_221),
.B2(n_217),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_456),
.B(n_195),
.C(n_198),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_480),
.B(n_275),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_579),
.B(n_276),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_579),
.B(n_277),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_581),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_581),
.B(n_277),
.Y(n_711)
);

NOR2x1p5_ASAP7_75t_L g712 ( 
.A(n_577),
.B(n_202),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_582),
.Y(n_713)
);

BUFx8_ASAP7_75t_L g714 ( 
.A(n_516),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_462),
.A2(n_375),
.B1(n_203),
.B2(n_214),
.Y(n_715)
);

INVxp33_ASAP7_75t_L g716 ( 
.A(n_449),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_582),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_481),
.B(n_295),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_493),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_516),
.B(n_323),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_509),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_509),
.B(n_295),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_516),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_483),
.B(n_287),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_483),
.B(n_492),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_510),
.B(n_513),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_510),
.B(n_287),
.Y(n_727)
);

BUFx8_ASAP7_75t_L g728 ( 
.A(n_534),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_533),
.B(n_210),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_585),
.B(n_282),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_492),
.B(n_501),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_501),
.B(n_298),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_513),
.B(n_298),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_561),
.B(n_215),
.C(n_228),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_500),
.B(n_282),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_534),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_546),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_546),
.B(n_286),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_546),
.A2(n_303),
.B1(n_286),
.B2(n_299),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_546),
.A2(n_303),
.B1(n_252),
.B2(n_269),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_462),
.A2(n_237),
.B1(n_323),
.B2(n_322),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_511),
.B(n_322),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_511),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_454),
.B(n_321),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_493),
.B(n_2),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_540),
.B(n_2),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_464),
.B(n_321),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_544),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_621),
.B(n_611),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_607),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_671),
.B(n_544),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_614),
.A2(n_634),
.B(n_623),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_593),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_613),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_676),
.A2(n_576),
.B1(n_539),
.B2(n_574),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_599),
.B(n_468),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_603),
.Y(n_757)
);

NOR2x2_ASAP7_75t_L g758 ( 
.A(n_735),
.B(n_489),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_716),
.B(n_737),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_664),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_743),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_594),
.B(n_564),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_721),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_723),
.B(n_487),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_748),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_713),
.Y(n_766)
);

NOR2x2_ASAP7_75t_L g767 ( 
.A(n_735),
.B(n_489),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_R g768 ( 
.A(n_618),
.B(n_530),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_632),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_599),
.B(n_566),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_676),
.A2(n_489),
.B1(n_524),
.B2(n_518),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_616),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_710),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_653),
.B(n_597),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_631),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_677),
.B(n_545),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_717),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_645),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_597),
.B(n_530),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_631),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_634),
.A2(n_518),
.B(n_524),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_659),
.B(n_545),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_694),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_678),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_688),
.B(n_530),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_594),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_696),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_658),
.B(n_550),
.Y(n_788)
);

AND3x1_ASAP7_75t_L g789 ( 
.A(n_745),
.B(n_311),
.C(n_312),
.Y(n_789)
);

BUFx5_ASAP7_75t_L g790 ( 
.A(n_674),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_648),
.B(n_312),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_726),
.B(n_549),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_657),
.B(n_549),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_648),
.B(n_550),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_649),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_704),
.B(n_549),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_657),
.B(n_552),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_730),
.B(n_448),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_694),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_730),
.A2(n_569),
.B1(n_552),
.B2(n_520),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_591),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_736),
.A2(n_569),
.B1(n_552),
.B2(n_520),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_744),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_598),
.B(n_569),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_747),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_647),
.B(n_520),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_631),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_600),
.B(n_551),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_600),
.B(n_551),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_SL g811 ( 
.A(n_745),
.B(n_571),
.C(n_5),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_629),
.B(n_572),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_603),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_627),
.A2(n_460),
.B1(n_526),
.B2(n_559),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_674),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_654),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_654),
.B(n_683),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_592),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_683),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_SL g820 ( 
.A(n_705),
.B(n_4),
.C(n_6),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_670),
.A2(n_460),
.B1(n_526),
.B2(n_559),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_662),
.A2(n_460),
.B(n_526),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_742),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_629),
.B(n_560),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_714),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_674),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_SL g827 ( 
.A1(n_646),
.A2(n_478),
.B1(n_563),
.B2(n_562),
.C(n_560),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_702),
.B(n_448),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_643),
.A2(n_526),
.B(n_488),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_658),
.B(n_526),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_674),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_612),
.B(n_559),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_714),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_612),
.Y(n_834)
);

NOR2x1p5_ASAP7_75t_L g835 ( 
.A(n_729),
.B(n_575),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_712),
.Y(n_836)
);

NAND2x1p5_ASAP7_75t_L g837 ( 
.A(n_643),
.B(n_448),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_615),
.B(n_550),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_596),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_719),
.B(n_575),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_728),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_615),
.B(n_570),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_602),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_650),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_670),
.B(n_558),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_737),
.B(n_570),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_605),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_725),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_651),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_689),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_741),
.B(n_562),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_741),
.B(n_563),
.Y(n_852)
);

NOR2x2_ASAP7_75t_L g853 ( 
.A(n_680),
.B(n_558),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_608),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_619),
.B(n_488),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_610),
.Y(n_856)
);

INVx6_ASAP7_75t_L g857 ( 
.A(n_728),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_617),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_619),
.B(n_488),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_674),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_734),
.B(n_679),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_642),
.B(n_567),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_622),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_725),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_731),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_682),
.B(n_572),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_692),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_669),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_601),
.B(n_531),
.Y(n_869)
);

CKINVDCx14_ASAP7_75t_R g870 ( 
.A(n_695),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_669),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_626),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_731),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_638),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_699),
.B(n_531),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_652),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_681),
.B(n_567),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_695),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_681),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_625),
.B(n_590),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_687),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_625),
.B(n_590),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_715),
.B(n_746),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_746),
.A2(n_478),
.B(n_588),
.C(n_587),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_706),
.B(n_531),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_715),
.B(n_589),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_661),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_623),
.B(n_589),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_665),
.A2(n_588),
.B1(n_587),
.B2(n_531),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_668),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_672),
.B(n_508),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_690),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_697),
.Y(n_893)
);

BUFx12f_ASAP7_75t_L g894 ( 
.A(n_595),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_665),
.A2(n_666),
.B1(n_686),
.B2(n_606),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_703),
.B(n_7),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_624),
.B(n_687),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_738),
.B(n_508),
.Y(n_898)
);

NOR2x2_ASAP7_75t_L g899 ( 
.A(n_656),
.B(n_8),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_635),
.B(n_514),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_698),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_701),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_666),
.B(n_606),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_628),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_640),
.B(n_508),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_SL g907 ( 
.A(n_691),
.B(n_8),
.C(n_9),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_604),
.A2(n_508),
.B1(n_488),
.B2(n_514),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_630),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_673),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_722),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_595),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_739),
.B(n_9),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_691),
.B(n_10),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_700),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_SL g916 ( 
.A1(n_740),
.A2(n_667),
.B1(n_686),
.B2(n_727),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_644),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_620),
.B(n_637),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_675),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_733),
.B(n_11),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_693),
.B(n_508),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_620),
.B(n_639),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_684),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_655),
.B(n_488),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_708),
.B(n_711),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_707),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_660),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_685),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_786),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_817),
.A2(n_707),
.B(n_732),
.C(n_724),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_749),
.B(n_732),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_780),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_813),
.Y(n_933)
);

BUFx12f_ASAP7_75t_L g934 ( 
.A(n_825),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_759),
.B(n_709),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_795),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_819),
.B(n_724),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_787),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_756),
.B(n_718),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_753),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_774),
.B(n_718),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_769),
.B(n_750),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_803),
.B(n_693),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_786),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_791),
.B(n_663),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_765),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_860),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_896),
.A2(n_641),
.B(n_636),
.C(n_633),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_780),
.A2(n_633),
.B(n_609),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_754),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_792),
.A2(n_71),
.B(n_150),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_786),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_883),
.A2(n_12),
.B(n_15),
.C(n_16),
.Y(n_953)
);

AOI222xp33_ASAP7_75t_L g954 ( 
.A1(n_913),
.A2(n_12),
.B1(n_17),
.B2(n_20),
.C1(n_21),
.C2(n_25),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_904),
.A2(n_895),
.B1(n_788),
.B2(n_779),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_SL g956 ( 
.A1(n_886),
.A2(n_83),
.B(n_140),
.C(n_128),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_857),
.B(n_81),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_904),
.A2(n_77),
.B(n_122),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_772),
.Y(n_959)
);

INVx3_ASAP7_75t_SL g960 ( 
.A(n_857),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_822),
.A2(n_66),
.B(n_116),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_920),
.A2(n_27),
.B(n_34),
.C(n_37),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_SL g963 ( 
.A1(n_770),
.A2(n_34),
.B1(n_41),
.B2(n_44),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_862),
.A2(n_86),
.B(n_49),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_878),
.B(n_41),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_870),
.B(n_55),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_752),
.A2(n_58),
.B(n_84),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_850),
.B(n_153),
.Y(n_968)
);

AOI21x1_ASAP7_75t_L g969 ( 
.A1(n_798),
.A2(n_90),
.B(n_100),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_850),
.B(n_102),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_926),
.A2(n_115),
.B(n_897),
.C(n_794),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_803),
.B(n_806),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_806),
.B(n_917),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_916),
.A2(n_897),
.B1(n_832),
.B2(n_881),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_860),
.Y(n_975)
);

AOI22x1_ASAP7_75t_SL g976 ( 
.A1(n_778),
.A2(n_772),
.B1(n_787),
.B2(n_881),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_927),
.B(n_867),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_903),
.B(n_901),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_841),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_879),
.B(n_911),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_816),
.B(n_893),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_SL g982 ( 
.A(n_768),
.B(n_914),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_793),
.A2(n_797),
.B1(n_830),
.B2(n_771),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_849),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_872),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_775),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_760),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_855),
.A2(n_859),
.B(n_875),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_804),
.B(n_823),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_879),
.B(n_816),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_915),
.B(n_845),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_801),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_886),
.A2(n_763),
.B1(n_784),
.B2(n_925),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_862),
.A2(n_837),
.B(n_906),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_818),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_752),
.A2(n_888),
.B(n_852),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_821),
.A2(n_814),
.B1(n_757),
.B2(n_838),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_834),
.B(n_764),
.Y(n_998)
);

AND2x2_ASAP7_75t_SL g999 ( 
.A(n_783),
.B(n_833),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_837),
.A2(n_906),
.B(n_922),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_762),
.B(n_861),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_853),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_813),
.B(n_796),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_762),
.B(n_861),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_851),
.A2(n_852),
.B(n_755),
.C(n_877),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_775),
.B(n_808),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_918),
.A2(n_922),
.B(n_924),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_846),
.B(n_805),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_921),
.A2(n_851),
.B1(n_835),
.B2(n_766),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_796),
.B(n_812),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_812),
.B(n_824),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_910),
.A2(n_928),
.B(n_923),
.C(n_919),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_L g1013 ( 
.A1(n_885),
.A2(n_828),
.B(n_898),
.C(n_869),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_860),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_840),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_846),
.B(n_805),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_789),
.B(n_838),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_918),
.A2(n_924),
.B(n_888),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_824),
.B(n_848),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_751),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_864),
.B(n_865),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_907),
.A2(n_811),
.B(n_840),
.C(n_836),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_866),
.A2(n_840),
.B1(n_909),
.B2(n_905),
.Y(n_1023)
);

CKINVDCx8_ASAP7_75t_R g1024 ( 
.A(n_782),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_782),
.B(n_810),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_894),
.B(n_868),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_829),
.A2(n_844),
.B(n_882),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_912),
.A2(n_831),
.B(n_826),
.C(n_815),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_884),
.A2(n_820),
.B(n_807),
.C(n_777),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_751),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_868),
.B(n_871),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_873),
.B(n_809),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_807),
.A2(n_776),
.B(n_785),
.C(n_890),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_782),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_842),
.B(n_773),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_868),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_776),
.A2(n_785),
.B(n_902),
.C(n_810),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_844),
.B(n_826),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_880),
.A2(n_882),
.B(n_891),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_880),
.A2(n_891),
.B(n_781),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_781),
.A2(n_921),
.B(n_809),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_871),
.B(n_842),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_866),
.A2(n_856),
.B(n_843),
.C(n_854),
.Y(n_1043)
);

OAI22x1_ASAP7_75t_L g1044 ( 
.A1(n_758),
.A2(n_767),
.B1(n_899),
.B2(n_802),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_912),
.A2(n_761),
.B(n_892),
.C(n_887),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_839),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_799),
.B(n_815),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_847),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_800),
.A2(n_874),
.B1(n_876),
.B2(n_858),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_863),
.B(n_900),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_900),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_908),
.A2(n_889),
.B(n_900),
.Y(n_1052)
);

OA22x2_ASAP7_75t_L g1053 ( 
.A1(n_827),
.A2(n_497),
.B1(n_394),
.B2(n_528),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_790),
.A2(n_827),
.B(n_643),
.Y(n_1054)
);

O2A1O1Ixp5_ASAP7_75t_L g1055 ( 
.A1(n_790),
.A2(n_817),
.B(n_676),
.C(n_657),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_790),
.A2(n_650),
.B(n_643),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_817),
.A2(n_896),
.B(n_756),
.C(n_819),
.Y(n_1057)
);

NAND3x1_ASAP7_75t_L g1058 ( 
.A(n_990),
.B(n_1004),
.C(n_931),
.Y(n_1058)
);

OA22x2_ASAP7_75t_L g1059 ( 
.A1(n_963),
.A2(n_1044),
.B1(n_959),
.B2(n_936),
.Y(n_1059)
);

O2A1O1Ixp5_ASAP7_75t_L g1060 ( 
.A1(n_1055),
.A2(n_983),
.B(n_939),
.C(n_967),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_991),
.B(n_1057),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_938),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_940),
.Y(n_1063)
);

AO31x2_ASAP7_75t_L g1064 ( 
.A1(n_997),
.A2(n_955),
.A3(n_1005),
.B(n_1054),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_950),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_941),
.B(n_945),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1056),
.A2(n_1007),
.B(n_994),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_973),
.B(n_977),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_937),
.B(n_1020),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_987),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_934),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_929),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_974),
.A2(n_1023),
.B1(n_1009),
.B2(n_1030),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_932),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1018),
.A2(n_1041),
.B(n_1000),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1027),
.A2(n_1039),
.B(n_1040),
.Y(n_1076)
);

AO32x2_ASAP7_75t_L g1077 ( 
.A1(n_963),
.A2(n_1049),
.A3(n_1053),
.B1(n_954),
.B2(n_1009),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_986),
.B(n_932),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_929),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_957),
.B(n_1051),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_972),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_989),
.B(n_1008),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_1052),
.A2(n_971),
.A3(n_1045),
.B(n_1050),
.Y(n_1083)
);

INVx8_ASAP7_75t_L g1084 ( 
.A(n_947),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1016),
.B(n_1011),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_947),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_984),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1010),
.B(n_943),
.Y(n_1088)
);

BUFx12f_ASAP7_75t_L g1089 ( 
.A(n_1002),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_993),
.A2(n_1025),
.B1(n_930),
.B2(n_980),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_996),
.A2(n_948),
.B(n_1029),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_946),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1021),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_970),
.B(n_942),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_992),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_1013),
.A2(n_993),
.B(n_958),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1033),
.A2(n_1037),
.B(n_1012),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_995),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_978),
.B(n_1001),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_SL g1100 ( 
.A1(n_954),
.A2(n_953),
.B(n_965),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1019),
.B(n_1046),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_L g1102 ( 
.A(n_998),
.B(n_968),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_976),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1022),
.A2(n_1043),
.B(n_962),
.C(n_982),
.Y(n_1104)
);

AOI21xp33_ASAP7_75t_L g1105 ( 
.A1(n_1017),
.A2(n_1032),
.B(n_1015),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1048),
.B(n_1035),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_981),
.B(n_964),
.C(n_951),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_SL g1108 ( 
.A(n_935),
.B(n_966),
.C(n_1024),
.Y(n_1108)
);

CKINVDCx16_ASAP7_75t_R g1109 ( 
.A(n_979),
.Y(n_1109)
);

BUFx12f_ASAP7_75t_L g1110 ( 
.A(n_944),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1036),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_988),
.A2(n_949),
.B(n_969),
.Y(n_1112)
);

BUFx2_ASAP7_75t_SL g1113 ( 
.A(n_944),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1035),
.B(n_1003),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_985),
.B(n_952),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_952),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_SL g1117 ( 
.A1(n_1028),
.A2(n_956),
.B(n_961),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_957),
.B(n_999),
.Y(n_1118)
);

AO21x2_ASAP7_75t_L g1119 ( 
.A1(n_1042),
.A2(n_1031),
.B(n_933),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_952),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_1026),
.A2(n_1038),
.B(n_1006),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1006),
.A2(n_1036),
.B(n_975),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1036),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_960),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_975),
.B(n_1014),
.Y(n_1125)
);

AOI211x1_ASAP7_75t_L g1126 ( 
.A1(n_975),
.A2(n_1014),
.B(n_957),
.C(n_1047),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1034),
.B(n_817),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_1034),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1054),
.A2(n_1000),
.B(n_1056),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_938),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1057),
.A2(n_817),
.B(n_756),
.Y(n_1131)
);

AOI221x1_ASAP7_75t_L g1132 ( 
.A1(n_983),
.A2(n_817),
.B1(n_971),
.B2(n_967),
.C(n_953),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_957),
.B(n_857),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_939),
.A2(n_817),
.B1(n_883),
.B2(n_896),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_939),
.A2(n_817),
.B1(n_974),
.B2(n_883),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_940),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_938),
.Y(n_1137)
);

BUFx8_ASAP7_75t_L g1138 ( 
.A(n_934),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1034),
.B(n_786),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_942),
.B(n_774),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1054),
.A2(n_1000),
.B(n_1056),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_939),
.B(n_817),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_932),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_939),
.A2(n_817),
.B1(n_883),
.B2(n_896),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_939),
.B(n_817),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_939),
.B(n_817),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_940),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_929),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_SL g1149 ( 
.A1(n_1029),
.A2(n_993),
.B(n_967),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_942),
.B(n_774),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_940),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_939),
.B(n_817),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1057),
.B(n_817),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1057),
.B(n_817),
.Y(n_1154)
);

AO32x2_ASAP7_75t_L g1155 ( 
.A1(n_955),
.A2(n_997),
.A3(n_983),
.B1(n_963),
.B2(n_916),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_947),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_983),
.A2(n_997),
.A3(n_955),
.B(n_1005),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1057),
.B(n_817),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1055),
.A2(n_817),
.B(n_939),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1055),
.A2(n_955),
.B(n_983),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_983),
.A2(n_997),
.A3(n_955),
.B(n_1005),
.Y(n_1161)
);

BUFx2_ASAP7_75t_SL g1162 ( 
.A(n_929),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_973),
.B(n_450),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_942),
.B(n_774),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1057),
.B(n_817),
.C(n_676),
.Y(n_1165)
);

NAND3x1_ASAP7_75t_L g1166 ( 
.A(n_990),
.B(n_913),
.C(n_745),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1057),
.B(n_817),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_940),
.Y(n_1168)
);

AOI21xp33_ASAP7_75t_L g1169 ( 
.A1(n_1057),
.A2(n_817),
.B(n_756),
.Y(n_1169)
);

NAND3x1_ASAP7_75t_L g1170 ( 
.A(n_990),
.B(n_913),
.C(n_745),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_940),
.Y(n_1171)
);

AND2x2_ASAP7_75t_SL g1172 ( 
.A(n_939),
.B(n_883),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_939),
.B(n_817),
.Y(n_1173)
);

OAI21xp33_ASAP7_75t_SL g1174 ( 
.A1(n_954),
.A2(n_904),
.B(n_895),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_983),
.A2(n_997),
.A3(n_955),
.B(n_1005),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_940),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_942),
.B(n_774),
.Y(n_1177)
);

INVx6_ASAP7_75t_L g1178 ( 
.A(n_929),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1132),
.A2(n_1075),
.A3(n_1097),
.B(n_1067),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1084),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1130),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1142),
.B(n_1145),
.Y(n_1182)
);

BUFx4_ASAP7_75t_SL g1183 ( 
.A(n_1133),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1165),
.A2(n_1169),
.B(n_1154),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1110),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1134),
.A2(n_1144),
.B1(n_1173),
.B2(n_1146),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1084),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1160),
.A2(n_1060),
.B(n_1091),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1134),
.A2(n_1144),
.B1(n_1135),
.B2(n_1172),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1139),
.B(n_1114),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1131),
.B(n_1152),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1124),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1165),
.A2(n_1167),
.B1(n_1158),
.B2(n_1153),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1100),
.A2(n_1131),
.B1(n_1059),
.B2(n_1066),
.Y(n_1194)
);

AND2x6_ASAP7_75t_L g1195 ( 
.A(n_1093),
.B(n_1088),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1084),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1160),
.A2(n_1076),
.B(n_1129),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1140),
.B(n_1150),
.Y(n_1198)
);

AO21x2_ASAP7_75t_L g1199 ( 
.A1(n_1159),
.A2(n_1149),
.B(n_1107),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1100),
.B(n_1061),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1117),
.A2(n_1107),
.B(n_1096),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1147),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1096),
.A2(n_1090),
.B(n_1122),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1085),
.A2(n_1174),
.B(n_1082),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1174),
.A2(n_1104),
.B(n_1069),
.C(n_1155),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1073),
.A2(n_1094),
.B1(n_1081),
.B2(n_1099),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_SL g1207 ( 
.A(n_1124),
.B(n_1109),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1171),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1130),
.B(n_1137),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1127),
.B(n_1163),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1074),
.A2(n_1143),
.B(n_1176),
.Y(n_1211)
);

BUFx2_ASAP7_75t_SL g1212 ( 
.A(n_1128),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1063),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1074),
.A2(n_1143),
.B(n_1151),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1138),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1166),
.A2(n_1170),
.B1(n_1058),
.B2(n_1108),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_1089),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1105),
.A2(n_1133),
.B1(n_1102),
.B2(n_1164),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1177),
.B(n_1118),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1068),
.B(n_1137),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1138),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1102),
.A2(n_1136),
.B(n_1168),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1065),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1087),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1101),
.A2(n_1064),
.B(n_1098),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1119),
.A2(n_1133),
.B(n_1175),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1086),
.Y(n_1227)
);

NAND2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1156),
.B(n_1139),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1078),
.A2(n_1095),
.B(n_1115),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1092),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1157),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1106),
.B(n_1062),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1156),
.A2(n_1126),
.B(n_1155),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1119),
.A2(n_1125),
.B(n_1155),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1126),
.B(n_1080),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1116),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1111),
.A2(n_1123),
.B(n_1083),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1157),
.A2(n_1161),
.B(n_1175),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1157),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1072),
.B(n_1148),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1080),
.A2(n_1120),
.B1(n_1103),
.B2(n_1178),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1077),
.A2(n_1113),
.B(n_1162),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1071),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1080),
.A2(n_1077),
.B(n_1178),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1072),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1077),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1079),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1079),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1148),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1134),
.A2(n_1144),
.B1(n_817),
.B2(n_1142),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1130),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1124),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1140),
.B(n_1150),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1165),
.A2(n_817),
.B(n_676),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1070),
.Y(n_1255)
);

INVx8_ASAP7_75t_L g1256 ( 
.A(n_1084),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1134),
.A2(n_1144),
.B1(n_1145),
.B2(n_1142),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1066),
.B(n_1130),
.Y(n_1258)
);

O2A1O1Ixp5_ASAP7_75t_L g1259 ( 
.A1(n_1169),
.A2(n_1060),
.B(n_1160),
.C(n_1158),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1134),
.A2(n_1144),
.B1(n_817),
.B2(n_1142),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1172),
.A2(n_883),
.B1(n_963),
.B2(n_1135),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1139),
.B(n_1114),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1154),
.A2(n_883),
.B1(n_1144),
.B2(n_1134),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1112),
.A2(n_1141),
.B(n_1129),
.Y(n_1264)
);

AOI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1165),
.A2(n_817),
.B(n_1154),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1070),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1084),
.Y(n_1267)
);

AND2x2_ASAP7_75t_SL g1268 ( 
.A(n_1172),
.B(n_1144),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1140),
.B(n_1150),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1154),
.A2(n_883),
.B1(n_1144),
.B2(n_1134),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1084),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1070),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1121),
.B(n_932),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1070),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1132),
.A2(n_1075),
.A3(n_1097),
.B(n_1067),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1134),
.B(n_1144),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1067),
.A2(n_1075),
.B(n_1097),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1070),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1134),
.A2(n_1144),
.B(n_817),
.C(n_1174),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1070),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1134),
.A2(n_1144),
.B1(n_817),
.B2(n_1142),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1110),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1070),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1070),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1070),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1138),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1160),
.A2(n_1097),
.B(n_1075),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1204),
.B(n_1200),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1181),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1258),
.B(n_1209),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1279),
.A2(n_1254),
.B(n_1250),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1213),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1219),
.B(n_1198),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1201),
.A2(n_1259),
.B(n_1203),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1253),
.B(n_1269),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1232),
.B(n_1210),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1210),
.B(n_1220),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1251),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1200),
.B(n_1191),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1265),
.A2(n_1184),
.B(n_1279),
.C(n_1281),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1223),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1193),
.A2(n_1244),
.B(n_1226),
.C(n_1218),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1259),
.A2(n_1277),
.B(n_1264),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1185),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1215),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1260),
.A2(n_1194),
.B(n_1186),
.C(n_1257),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1235),
.B(n_1190),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1251),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1261),
.A2(n_1263),
.B1(n_1270),
.B2(n_1189),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1194),
.A2(n_1257),
.B(n_1205),
.C(n_1182),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1205),
.B(n_1276),
.Y(n_1312)
);

O2A1O1Ixp5_ASAP7_75t_L g1313 ( 
.A1(n_1276),
.A2(n_1238),
.B(n_1231),
.C(n_1239),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1224),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1236),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1193),
.B(n_1206),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1206),
.B(n_1263),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1235),
.A2(n_1216),
.B(n_1187),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1262),
.B(n_1268),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1261),
.A2(n_1189),
.B(n_1268),
.C(n_1218),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1241),
.A2(n_1252),
.B(n_1192),
.C(n_1233),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1221),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1221),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1235),
.A2(n_1242),
.B1(n_1246),
.B2(n_1280),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1207),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1246),
.B(n_1195),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1243),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1215),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1199),
.A2(n_1274),
.B(n_1283),
.C(n_1255),
.Y(n_1329)
);

O2A1O1Ixp5_ASAP7_75t_L g1330 ( 
.A1(n_1284),
.A2(n_1285),
.B(n_1278),
.C(n_1208),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1271),
.B(n_1245),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1202),
.B(n_1272),
.Y(n_1332)
);

O2A1O1Ixp5_ASAP7_75t_L g1333 ( 
.A1(n_1266),
.A2(n_1267),
.B(n_1230),
.C(n_1247),
.Y(n_1333)
);

AOI221xp5_ASAP7_75t_L g1334 ( 
.A1(n_1199),
.A2(n_1212),
.B1(n_1185),
.B2(n_1282),
.C(n_1286),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1183),
.A2(n_1267),
.B(n_1287),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1195),
.B(n_1225),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1282),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1195),
.B(n_1225),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1242),
.A2(n_1188),
.B1(n_1222),
.B2(n_1228),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1195),
.B(n_1188),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1229),
.A2(n_1211),
.B(n_1214),
.C(n_1237),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1234),
.B(n_1179),
.Y(n_1342)
);

OA22x2_ASAP7_75t_L g1343 ( 
.A1(n_1248),
.A2(n_1249),
.B1(n_1243),
.B2(n_1217),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1228),
.B(n_1240),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1227),
.A2(n_1180),
.B1(n_1196),
.B2(n_1256),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1180),
.B(n_1196),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1179),
.A2(n_1275),
.B(n_1197),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1273),
.A2(n_1275),
.B(n_1227),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1273),
.A2(n_1227),
.B(n_1256),
.Y(n_1349)
);

AND2x6_ASAP7_75t_L g1350 ( 
.A(n_1231),
.B(n_1239),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1221),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1224),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1204),
.B(n_1200),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1204),
.B(n_1200),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1201),
.A2(n_1259),
.B(n_1203),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1204),
.B(n_1200),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1258),
.B(n_1209),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1310),
.A2(n_1317),
.B1(n_1299),
.B2(n_1316),
.Y(n_1358)
);

INVxp33_ASAP7_75t_L g1359 ( 
.A(n_1296),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1308),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1340),
.B(n_1347),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1350),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1308),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1350),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1292),
.Y(n_1365)
);

CKINVDCx14_ASAP7_75t_R g1366 ( 
.A(n_1306),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1310),
.A2(n_1312),
.B1(n_1317),
.B2(n_1353),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1347),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1288),
.B(n_1353),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1327),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1339),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1342),
.B(n_1336),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1339),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1335),
.B(n_1348),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1336),
.B(n_1338),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1288),
.A2(n_1354),
.B1(n_1356),
.B2(n_1312),
.Y(n_1377)
);

BUFx2_ASAP7_75t_SL g1378 ( 
.A(n_1343),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1326),
.B(n_1338),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1307),
.A2(n_1311),
.B(n_1301),
.Y(n_1380)
);

NAND2xp33_ASAP7_75t_SL g1381 ( 
.A(n_1354),
.B(n_1356),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1326),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1313),
.A2(n_1341),
.B(n_1324),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1289),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1316),
.A2(n_1297),
.B1(n_1334),
.B2(n_1357),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1307),
.A2(n_1320),
.B(n_1345),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1324),
.A2(n_1333),
.B(n_1330),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1298),
.B(n_1309),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1303),
.A2(n_1329),
.B(n_1291),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_1315),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1290),
.A2(n_1295),
.B1(n_1293),
.B2(n_1325),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1294),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1294),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1332),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1355),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1379),
.B(n_1355),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1370),
.B(n_1300),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1376),
.B(n_1304),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1376),
.B(n_1314),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1370),
.B(n_1319),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1369),
.Y(n_1401)
);

NOR2x1_ASAP7_75t_SL g1402 ( 
.A(n_1375),
.B(n_1345),
.Y(n_1402)
);

CKINVDCx6p67_ASAP7_75t_R g1403 ( 
.A(n_1378),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1365),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1375),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1365),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1376),
.B(n_1352),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1367),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1379),
.B(n_1343),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1361),
.B(n_1318),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1362),
.B(n_1349),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1377),
.B(n_1321),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1361),
.B(n_1344),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1373),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1364),
.B(n_1346),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1361),
.B(n_1331),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1413),
.B(n_1382),
.Y(n_1417)
);

AOI21xp33_ASAP7_75t_L g1418 ( 
.A1(n_1412),
.A2(n_1368),
.B(n_1389),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1404),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1412),
.A2(n_1380),
.B1(n_1358),
.B2(n_1368),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1403),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1403),
.A2(n_1358),
.B1(n_1386),
.B2(n_1385),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1414),
.B(n_1373),
.Y(n_1423)
);

OAI211xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1399),
.A2(n_1377),
.B(n_1385),
.C(n_1391),
.Y(n_1424)
);

OAI31xp33_ASAP7_75t_L g1425 ( 
.A1(n_1405),
.A2(n_1381),
.A3(n_1372),
.B(n_1374),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1403),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1404),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1405),
.B(n_1375),
.Y(n_1428)
);

AND2x2_ASAP7_75t_SL g1429 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1406),
.Y(n_1430)
);

OAI211xp5_ASAP7_75t_L g1431 ( 
.A1(n_1399),
.A2(n_1374),
.B(n_1372),
.C(n_1381),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1407),
.A2(n_1378),
.B1(n_1366),
.B2(n_1391),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1410),
.A2(n_1366),
.B(n_1359),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1414),
.Y(n_1434)
);

AOI211xp5_ASAP7_75t_L g1435 ( 
.A1(n_1410),
.A2(n_1359),
.B(n_1382),
.C(n_1388),
.Y(n_1435)
);

OAI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1405),
.A2(n_1375),
.B1(n_1305),
.B2(n_1390),
.C(n_1373),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_SL g1437 ( 
.A(n_1399),
.B(n_1328),
.C(n_1388),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1401),
.A2(n_1395),
.B(n_1393),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1407),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1407),
.A2(n_1375),
.B1(n_1400),
.B2(n_1397),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1415),
.Y(n_1441)
);

OAI211xp5_ASAP7_75t_L g1442 ( 
.A1(n_1397),
.A2(n_1383),
.B(n_1387),
.C(n_1384),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1408),
.Y(n_1443)
);

OAI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1405),
.A2(n_1383),
.B(n_1387),
.C(n_1384),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1400),
.A2(n_1375),
.B1(n_1360),
.B2(n_1363),
.Y(n_1445)
);

INVx5_ASAP7_75t_SL g1446 ( 
.A(n_1411),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1413),
.B(n_1416),
.Y(n_1447)
);

OAI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1398),
.A2(n_1360),
.B1(n_1363),
.B2(n_1394),
.C(n_1337),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1418),
.B(n_1409),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1421),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1428),
.B(n_1402),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1444),
.A2(n_1392),
.B(n_1393),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1419),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1427),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1434),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1421),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1438),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1426),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1428),
.B(n_1383),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1429),
.B(n_1396),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1426),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1430),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1428),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1443),
.Y(n_1464)
);

INVx4_ASAP7_75t_SL g1465 ( 
.A(n_1441),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1429),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1423),
.B(n_1398),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1447),
.B(n_1409),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1423),
.Y(n_1469)
);

INVx5_ASAP7_75t_L g1470 ( 
.A(n_1446),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1453),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1453),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1466),
.B(n_1468),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1449),
.A2(n_1420),
.B1(n_1422),
.B2(n_1442),
.C(n_1440),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1454),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1458),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1449),
.A2(n_1424),
.B(n_1431),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_L g1479 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1469),
.B(n_1455),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1450),
.B(n_1435),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1455),
.B(n_1417),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1456),
.B(n_1433),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1457),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1458),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1462),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1457),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1466),
.B(n_1441),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1470),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1464),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1450),
.B(n_1439),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1457),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1466),
.B(n_1447),
.Y(n_1494)
);

BUFx2_ASAP7_75t_SL g1495 ( 
.A(n_1470),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1458),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1456),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1463),
.A2(n_1389),
.B1(n_1432),
.B2(n_1425),
.Y(n_1498)
);

AND2x2_ASAP7_75t_SL g1499 ( 
.A(n_1452),
.B(n_1383),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1461),
.B(n_1371),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1468),
.B(n_1439),
.Y(n_1501)
);

AOI31xp33_ASAP7_75t_L g1502 ( 
.A1(n_1451),
.A2(n_1436),
.A3(n_1445),
.B(n_1448),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1471),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1471),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1477),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1472),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1480),
.B(n_1467),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1479),
.A2(n_1461),
.B(n_1452),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1472),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1480),
.B(n_1467),
.Y(n_1512)
);

NOR2xp67_ASAP7_75t_SL g1513 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1475),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1478),
.B(n_1468),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1475),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1482),
.B(n_1467),
.Y(n_1517)
);

NAND2xp33_ASAP7_75t_L g1518 ( 
.A(n_1474),
.B(n_1470),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1498),
.A2(n_1483),
.B1(n_1481),
.B2(n_1492),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1483),
.A2(n_1463),
.B1(n_1459),
.B2(n_1470),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1486),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1477),
.B(n_1465),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1473),
.B(n_1465),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1497),
.B(n_1465),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1487),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1501),
.B(n_1460),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1473),
.B(n_1460),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1497),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_SL g1529 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1476),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1494),
.B(n_1465),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1506),
.B(n_1500),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1506),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1521),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1528),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1505),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1504),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1511),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1530),
.B(n_1515),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1529),
.B(n_1496),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1524),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1522),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1518),
.A2(n_1389),
.B1(n_1499),
.B2(n_1484),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1528),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1511),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1523),
.B(n_1494),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1509),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1512),
.B(n_1491),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1514),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1517),
.B(n_1527),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1522),
.B(n_1470),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1523),
.B(n_1476),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1531),
.B(n_1484),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1544),
.A2(n_1519),
.B(n_1510),
.Y(n_1556)
);

XNOR2xp5_ASAP7_75t_L g1557 ( 
.A(n_1554),
.B(n_1322),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1541),
.A2(n_1529),
.B(n_1520),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1547),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1547),
.Y(n_1560)
);

AOI31xp33_ASAP7_75t_L g1561 ( 
.A1(n_1532),
.A2(n_1504),
.A3(n_1508),
.B(n_1531),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1549),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1549),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1533),
.B(n_1508),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1552),
.B(n_1526),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1534),
.B(n_1503),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1532),
.A2(n_1518),
.B(n_1502),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1548),
.A2(n_1522),
.B1(n_1524),
.B2(n_1489),
.Y(n_1568)
);

OAI21xp33_ASAP7_75t_L g1569 ( 
.A1(n_1540),
.A2(n_1499),
.B(n_1489),
.Y(n_1569)
);

OAI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1544),
.A2(n_1490),
.B1(n_1513),
.B2(n_1463),
.C(n_1517),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1535),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1565),
.B(n_1564),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1557),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1567),
.B(n_1524),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1571),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1561),
.B(n_1538),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1559),
.B(n_1555),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1560),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1562),
.B(n_1552),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1563),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1576),
.A2(n_1556),
.B1(n_1554),
.B2(n_1555),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1574),
.A2(n_1558),
.B(n_1553),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1573),
.A2(n_1568),
.B(n_1548),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1575),
.A2(n_1569),
.B1(n_1570),
.B2(n_1566),
.C(n_1542),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1573),
.B(n_1543),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1577),
.B(n_1543),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1579),
.B(n_1543),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1578),
.Y(n_1588)
);

NOR2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1572),
.B(n_1545),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1585),
.B(n_1580),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1589),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1587),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1583),
.B(n_1513),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1590),
.B(n_1581),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1591),
.B(n_1582),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1593),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1592),
.B(n_1584),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1592),
.B(n_1586),
.Y(n_1598)
);

OAI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1597),
.A2(n_1588),
.B1(n_1490),
.B2(n_1551),
.C(n_1536),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1598),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_SL g1601 ( 
.A(n_1596),
.B(n_1351),
.C(n_1323),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1595),
.Y(n_1602)
);

BUFx10_ASAP7_75t_L g1603 ( 
.A(n_1600),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1602),
.B(n_1594),
.Y(n_1604)
);

AOI31xp33_ASAP7_75t_L g1605 ( 
.A1(n_1601),
.A2(n_1541),
.A3(n_1551),
.B(n_1539),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1603),
.Y(n_1606)
);

AOI322xp5_ASAP7_75t_L g1607 ( 
.A1(n_1606),
.A2(n_1604),
.A3(n_1541),
.B1(n_1605),
.B2(n_1546),
.C1(n_1539),
.C2(n_1537),
.Y(n_1607)
);

XNOR2xp5_ASAP7_75t_L g1608 ( 
.A(n_1607),
.B(n_1599),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1608),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1609),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1610),
.B(n_1606),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1611),
.A2(n_1606),
.B(n_1546),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1612),
.B(n_1550),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1613),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1614),
.A2(n_1516),
.B1(n_1525),
.B2(n_1507),
.Y(n_1615)
);

AOI211xp5_ASAP7_75t_L g1616 ( 
.A1(n_1615),
.A2(n_1485),
.B(n_1493),
.C(n_1488),
.Y(n_1616)
);


endmodule