module fake_jpeg_13470_n_77 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_16),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_49),
.B1(n_54),
.B2(n_41),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_53),
.B(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_60),
.B(n_51),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

OAI321xp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_51),
.A3(n_24),
.B1(n_38),
.B2(n_28),
.C(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_39),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_66),
.A2(n_45),
.B1(n_23),
.B2(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_22),
.C(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_42),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_43),
.A3(n_31),
.B1(n_34),
.B2(n_52),
.C1(n_27),
.C2(n_32),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_74),
.B1(n_56),
.B2(n_48),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_40),
.CI(n_26),
.CON(n_74),
.SN(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_55),
.C(n_59),
.Y(n_76)
);

BUFx24_ASAP7_75t_SL g77 ( 
.A(n_76),
.Y(n_77)
);


endmodule