module fake_netlist_6_1701_n_63 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_10, n_63);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_63;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_24;
wire n_21;
wire n_18;
wire n_37;
wire n_33;
wire n_54;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_60;
wire n_59;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_17;
wire n_58;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_43;
wire n_19;
wire n_47;
wire n_48;
wire n_29;
wire n_62;
wire n_31;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_16),
.B(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AND2x6_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_29),
.B1(n_23),
.B2(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_25),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_18),
.B(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_21),
.Y(n_38)
);

AO22x2_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI21x1_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_28),
.B(n_27),
.Y(n_45)
);

AO21x2_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_30),
.B(n_28),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_31),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_41),
.B(n_43),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_49),
.C(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_46),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_55),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_46),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_22),
.B1(n_45),
.B2(n_46),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_R g60 ( 
.A(n_57),
.B(n_45),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

OR2x6_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_59),
.Y(n_63)
);


endmodule