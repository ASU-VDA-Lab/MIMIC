module real_aes_7533_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_252;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g481 ( .A1(n_0), .A2(n_136), .B(n_482), .C(n_485), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_1), .B(n_476), .Y(n_487) );
INVx1_ASAP7_75t_L g429 ( .A(n_2), .Y(n_429) );
INVx1_ASAP7_75t_L g174 ( .A(n_3), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_4), .B(n_137), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g113 ( .A1(n_5), .A2(n_97), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_5), .Y(n_115) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_5), .A2(n_115), .B1(n_116), .B2(n_447), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_6), .A2(n_461), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_7), .A2(n_143), .B(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_8), .A2(n_40), .B1(n_140), .B2(n_192), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_9), .B(n_143), .Y(n_160) );
AND2x6_ASAP7_75t_L g145 ( .A(n_10), .B(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_11), .A2(n_145), .B(n_464), .C(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_12), .B(n_41), .Y(n_430) );
INVx1_ASAP7_75t_L g748 ( .A(n_12), .Y(n_748) );
INVx1_ASAP7_75t_L g127 ( .A(n_13), .Y(n_127) );
INVx1_ASAP7_75t_L g166 ( .A(n_14), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_15), .B(n_133), .Y(n_186) );
AOI321xp33_ASAP7_75t_L g110 ( .A1(n_16), .A2(n_111), .A3(n_424), .B1(n_431), .B2(n_432), .C(n_434), .Y(n_110) );
INVx1_ASAP7_75t_L g431 ( .A(n_16), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_17), .B(n_137), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_18), .B(n_123), .Y(n_122) );
AO32x2_ASAP7_75t_L g203 ( .A1(n_19), .A2(n_143), .A3(n_144), .B1(n_163), .B2(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_20), .B(n_140), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_21), .B(n_123), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_22), .A2(n_56), .B1(n_140), .B2(n_192), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g200 ( .A1(n_23), .A2(n_81), .B1(n_133), .B2(n_140), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_24), .B(n_140), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_25), .A2(n_144), .B(n_464), .C(n_466), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_26), .A2(n_144), .B(n_464), .C(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_27), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_28), .A2(n_98), .B1(n_441), .B2(n_442), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_28), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_29), .B(n_182), .Y(n_240) );
AOI222xp33_ASAP7_75t_SL g438 ( .A1(n_30), .A2(n_439), .B1(n_445), .B2(n_737), .C1(n_738), .C2(n_740), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_31), .A2(n_461), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_32), .B(n_182), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g104 ( .A1(n_33), .A2(n_105), .B1(n_743), .B2(n_754), .Y(n_104) );
INVx2_ASAP7_75t_L g135 ( .A(n_34), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_35), .A2(n_496), .B(n_497), .C(n_501), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_36), .B(n_140), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_37), .B(n_182), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g439 ( .A1(n_38), .A2(n_440), .B1(n_443), .B2(n_444), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_38), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_39), .B(n_188), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_41), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_42), .B(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_43), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_44), .B(n_137), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_45), .B(n_461), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_46), .A2(n_496), .B(n_501), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_47), .B(n_140), .Y(n_153) );
INVx1_ASAP7_75t_L g483 ( .A(n_48), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g111 ( .A1(n_49), .A2(n_112), .B1(n_422), .B2(n_423), .Y(n_111) );
INVx1_ASAP7_75t_L g423 ( .A(n_49), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_50), .A2(n_89), .B1(n_192), .B2(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g522 ( .A(n_51), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_52), .B(n_140), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_53), .B(n_140), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_54), .B(n_461), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_55), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_SL g139 ( .A1(n_57), .A2(n_61), .B1(n_133), .B2(n_140), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_58), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_59), .B(n_140), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_60), .B(n_140), .Y(n_239) );
INVx1_ASAP7_75t_L g146 ( .A(n_62), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_63), .B(n_461), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_64), .B(n_476), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_65), .A2(n_158), .B(n_169), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_66), .B(n_140), .Y(n_175) );
INVx1_ASAP7_75t_L g126 ( .A(n_67), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_68), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_69), .B(n_137), .Y(n_499) );
AO32x2_ASAP7_75t_L g196 ( .A1(n_70), .A2(n_143), .A3(n_144), .B1(n_197), .B2(n_201), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_71), .B(n_138), .Y(n_533) );
INVx1_ASAP7_75t_L g238 ( .A(n_72), .Y(n_238) );
INVx1_ASAP7_75t_L g214 ( .A(n_73), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_74), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_75), .B(n_468), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_76), .A2(n_464), .B(n_501), .C(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_77), .B(n_133), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_78), .Y(n_509) );
INVx1_ASAP7_75t_L g753 ( .A(n_79), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_80), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_82), .B(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_83), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_84), .B(n_133), .Y(n_218) );
INVx2_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_86), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_87), .B(n_130), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_88), .B(n_133), .Y(n_154) );
OR2x2_ASAP7_75t_L g426 ( .A(n_90), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g450 ( .A(n_90), .B(n_428), .Y(n_450) );
INVx2_ASAP7_75t_L g736 ( .A(n_90), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_91), .A2(n_103), .B1(n_133), .B2(n_134), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_92), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_93), .B(n_461), .Y(n_494) );
INVx1_ASAP7_75t_L g498 ( .A(n_94), .Y(n_498) );
INVxp67_ASAP7_75t_L g512 ( .A(n_95), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_96), .B(n_133), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_97), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_98), .Y(n_441) );
INVx1_ASAP7_75t_L g529 ( .A(n_99), .Y(n_529) );
INVx1_ASAP7_75t_L g558 ( .A(n_100), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_101), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g524 ( .A(n_102), .B(n_182), .Y(n_524) );
AOI22x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B1(n_436), .B2(n_438), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_SL g437 ( .A(n_108), .Y(n_437) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_111), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g422 ( .A(n_112), .Y(n_422) );
XNOR2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
INVx2_ASAP7_75t_L g447 ( .A(n_116), .Y(n_447) );
AND2x2_ASAP7_75t_SL g116 ( .A(n_117), .B(n_356), .Y(n_116) );
NOR5xp2_ASAP7_75t_L g117 ( .A(n_118), .B(n_269), .C(n_315), .D(n_328), .E(n_340), .Y(n_117) );
OAI211xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_177), .B(n_223), .C(n_250), .Y(n_118) );
INVx1_ASAP7_75t_SL g351 ( .A(n_119), .Y(n_351) );
OR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_147), .Y(n_119) );
AND2x2_ASAP7_75t_L g275 ( .A(n_120), .B(n_148), .Y(n_275) );
AND2x2_ASAP7_75t_L g303 ( .A(n_120), .B(n_249), .Y(n_303) );
AND2x2_ASAP7_75t_L g311 ( .A(n_120), .B(n_254), .Y(n_311) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g241 ( .A(n_121), .B(n_149), .Y(n_241) );
INVx2_ASAP7_75t_L g253 ( .A(n_121), .Y(n_253) );
AND2x2_ASAP7_75t_L g378 ( .A(n_121), .B(n_320), .Y(n_378) );
OR2x2_ASAP7_75t_L g380 ( .A(n_121), .B(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_128), .Y(n_121) );
INVx1_ASAP7_75t_L g247 ( .A(n_122), .Y(n_247) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
INVx1_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_124), .B(n_125), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
NAND3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_142), .C(n_144), .Y(n_128) );
AO21x1_ASAP7_75t_L g246 ( .A1(n_129), .A2(n_142), .B(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_132), .B1(n_136), .B2(n_139), .Y(n_129) );
INVx2_ASAP7_75t_L g193 ( .A(n_130), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_130), .A2(n_138), .B1(n_198), .B2(n_200), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_130), .A2(n_136), .B1(n_205), .B2(n_206), .Y(n_204) );
INVx4_ASAP7_75t_L g484 ( .A(n_130), .Y(n_484) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx3_ASAP7_75t_L g138 ( .A(n_131), .Y(n_138) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
INVx1_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
AND2x2_ASAP7_75t_L g462 ( .A(n_131), .B(n_159), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_131), .Y(n_465) );
INVx2_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_136), .A2(n_156), .B(n_157), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_136), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_137), .A2(n_153), .B(n_154), .Y(n_152) );
O2A1O1Ixp5_ASAP7_75t_SL g212 ( .A1(n_137), .A2(n_213), .B(n_214), .C(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_137), .A2(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_137), .B(n_512), .Y(n_511) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_140), .Y(n_560) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
BUFx3_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
AND2x6_ASAP7_75t_L g464 ( .A(n_141), .B(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g476 ( .A(n_142), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_142), .B(n_503), .Y(n_502) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_142), .A2(n_528), .B(n_535), .Y(n_527) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_142), .A2(n_555), .B(n_562), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_142), .B(n_563), .Y(n_562) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_143), .A2(n_151), .B(n_160), .Y(n_150) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_143), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_143), .A2(n_540), .B(n_541), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_144), .A2(n_234), .B(n_237), .Y(n_233) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g151 ( .A1(n_145), .A2(n_152), .B(n_155), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_145), .A2(n_165), .B(n_172), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_145), .A2(n_184), .B(n_189), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_145), .A2(n_212), .B(n_216), .Y(n_211) );
AND2x4_ASAP7_75t_L g461 ( .A(n_145), .B(n_462), .Y(n_461) );
INVx4_ASAP7_75t_SL g486 ( .A(n_145), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_145), .B(n_462), .Y(n_530) );
INVx2_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g291 ( .A(n_148), .B(n_263), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_148), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g405 ( .A(n_148), .B(n_245), .Y(n_405) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_161), .Y(n_148) );
AND2x2_ASAP7_75t_L g248 ( .A(n_149), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g295 ( .A(n_149), .Y(n_295) );
AND2x2_ASAP7_75t_L g320 ( .A(n_149), .B(n_232), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_149), .B(n_353), .Y(n_390) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g254 ( .A(n_150), .B(n_232), .Y(n_254) );
AND2x2_ASAP7_75t_L g268 ( .A(n_150), .B(n_231), .Y(n_268) );
AND2x2_ASAP7_75t_L g285 ( .A(n_150), .B(n_161), .Y(n_285) );
AND2x2_ASAP7_75t_L g342 ( .A(n_150), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_150), .B(n_249), .Y(n_355) );
AND2x2_ASAP7_75t_L g407 ( .A(n_150), .B(n_332), .Y(n_407) );
INVx2_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g230 ( .A(n_161), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g249 ( .A(n_161), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_161), .B(n_232), .Y(n_326) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_176), .Y(n_161) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_162), .A2(n_233), .B(n_240), .Y(n_232) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_163), .B(n_536), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_169), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_167), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_167), .A2(n_543), .B(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_169), .A2(n_558), .B(n_559), .C(n_560), .Y(n_557) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_170), .A2(n_217), .B(n_218), .Y(n_216) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g468 ( .A(n_171), .Y(n_468) );
O2A1O1Ixp5_ASAP7_75t_L g237 ( .A1(n_173), .A2(n_193), .B(n_238), .C(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_173), .A2(n_467), .B(n_469), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_207), .B(n_220), .Y(n_177) );
INVx1_ASAP7_75t_SL g339 ( .A(n_178), .Y(n_339) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_195), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_SL g227 ( .A(n_180), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g222 ( .A(n_181), .Y(n_222) );
INVx1_ASAP7_75t_L g259 ( .A(n_181), .Y(n_259) );
AND2x2_ASAP7_75t_L g280 ( .A(n_181), .B(n_202), .Y(n_280) );
AND2x2_ASAP7_75t_L g314 ( .A(n_181), .B(n_203), .Y(n_314) );
OR2x2_ASAP7_75t_L g333 ( .A(n_181), .B(n_209), .Y(n_333) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_181), .Y(n_347) );
AND2x2_ASAP7_75t_L g360 ( .A(n_181), .B(n_361), .Y(n_360) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_194), .Y(n_181) );
INVx2_ASAP7_75t_L g201 ( .A(n_182), .Y(n_201) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_182), .A2(n_211), .B(n_219), .Y(n_210) );
INVx1_ASAP7_75t_L g474 ( .A(n_182), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_182), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_182), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_193), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_195), .A2(n_282), .B1(n_283), .B2(n_292), .Y(n_281) );
AND2x2_ASAP7_75t_L g365 ( .A(n_195), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_202), .Y(n_195) );
INVx1_ASAP7_75t_L g226 ( .A(n_196), .Y(n_226) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
INVx1_ASAP7_75t_L g274 ( .A(n_196), .Y(n_274) );
AND2x2_ASAP7_75t_L g289 ( .A(n_196), .B(n_203), .Y(n_289) );
INVx2_ASAP7_75t_L g485 ( .A(n_199), .Y(n_485) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_199), .Y(n_500) );
INVx1_ASAP7_75t_L g471 ( .A(n_201), .Y(n_471) );
OR2x2_ASAP7_75t_L g243 ( .A(n_202), .B(n_228), .Y(n_243) );
AND2x2_ASAP7_75t_L g273 ( .A(n_202), .B(n_274), .Y(n_273) );
NOR2xp67_ASAP7_75t_L g361 ( .A(n_202), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g221 ( .A(n_203), .B(n_222), .Y(n_221) );
BUFx2_ASAP7_75t_L g330 ( .A(n_203), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_207), .B(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g308 ( .A(n_208), .B(n_274), .Y(n_308) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g220 ( .A(n_209), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
OR2x2_ASAP7_75t_L g258 ( .A(n_210), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_210), .Y(n_313) );
AOI32xp33_ASAP7_75t_L g350 ( .A1(n_220), .A2(n_280), .A3(n_351), .B1(n_352), .B2(n_354), .Y(n_350) );
AND2x2_ASAP7_75t_L g276 ( .A(n_221), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_221), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_221), .B(n_308), .Y(n_394) );
INVx1_ASAP7_75t_L g399 ( .A(n_221), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_229), .B1(n_242), .B2(n_244), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
AND2x2_ASAP7_75t_L g329 ( .A(n_225), .B(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_226), .B(n_228), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_251), .B1(n_255), .B2(n_265), .Y(n_250) );
AND2x2_ASAP7_75t_L g272 ( .A(n_227), .B(n_273), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_227), .A2(n_241), .B(n_289), .C(n_324), .Y(n_323) );
OAI332xp33_ASAP7_75t_L g328 ( .A1(n_227), .A2(n_329), .A3(n_331), .B1(n_333), .B2(n_334), .B3(n_336), .C1(n_337), .C2(n_339), .Y(n_328) );
INVx2_ASAP7_75t_L g369 ( .A(n_227), .Y(n_369) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_228), .Y(n_287) );
INVx1_ASAP7_75t_L g362 ( .A(n_228), .Y(n_362) );
AND2x2_ASAP7_75t_L g416 ( .A(n_228), .B(n_280), .Y(n_416) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_241), .Y(n_229) );
AND2x2_ASAP7_75t_L g296 ( .A(n_231), .B(n_246), .Y(n_296) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g245 ( .A(n_232), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g344 ( .A(n_232), .B(n_246), .Y(n_344) );
INVx1_ASAP7_75t_L g353 ( .A(n_232), .Y(n_353) );
INVx1_ASAP7_75t_L g327 ( .A(n_241), .Y(n_327) );
INVxp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g411 ( .A(n_243), .B(n_263), .Y(n_411) );
INVx1_ASAP7_75t_SL g322 ( .A(n_244), .Y(n_322) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
AND2x2_ASAP7_75t_L g349 ( .A(n_245), .B(n_307), .Y(n_349) );
INVx1_ASAP7_75t_L g368 ( .A(n_245), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_245), .B(n_335), .Y(n_370) );
INVx1_ASAP7_75t_L g267 ( .A(n_246), .Y(n_267) );
AND2x2_ASAP7_75t_L g271 ( .A(n_248), .B(n_252), .Y(n_271) );
AND2x2_ASAP7_75t_L g338 ( .A(n_248), .B(n_296), .Y(n_338) );
INVx2_ASAP7_75t_L g381 ( .A(n_248), .Y(n_381) );
INVx2_ASAP7_75t_L g264 ( .A(n_249), .Y(n_264) );
AND2x2_ASAP7_75t_L g266 ( .A(n_249), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g282 ( .A(n_252), .Y(n_282) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_253), .B(n_326), .Y(n_332) );
OR2x2_ASAP7_75t_L g396 ( .A(n_253), .B(n_355), .Y(n_396) );
INVx1_ASAP7_75t_L g420 ( .A(n_253), .Y(n_420) );
INVx1_ASAP7_75t_L g376 ( .A(n_254), .Y(n_376) );
AND2x2_ASAP7_75t_L g421 ( .A(n_254), .B(n_264), .Y(n_421) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_284), .B1(n_286), .B2(n_290), .Y(n_283) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI322xp33_ASAP7_75t_SL g367 ( .A1(n_261), .A2(n_368), .A3(n_369), .B1(n_370), .B2(n_371), .C1(n_374), .C2(n_376), .Y(n_367) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g364 ( .A(n_262), .B(n_280), .Y(n_364) );
OR2x2_ASAP7_75t_L g398 ( .A(n_262), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g401 ( .A(n_262), .B(n_333), .Y(n_401) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g346 ( .A(n_263), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g402 ( .A(n_263), .B(n_333), .Y(n_402) );
INVx3_ASAP7_75t_L g335 ( .A(n_264), .Y(n_335) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g391 ( .A(n_266), .Y(n_391) );
AOI222xp33_ASAP7_75t_L g270 ( .A1(n_268), .A2(n_271), .B1(n_272), .B2(n_275), .C1(n_276), .C2(n_278), .Y(n_270) );
INVx1_ASAP7_75t_L g301 ( .A(n_268), .Y(n_301) );
NAND3xp33_ASAP7_75t_SL g269 ( .A(n_270), .B(n_281), .C(n_298), .Y(n_269) );
AND2x2_ASAP7_75t_L g386 ( .A(n_273), .B(n_287), .Y(n_386) );
BUFx2_ASAP7_75t_L g277 ( .A(n_274), .Y(n_277) );
INVx1_ASAP7_75t_L g318 ( .A(n_274), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_275), .A2(n_311), .B1(n_364), .B2(n_365), .C(n_367), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_277), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_280), .Y(n_304) );
AND2x2_ASAP7_75t_L g317 ( .A(n_280), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_285), .B(n_296), .Y(n_297) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
OAI21xp33_ASAP7_75t_L g292 ( .A1(n_287), .A2(n_293), .B(n_297), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_287), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g384 ( .A(n_289), .B(n_366), .Y(n_384) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g307 ( .A(n_295), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_296), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g413 ( .A(n_296), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_304), .B1(n_305), .B2(n_308), .C(n_309), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_300), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g409 ( .A(n_308), .B(n_314), .Y(n_409) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
OAI31xp33_ASAP7_75t_SL g377 ( .A1(n_312), .A2(n_351), .A3(n_378), .B(n_379), .Y(n_377) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g366 ( .A(n_313), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_314), .B(n_318), .Y(n_417) );
OAI221xp5_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_319), .B1(n_321), .B2(n_322), .C(n_323), .Y(n_315) );
INVx1_ASAP7_75t_L g321 ( .A(n_317), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_320), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g336 ( .A(n_329), .Y(n_336) );
INVx2_ASAP7_75t_L g372 ( .A(n_330), .Y(n_372) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g358 ( .A(n_335), .B(n_344), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_335), .A2(n_352), .B(n_409), .C(n_410), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g340 ( .A1(n_336), .A2(n_341), .B1(n_345), .B2(n_348), .C(n_350), .Y(n_340) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_339), .A2(n_404), .B(n_406), .C(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_342), .A2(n_393), .B1(n_395), .B2(n_397), .C(n_400), .Y(n_392) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
NOR4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_382), .C(n_403), .D(n_414), .Y(n_356) );
OAI211xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_359), .B(n_363), .C(n_377), .Y(n_357) );
INVx1_ASAP7_75t_SL g412 ( .A(n_364), .Y(n_412) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_SL g375 ( .A(n_373), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_380), .A2(n_389), .B1(n_401), .B2(n_402), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B(n_387), .C(n_392), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI31xp33_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_415), .A3(n_417), .B(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g433 ( .A(n_426), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_426), .B(n_435), .Y(n_434) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_427), .B(n_736), .Y(n_742) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g735 ( .A(n_428), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
NAND3xp33_ASAP7_75t_SL g750 ( .A(n_429), .B(n_736), .C(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_434), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g737 ( .A(n_439), .Y(n_737) );
INVx1_ASAP7_75t_L g443 ( .A(n_440), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_448), .B1(n_451), .B2(n_733), .Y(n_445) );
INVx1_ASAP7_75t_L g739 ( .A(n_446), .Y(n_739) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_450), .A2(n_452), .B1(n_735), .B2(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_453), .B(n_669), .Y(n_452) );
NOR5xp2_ASAP7_75t_L g453 ( .A(n_454), .B(n_600), .C(n_629), .D(n_649), .E(n_656), .Y(n_453) );
OAI211xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_488), .B(n_545), .C(n_587), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_456), .A2(n_672), .B1(n_674), .B2(n_675), .Y(n_671) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_475), .Y(n_456) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_457), .Y(n_548) );
AND2x4_ASAP7_75t_L g580 ( .A(n_457), .B(n_581), .Y(n_580) );
INVx5_ASAP7_75t_L g598 ( .A(n_457), .Y(n_598) );
AND2x2_ASAP7_75t_L g607 ( .A(n_457), .B(n_599), .Y(n_607) );
AND2x2_ASAP7_75t_L g619 ( .A(n_457), .B(n_492), .Y(n_619) );
AND2x2_ASAP7_75t_L g715 ( .A(n_457), .B(n_583), .Y(n_715) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_472), .Y(n_457) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_463), .B(n_471), .Y(n_458) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx5_ASAP7_75t_L g480 ( .A(n_464), .Y(n_480) );
INVx2_ASAP7_75t_L g470 ( .A(n_468), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_470), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_470), .A2(n_500), .B(n_522), .C(n_523), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g581 ( .A(n_475), .Y(n_581) );
AND2x2_ASAP7_75t_L g599 ( .A(n_475), .B(n_554), .Y(n_599) );
AND2x2_ASAP7_75t_L g618 ( .A(n_475), .B(n_553), .Y(n_618) );
AND2x2_ASAP7_75t_L g658 ( .A(n_475), .B(n_598), .Y(n_658) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_487), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .B(n_481), .C(n_486), .Y(n_478) );
INVx2_ASAP7_75t_L g496 ( .A(n_480), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_480), .A2(n_486), .B(n_509), .C(n_510), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g501 ( .A(n_486), .Y(n_501) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_514), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI322xp5_ASAP7_75t_L g717 ( .A1(n_491), .A2(n_525), .A3(n_572), .B1(n_580), .B2(n_634), .C1(n_718), .C2(n_721), .Y(n_717) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_504), .Y(n_491) );
INVx5_ASAP7_75t_L g550 ( .A(n_492), .Y(n_550) );
AND2x2_ASAP7_75t_L g566 ( .A(n_492), .B(n_552), .Y(n_566) );
BUFx2_ASAP7_75t_L g644 ( .A(n_492), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_492), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g721 ( .A(n_492), .B(n_628), .Y(n_721) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_504), .B(n_516), .Y(n_575) );
INVx1_ASAP7_75t_L g602 ( .A(n_504), .Y(n_602) );
AND2x2_ASAP7_75t_L g615 ( .A(n_504), .B(n_537), .Y(n_615) );
AND2x2_ASAP7_75t_L g716 ( .A(n_504), .B(n_634), .Y(n_716) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g570 ( .A(n_505), .B(n_516), .Y(n_570) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_505), .Y(n_578) );
OR2x2_ASAP7_75t_L g585 ( .A(n_505), .B(n_537), .Y(n_585) );
AND2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_505), .B(n_527), .Y(n_624) );
INVxp67_ASAP7_75t_L g648 ( .A(n_505), .Y(n_648) );
AND2x2_ASAP7_75t_L g655 ( .A(n_505), .B(n_525), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_505), .B(n_537), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_505), .B(n_526), .Y(n_681) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_513), .Y(n_505) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_516), .B(n_538), .Y(n_625) );
OR2x2_ASAP7_75t_L g647 ( .A(n_516), .B(n_526), .Y(n_647) );
AND2x2_ASAP7_75t_L g660 ( .A(n_516), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_516), .B(n_615), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_516), .A2(n_671), .B(n_676), .C(n_685), .Y(n_670) );
AND2x2_ASAP7_75t_L g731 ( .A(n_516), .B(n_537), .Y(n_731) );
INVx5_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g584 ( .A(n_517), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_517), .B(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_517), .B(n_579), .Y(n_591) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_517), .Y(n_593) );
OR2x2_ASAP7_75t_L g604 ( .A(n_517), .B(n_526), .Y(n_604) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_517), .B(n_595), .Y(n_609) );
AND2x2_ASAP7_75t_L g634 ( .A(n_517), .B(n_526), .Y(n_634) );
AND2x2_ASAP7_75t_L g654 ( .A(n_517), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g692 ( .A(n_517), .B(n_525), .Y(n_692) );
OR2x2_ASAP7_75t_L g695 ( .A(n_517), .B(n_681), .Y(n_695) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_526), .A2(n_639), .B(n_642), .C(n_648), .Y(n_638) );
INVx5_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_527), .B(n_537), .Y(n_569) );
AND2x2_ASAP7_75t_L g573 ( .A(n_527), .B(n_538), .Y(n_573) );
OR2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_537), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_SL g596 ( .A(n_537), .Y(n_596) );
OR2x2_ASAP7_75t_L g724 ( .A(n_537), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_564), .B(n_567), .C(n_576), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI31xp33_ASAP7_75t_L g649 ( .A1(n_547), .A2(n_650), .A3(n_652), .B(n_653), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_548), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_549), .B(n_580), .Y(n_586) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_550), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g606 ( .A(n_550), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_550), .B(n_581), .Y(n_611) );
AND2x2_ASAP7_75t_L g621 ( .A(n_550), .B(n_580), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_550), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g641 ( .A(n_550), .B(n_598), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_550), .B(n_618), .Y(n_646) );
OR2x2_ASAP7_75t_L g665 ( .A(n_550), .B(n_552), .Y(n_665) );
OR2x2_ASAP7_75t_L g667 ( .A(n_550), .B(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_550), .Y(n_714) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g614 ( .A(n_552), .B(n_581), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_552), .B(n_598), .Y(n_637) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g583 ( .A(n_554), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g674 ( .A(n_566), .B(n_598), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_566), .A2(n_580), .A3(n_618), .B1(n_677), .B2(n_678), .C1(n_679), .C2(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g684 ( .A(n_566), .Y(n_684) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_SL g678 ( .A(n_568), .Y(n_678) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
OR2x2_ASAP7_75t_L g630 ( .A(n_569), .B(n_575), .Y(n_630) );
INVx1_ASAP7_75t_L g661 ( .A(n_569), .Y(n_661) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI32xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .A3(n_582), .B1(n_584), .B2(n_586), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI21xp33_ASAP7_75t_SL g616 ( .A1(n_579), .A2(n_594), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g631 ( .A(n_580), .Y(n_631) );
AND2x4_ASAP7_75t_L g628 ( .A(n_581), .B(n_598), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_581), .B(n_664), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_582), .A2(n_609), .A3(n_628), .B1(n_661), .B2(n_694), .C1(n_696), .C2(n_697), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_582), .A2(n_659), .B1(n_723), .B2(n_724), .C(n_726), .Y(n_722) );
AND2x2_ASAP7_75t_L g610 ( .A(n_583), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g590 ( .A(n_585), .Y(n_590) );
OR2x2_ASAP7_75t_L g662 ( .A(n_585), .B(n_647), .Y(n_662) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .A3(n_592), .B(n_597), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_588), .A2(n_621), .B1(n_622), .B2(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g633 ( .A(n_590), .B(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_592), .A2(n_633), .B1(n_686), .B2(n_689), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g675 ( .A(n_595), .B(n_644), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_595), .B(n_634), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_596), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g709 ( .A(n_596), .B(n_647), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_597), .A2(n_692), .B1(n_705), .B2(n_708), .Y(n_704) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g613 ( .A(n_598), .Y(n_613) );
AND2x2_ASAP7_75t_L g696 ( .A(n_598), .B(n_618), .Y(n_696) );
OR2x2_ASAP7_75t_L g698 ( .A(n_598), .B(n_665), .Y(n_698) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_598), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_599), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_599), .B(n_644), .Y(n_652) );
OAI211xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_605), .B(n_608), .C(n_620), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_612), .B2(n_615), .C(n_616), .Y(n_608) );
INVxp67_ASAP7_75t_L g720 ( .A(n_611), .Y(n_720) );
INVx1_ASAP7_75t_L g687 ( .A(n_612), .Y(n_687) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g651 ( .A(n_613), .B(n_618), .Y(n_651) );
INVx1_ASAP7_75t_L g668 ( .A(n_614), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_614), .B(n_641), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g683 ( .A(n_618), .Y(n_683) );
AND2x2_ASAP7_75t_L g689 ( .A(n_618), .B(n_644), .Y(n_689) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_SL g677 ( .A(n_625), .Y(n_677) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_628), .B(n_664), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_635), .C(n_638), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g725 ( .A(n_634), .Y(n_725) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g643 ( .A(n_637), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_641), .B(n_700), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_647), .Y(n_642) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_645), .A2(n_691), .B(n_693), .C(n_699), .Y(n_690) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g702 ( .A(n_647), .Y(n_702) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI222xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B1(n_662), .B2(n_663), .C1(n_666), .C2(n_667), .Y(n_656) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g732 ( .A(n_663), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_664), .B(n_707), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_664), .A2(n_711), .B1(n_713), .B2(n_716), .Y(n_710) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NOR4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_690), .C(n_703), .D(n_722), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_672), .B(n_702), .Y(n_712) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g679 ( .A(n_677), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_680), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_710), .C(n_717), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx2_ASAP7_75t_L g719 ( .A(n_715), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_729), .B(n_732), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_SL g756 ( .A(n_745), .Y(n_756) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx14_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
endmodule