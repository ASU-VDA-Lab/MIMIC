module fake_netlist_6_3999_n_87 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_87);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_87;

wire n_52;
wire n_46;
wire n_21;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_86;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_19),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_7),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_2),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_23),
.B(n_24),
.Y(n_41)
);

AO21x2_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_24),
.B(n_20),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_27),
.B(n_25),
.C(n_34),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_40),
.B(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI211xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_28),
.B(n_38),
.C(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AO21x2_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_20),
.B(n_27),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_42),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_46),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_42),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_46),
.Y(n_57)
);

AND2x4_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_25),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

AOI221x1_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_33),
.B1(n_21),
.B2(n_29),
.C(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_53),
.B(n_51),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_53),
.Y(n_64)
);

OAI31xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_51),
.A3(n_21),
.B(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_56),
.Y(n_66)
);

O2A1O1Ixp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_59),
.B(n_50),
.C(n_47),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_34),
.A3(n_31),
.B1(n_30),
.B2(n_6),
.C1(n_13),
.C2(n_11),
.Y(n_68)
);

AOI221xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_34),
.B1(n_31),
.B2(n_58),
.C(n_53),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_62),
.B1(n_66),
.B2(n_60),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_50),
.C(n_47),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_50),
.B(n_47),
.C(n_49),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_53),
.B1(n_49),
.B2(n_47),
.Y(n_73)
);

AOI211xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_65),
.B(n_63),
.C(n_30),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_61),
.C(n_49),
.Y(n_75)
);

OAI221xp5_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_60),
.B1(n_66),
.B2(n_53),
.C(n_6),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_60),
.B1(n_13),
.B2(n_11),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_49),
.Y(n_78)
);

AND4x1_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_30),
.C(n_15),
.D(n_49),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_30),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_67),
.C(n_30),
.Y(n_82)
);

XOR2x1_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_77),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_75),
.Y(n_84)
);

AOI222xp33_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_74),
.B1(n_78),
.B2(n_81),
.C1(n_82),
.C2(n_83),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2x2_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_85),
.Y(n_87)
);


endmodule