module real_jpeg_23262_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_59),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_1),
.A2(n_59),
.B1(n_65),
.B2(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_2),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_5),
.A2(n_47),
.B1(n_65),
.B2(n_66),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_5),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_71),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_7),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_7),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_10),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_10),
.B(n_66),
.C(n_88),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_10),
.B(n_60),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_103),
.B1(n_172),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_99),
.Y(n_209)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_13),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_94),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_94),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_77),
.Y(n_124)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_137),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_19),
.B(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_101),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_20),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_61),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_44),
.C(n_82),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_38),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_25),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_25),
.A2(n_41),
.B1(n_99),
.B2(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_27),
.A2(n_30),
.B(n_79),
.C(n_81),
.Y(n_78)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_32),
.C(n_35),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_29),
.B(n_51),
.C(n_55),
.Y(n_188)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g187 ( 
.A(n_30),
.B(n_80),
.CON(n_187),
.SN(n_187)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_35),
.B(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_37),
.A2(n_79),
.B(n_80),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_38),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_57),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_49),
.B1(n_60),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_48),
.A2(n_53),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_49),
.A2(n_58),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_49),
.A2(n_60),
.B1(n_187),
.B2(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_52),
.A2(n_54),
.B(n_186),
.C(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_53),
.B(n_133),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_55),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_55),
.B(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_78),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_62),
.A2(n_63),
.B1(n_78),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_76),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_117),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_66),
.B1(n_88),
.B2(n_89),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_65),
.B(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_68),
.B(n_80),
.Y(n_177)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_68),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_70),
.A2(n_120),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_73),
.A2(n_103),
.B1(n_165),
.B2(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_75),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_78),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_80),
.B(n_90),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_83),
.B(n_101),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.C(n_97),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_84),
.B(n_95),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_91),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_85),
.A2(n_123),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_85),
.A2(n_123),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_86),
.A2(n_90),
.B1(n_151),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_86),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_91),
.B(n_123),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_96),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_97),
.B(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_116),
.B(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_103),
.A2(n_105),
.B(n_119),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_134),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_126),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_121),
.B2(n_125),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_237),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_233),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_223),
.B(n_232),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_199),
.B(n_222),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_181),
.B(n_198),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_161),
.B(n_180),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_152),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_148),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_156),
.C(n_159),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_168),
.B(n_179),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_167),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_173),
.B(n_178),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_197),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_197),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_192),
.C(n_194),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_196),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_201),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_214),
.B2(n_215),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_217),
.C(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_208),
.C(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_231),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_228),
.C(n_229),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);


endmodule