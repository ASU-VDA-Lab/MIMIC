module fake_jpeg_5895_n_299 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_15),
.B(n_21),
.Y(n_49)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_39),
.Y(n_59)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_35),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_61),
.B1(n_26),
.B2(n_35),
.Y(n_72)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_23),
.B1(n_16),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_39),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_32),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_23),
.B1(n_16),
.B2(n_19),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_19),
.B1(n_23),
.B2(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_39),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_39),
.B1(n_36),
.B2(n_28),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_72),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_32),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_59),
.C(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_35),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_39),
.B1(n_34),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_73),
.B1(n_79),
.B2(n_46),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_71),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_39),
.B1(n_34),
.B2(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_40),
.B(n_38),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_83),
.B(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_32),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_82),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_31),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_105),
.B(n_80),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_93),
.Y(n_125)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_90),
.Y(n_124)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_46),
.B1(n_52),
.B2(n_44),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_100),
.B1(n_73),
.B2(n_50),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_59),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_61),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_83),
.C(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_57),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_104),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_30),
.B(n_43),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_68),
.B(n_62),
.C(n_82),
.D(n_64),
.Y(n_122)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx11_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_115),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_81),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_68),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_122),
.B(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_83),
.B1(n_72),
.B2(n_80),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_131),
.B1(n_77),
.B2(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_108),
.Y(n_143)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_72),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_54),
.B1(n_78),
.B2(n_76),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_45),
.B1(n_51),
.B2(n_48),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_92),
.B1(n_86),
.B2(n_91),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_88),
.C(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_148),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_58),
.B(n_75),
.C(n_124),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_144),
.B1(n_146),
.B2(n_150),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_86),
.B(n_91),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_141),
.B(n_142),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_92),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_92),
.B(n_108),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_153),
.B(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_92),
.B1(n_76),
.B2(n_66),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_66),
.B1(n_69),
.B2(n_77),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_85),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_77),
.B1(n_52),
.B2(n_44),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_151),
.B(n_60),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_38),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_84),
.B(n_104),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_52),
.B1(n_60),
.B2(n_31),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_104),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_38),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_30),
.A3(n_17),
.B1(n_58),
.B2(n_18),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_158),
.B(n_126),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_165),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_119),
.B1(n_109),
.B2(n_115),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_162),
.B1(n_169),
.B2(n_177),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_123),
.B1(n_131),
.B2(n_116),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_167),
.B1(n_171),
.B2(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_112),
.B1(n_132),
.B2(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_112),
.B1(n_89),
.B2(n_128),
.Y(n_171)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_152),
.B1(n_143),
.B2(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_26),
.B1(n_18),
.B2(n_24),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_178),
.A2(n_184),
.B1(n_70),
.B2(n_24),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_99),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_183),
.B1(n_21),
.B2(n_15),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_99),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_173),
.B1(n_161),
.B2(n_174),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_189),
.A2(n_194),
.B1(n_206),
.B2(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_141),
.C(n_136),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_193),
.C(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_145),
.C(n_148),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_138),
.B1(n_150),
.B2(n_156),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_140),
.B1(n_139),
.B2(n_149),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_164),
.B1(n_21),
.B2(n_15),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_158),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_197),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_29),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_22),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_203),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_204),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_22),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_111),
.C(n_94),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_111),
.B1(n_70),
.B2(n_94),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_220),
.B1(n_202),
.B2(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_226),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_171),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_177),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_197),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_165),
.B1(n_180),
.B2(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_222),
.B1(n_24),
.B2(n_21),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_175),
.B1(n_164),
.B2(n_159),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_111),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_198),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_227),
.C(n_194),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_13),
.B(n_12),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_29),
.C(n_22),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_0),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_245),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_239),
.B(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_187),
.CI(n_199),
.CON(n_235),
.SN(n_235)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_242),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_29),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_216),
.C(n_213),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_238),
.C(n_29),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_213),
.C(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_199),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_222),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_1),
.B(n_2),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_210),
.B1(n_224),
.B2(n_211),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_15),
.B1(n_24),
.B2(n_22),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_214),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_242),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_255),
.C(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_244),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_11),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_1),
.C(n_2),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_13),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_259),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_240),
.B(n_235),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_231),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_3),
.C(n_4),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_12),
.Y(n_259)
);

AND2x4_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_3),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_6),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_267),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_234),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_251),
.A2(n_229),
.B1(n_11),
.B2(n_5),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_274),
.B1(n_5),
.B2(n_6),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_260),
.B1(n_261),
.B2(n_257),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_270),
.B1(n_271),
.B2(n_262),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_3),
.B(n_4),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_4),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_255),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_280),
.B(n_282),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_250),
.C(n_258),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_9),
.C(n_7),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_4),
.B(n_5),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_284),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_287),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_275),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_288),
.A2(n_290),
.B(n_285),
.Y(n_295)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_269),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_289),
.B(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_278),
.C(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_294),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_295),
.C(n_297),
.Y(n_299)
);


endmodule