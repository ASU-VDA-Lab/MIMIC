module fake_jpeg_12569_n_390 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_57),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_83),
.Y(n_127)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_89),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_6),
.CON(n_70),
.SN(n_70)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_109),
.Y(n_117)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_74),
.B(n_82),
.Y(n_168)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_7),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_23),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_100),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_54),
.B1(n_49),
.B2(n_27),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_54),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_14),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_96),
.B(n_105),
.Y(n_170)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_98),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_103),
.Y(n_130)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_106),
.Y(n_121)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_107),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_20),
.B(n_14),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_111),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_35),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_110),
.Y(n_124)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_44),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_113),
.A2(n_123),
.B1(n_129),
.B2(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_146),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_94),
.B1(n_107),
.B2(n_99),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_41),
.B1(n_45),
.B2(n_27),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_128),
.A2(n_123),
.B1(n_133),
.B2(n_174),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_28),
.B1(n_55),
.B2(n_26),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_131),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_28),
.B1(n_44),
.B2(n_52),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_138),
.B(n_140),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_59),
.B(n_55),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_52),
.B1(n_50),
.B2(n_39),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_147),
.B1(n_149),
.B2(n_153),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_105),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_61),
.A2(n_50),
.B1(n_39),
.B2(n_32),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_66),
.A2(n_31),
.B1(n_32),
.B2(n_41),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_72),
.A2(n_31),
.B1(n_45),
.B2(n_3),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_74),
.B(n_3),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_161),
.B(n_163),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_96),
.B(n_3),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_84),
.B(n_3),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_164),
.B(n_166),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_48),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_86),
.A2(n_48),
.B1(n_87),
.B2(n_88),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_176),
.B1(n_157),
.B2(n_158),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_91),
.B(n_48),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_98),
.B(n_48),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_62),
.A2(n_100),
.B1(n_93),
.B2(n_58),
.Y(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_147),
.B1(n_128),
.B2(n_145),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_183),
.A2(n_201),
.B1(n_215),
.B2(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_119),
.A2(n_125),
.B1(n_159),
.B2(n_151),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_187),
.A2(n_192),
.B1(n_226),
.B2(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_124),
.B(n_144),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_191),
.B(n_216),
.C(n_219),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_119),
.A2(n_169),
.B1(n_115),
.B2(n_168),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_206),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_198),
.A2(n_211),
.B1(n_213),
.B2(n_217),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_152),
.B(n_135),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_200),
.B(n_204),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_127),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_224),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_134),
.B1(n_128),
.B2(n_129),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_135),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_207),
.Y(n_246)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

BUFx24_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_218),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_130),
.B1(n_175),
.B2(n_165),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_165),
.A2(n_133),
.B1(n_174),
.B2(n_143),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_217),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_118),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_116),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_139),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_150),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_114),
.A2(n_117),
.B1(n_139),
.B2(n_156),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_150),
.B(n_156),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_221),
.B(n_222),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_150),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_167),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_144),
.A2(n_113),
.B1(n_124),
.B2(n_153),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_223),
.A3(n_227),
.B1(n_191),
.B2(n_182),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_232),
.A2(n_259),
.B(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_240),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_216),
.Y(n_240)
);

XOR2x1_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_216),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_179),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_257),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_242),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_198),
.A2(n_186),
.B1(n_190),
.B2(n_228),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_252),
.A2(n_258),
.B1(n_261),
.B2(n_267),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_181),
.C(n_180),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_270),
.C(n_264),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_178),
.B(n_218),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_206),
.B1(n_195),
.B2(n_196),
.Y(n_258)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_219),
.A2(n_177),
.A3(n_210),
.B1(n_224),
.B2(n_212),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_185),
.A2(n_194),
.B1(n_208),
.B2(n_214),
.Y(n_261)
);

AO22x2_ASAP7_75t_L g269 ( 
.A1(n_193),
.A2(n_183),
.B1(n_186),
.B2(n_201),
.Y(n_269)
);

AO21x2_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_241),
.B(n_238),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_193),
.B(n_144),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_244),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_186),
.A2(n_179),
.B(n_201),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_249),
.B1(n_269),
.B2(n_272),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_273),
.A2(n_297),
.B1(n_276),
.B2(n_287),
.Y(n_318)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_260),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_283),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_256),
.B1(n_298),
.B2(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_277),
.B(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_235),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_280),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_240),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_237),
.B(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_282),
.B(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_239),
.Y(n_284)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_295),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_289),
.A2(n_297),
.B(n_300),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_245),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_290),
.B(n_293),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_255),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_270),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_269),
.B(n_270),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_247),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_298),
.B(n_299),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_234),
.B(n_268),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_254),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_255),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_233),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_290),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_295),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_266),
.C(n_261),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_308),
.C(n_317),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_297),
.B(n_296),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_256),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_312),
.A2(n_317),
.B(n_276),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_281),
.B(n_300),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_314),
.A2(n_301),
.B(n_303),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_285),
.B1(n_281),
.B2(n_278),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_283),
.B1(n_286),
.B2(n_294),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_285),
.A2(n_291),
.B(n_276),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_296),
.B1(n_293),
.B2(n_302),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_280),
.A3(n_279),
.B1(n_297),
.B2(n_292),
.C1(n_274),
.C2(n_288),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_319),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_323),
.A2(n_330),
.B1(n_337),
.B2(n_312),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_275),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_324),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_327),
.A2(n_334),
.B1(n_338),
.B2(n_315),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_306),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_329),
.B(n_332),
.Y(n_341)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_308),
.B(n_316),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_320),
.Y(n_333)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_318),
.A2(n_320),
.B1(n_317),
.B2(n_314),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_307),
.Y(n_335)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_308),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_310),
.A2(n_309),
.B1(n_306),
.B2(n_321),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_311),
.B(n_304),
.Y(n_339)
);

OA21x2_ASAP7_75t_SL g344 ( 
.A1(n_339),
.A2(n_313),
.B(n_322),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_SL g363 ( 
.A(n_342),
.B(n_337),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_344),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_336),
.C(n_332),
.Y(n_355)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_348),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_350),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_323),
.A2(n_318),
.B1(n_312),
.B2(n_305),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_361),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_347),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_359),
.Y(n_367)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_358),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_326),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_346),
.A2(n_325),
.B(n_305),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_360),
.A2(n_362),
.B(n_363),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_345),
.A2(n_325),
.B(n_334),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_350),
.A2(n_328),
.B(n_327),
.Y(n_362)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_353),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_356),
.A2(n_323),
.B1(n_348),
.B2(n_351),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_368),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_356),
.A2(n_324),
.B1(n_340),
.B2(n_330),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_355),
.C(n_354),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_341),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_338),
.Y(n_372)
);

AOI21x1_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_359),
.B(n_352),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_354),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_373),
.B(n_375),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_339),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_333),
.Y(n_381)
);

AOI21x1_ASAP7_75t_SL g378 ( 
.A1(n_374),
.A2(n_371),
.B(n_360),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_378),
.A2(n_382),
.B(n_352),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_372),
.A2(n_369),
.B(n_371),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_381),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_384),
.A2(n_385),
.B(n_365),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_376),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_383),
.A2(n_370),
.B(n_331),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_386),
.A2(n_387),
.B(n_370),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_373),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_366),
.Y(n_390)
);


endmodule