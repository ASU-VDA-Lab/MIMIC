module fake_jpeg_11136_n_387 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_61),
.Y(n_119)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_59),
.Y(n_100)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_16),
.B(n_9),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_67),
.Y(n_120)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_31),
.CON(n_64),
.SN(n_64)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_2),
.B(n_3),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_2),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_27),
.B(n_10),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_76),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_32),
.Y(n_131)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_44),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_72),
.B1(n_57),
.B2(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_85),
.A2(n_101),
.B1(n_68),
.B2(n_65),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_89),
.B(n_127),
.Y(n_173)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_96),
.Y(n_138)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_49),
.Y(n_97)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_51),
.B1(n_53),
.B2(n_80),
.Y(n_101)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_41),
.B1(n_18),
.B2(n_42),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_25),
.B1(n_24),
.B2(n_17),
.Y(n_140)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_41),
.C(n_18),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_25),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_43),
.B1(n_42),
.B2(n_46),
.Y(n_139)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_43),
.B1(n_42),
.B2(n_29),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_129),
.B1(n_43),
.B2(n_33),
.Y(n_157)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

HAxp5_ASAP7_75t_SL g122 ( 
.A(n_81),
.B(n_31),
.CON(n_122),
.SN(n_122)
);

OR2x2_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_37),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_48),
.B(n_44),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_83),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_43),
.B1(n_42),
.B2(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_32),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_132),
.B(n_134),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_143),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_139),
.A2(n_160),
.B1(n_90),
.B2(n_105),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_157),
.B1(n_35),
.B2(n_17),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_29),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_147),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_34),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_144),
.B(n_153),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_155),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_33),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx2_ASAP7_75t_SL g186 ( 
.A(n_148),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_24),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_119),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_26),
.B(n_6),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_85),
.B1(n_101),
.B2(n_118),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_99),
.B(n_39),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_36),
.Y(n_178)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_39),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_94),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_116),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_37),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_110),
.B(n_36),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_35),
.Y(n_194)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_96),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_180),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_178),
.B(n_198),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_167),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_189),
.B1(n_212),
.B2(n_139),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_207),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_196),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_135),
.B(n_122),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_89),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_214),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_204),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_110),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_126),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_137),
.Y(n_208)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_145),
.B1(n_84),
.B2(n_111),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_26),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_154),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_108),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_222),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_160),
.B(n_147),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_219),
.B(n_220),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_205),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_149),
.B(n_161),
.Y(n_225)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_171),
.B1(n_84),
.B2(n_137),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_149),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_233),
.C(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_186),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_187),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_231),
.B(n_243),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_138),
.B1(n_172),
.B2(n_165),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_241),
.B1(n_245),
.B2(n_208),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_138),
.C(n_175),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_136),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_242),
.Y(n_250)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_240),
.B1(n_244),
.B2(n_196),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_177),
.A2(n_203),
.B1(n_206),
.B2(n_183),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_136),
.B1(n_145),
.B2(n_170),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_4),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_188),
.B(n_201),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_88),
.B1(n_102),
.B2(n_95),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_176),
.A2(n_150),
.B(n_74),
.C(n_4),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_195),
.A2(n_150),
.B(n_7),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_246),
.B(n_6),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_218),
.A2(n_195),
.B1(n_180),
.B2(n_184),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_248),
.A2(n_266),
.B1(n_251),
.B2(n_247),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_223),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_184),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_268),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_232),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_241),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_214),
.C(n_195),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_273),
.C(n_219),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_226),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_224),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_221),
.B(n_178),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_271),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_221),
.B1(n_225),
.B2(n_222),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_187),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_274),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_197),
.C(n_192),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_215),
.B(n_209),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_298),
.C(n_197),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_228),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_281),
.C(n_285),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_228),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_283),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_233),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_280),
.B(n_289),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_231),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_239),
.B(n_244),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_249),
.B1(n_270),
.B2(n_267),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_266),
.A2(n_226),
.B1(n_217),
.B2(n_235),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_251),
.B1(n_265),
.B2(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_271),
.C(n_256),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_263),
.C(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_217),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_270),
.B1(n_275),
.B2(n_258),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_302),
.A2(n_208),
.B1(n_245),
.B2(n_237),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_282),
.A2(n_290),
.B(n_297),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_309),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_306),
.C(n_310),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_250),
.C(n_272),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_307),
.A2(n_284),
.B1(n_257),
.B2(n_245),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_250),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_254),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_283),
.A2(n_249),
.B1(n_268),
.B2(n_254),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_286),
.B1(n_292),
.B2(n_294),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_299),
.B1(n_294),
.B2(n_279),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_278),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_192),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_318),
.C(n_319),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_190),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_257),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_291),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_320),
.B(n_327),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_321),
.A2(n_325),
.B1(n_332),
.B2(n_245),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_282),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_309),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_281),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_335),
.Y(n_337)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_329),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_311),
.A2(n_299),
.B(n_293),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_328),
.B(n_334),
.Y(n_346)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_305),
.B(n_287),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_331),
.B(n_190),
.Y(n_349)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_310),
.A3(n_315),
.B1(n_317),
.B2(n_318),
.C1(n_300),
.C2(n_191),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_341),
.B(n_343),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_300),
.C(n_202),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_345),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_209),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_322),
.Y(n_345)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_347),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_333),
.C(n_324),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_348),
.B(n_349),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_339),
.A2(n_340),
.B1(n_332),
.B2(n_333),
.Y(n_351)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_338),
.A2(n_321),
.B(n_323),
.Y(n_352)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_336),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_360),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_335),
.C(n_211),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_185),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_346),
.A2(n_245),
.B(n_191),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_339),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_361),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_355),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_369),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_344),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_10),
.B(n_11),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_364),
.B(n_360),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_6),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_368),
.A2(n_358),
.B1(n_359),
.B2(n_354),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_356),
.B(n_359),
.Y(n_369)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_373),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_367),
.A2(n_350),
.B(n_11),
.Y(n_373)
);

AOI21x1_ASAP7_75t_L g380 ( 
.A1(n_375),
.A2(n_368),
.B(n_361),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_10),
.C(n_11),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_12),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_380),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_374),
.B(n_372),
.Y(n_382)
);

AO221x1_ASAP7_75t_L g383 ( 
.A1(n_382),
.A2(n_377),
.B1(n_366),
.B2(n_380),
.C(n_371),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_381),
.B(n_365),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_12),
.B(n_14),
.Y(n_385)
);

AO21x1_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_14),
.B(n_15),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_386),
.B(n_15),
.Y(n_387)
);


endmodule