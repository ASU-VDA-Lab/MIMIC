module fake_jpeg_12473_n_592 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_592);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_592;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_9),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_38),
.B(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_61),
.B(n_88),
.Y(n_155)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_63),
.B(n_84),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_22),
.B(n_10),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_66),
.B(n_83),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_68),
.Y(n_204)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_71),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_24),
.B(n_18),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_77),
.B(n_125),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_80),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_82),
.B(n_92),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_22),
.B(n_10),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_11),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_11),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_31),
.B(n_9),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_117),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_43),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_12),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_94),
.B(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_97),
.B(n_109),
.Y(n_161)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_98),
.Y(n_129)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx9p33_ASAP7_75t_R g100 ( 
.A(n_23),
.Y(n_100)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx5_ASAP7_75t_SL g106 ( 
.A(n_23),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_106),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_49),
.B(n_12),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_54),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_127),
.Y(n_174)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_54),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_45),
.B(n_12),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_15),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_57),
.B1(n_48),
.B2(n_41),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_133),
.A2(n_156),
.B1(n_162),
.B2(n_164),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_77),
.A2(n_54),
.B1(n_35),
.B2(n_58),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_136),
.A2(n_137),
.B1(n_154),
.B2(n_160),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_48),
.B1(n_35),
.B2(n_58),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_48),
.B1(n_53),
.B2(n_41),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_140),
.A2(n_151),
.B1(n_153),
.B2(n_168),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_96),
.A2(n_26),
.B1(n_56),
.B2(n_30),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_103),
.A2(n_26),
.B1(n_56),
.B2(n_30),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_110),
.A2(n_57),
.B1(n_55),
.B2(n_50),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_29),
.B1(n_36),
.B2(n_28),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_55),
.B1(n_50),
.B2(n_44),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_69),
.A2(n_36),
.B1(n_29),
.B2(n_28),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_71),
.A2(n_36),
.B1(n_28),
.B2(n_39),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_166),
.B(n_187),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_64),
.A2(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_70),
.A2(n_85),
.B1(n_86),
.B2(n_36),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_172),
.A2(n_188),
.B1(n_197),
.B2(n_107),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_42),
.B1(n_28),
.B2(n_36),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_175),
.A2(n_200),
.B1(n_206),
.B2(n_98),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_95),
.B(n_62),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_181),
.B(n_189),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_65),
.B(n_8),
.C(n_17),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_14),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_8),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_70),
.A2(n_7),
.B1(n_17),
.B2(n_4),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_105),
.B(n_116),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_62),
.B(n_13),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_191),
.B(n_198),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_114),
.A2(n_13),
.B1(n_17),
.B2(n_4),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_120),
.B(n_126),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_104),
.A2(n_13),
.B1(n_16),
.B2(n_5),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_115),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_208),
.B(n_209),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_78),
.B(n_6),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_122),
.B(n_6),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_210),
.B(n_197),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_89),
.B(n_18),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_121),
.B(n_14),
.Y(n_216)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_214),
.B(n_216),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_2),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_215),
.B(n_226),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_173),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_217),
.B(n_223),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_218),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_222),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_73),
.Y(n_223)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_224),
.Y(n_325)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_136),
.B(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_136),
.B(n_3),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_227),
.B(n_249),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_228),
.Y(n_337)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_229),
.Y(n_326)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_233),
.Y(n_298)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_131),
.Y(n_234)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_234),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_72),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_161),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_237),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_174),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_145),
.Y(n_239)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_134),
.B(n_72),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_240),
.Y(n_316)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_243),
.Y(n_331)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_145),
.A2(n_74),
.B1(n_81),
.B2(n_118),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_246),
.A2(n_248),
.B1(n_267),
.B2(n_276),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_247),
.A2(n_253),
.B1(n_260),
.B2(n_261),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_16),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_146),
.B(n_73),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_250),
.Y(n_303)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_252),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_167),
.A2(n_113),
.B1(n_76),
.B2(n_90),
.Y(n_253)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_149),
.Y(n_254)
);

INVx11_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_255),
.Y(n_332)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_132),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_257),
.B(n_258),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_144),
.B(n_78),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_201),
.B(n_90),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_262),
.Y(n_328)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_132),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

BUFx4f_ASAP7_75t_SL g262 ( 
.A(n_149),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_170),
.A2(n_108),
.B1(n_124),
.B2(n_123),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_164),
.B(n_188),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_149),
.B(n_212),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_269),
.Y(n_308)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_185),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_266),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_167),
.A2(n_108),
.B1(n_124),
.B2(n_101),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_150),
.B(n_125),
.Y(n_269)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_142),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_176),
.Y(n_273)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_142),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_150),
.B(n_205),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_207),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_157),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_190),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_282),
.B1(n_283),
.B2(n_148),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_151),
.B(n_153),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_281),
.C(n_284),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_156),
.B(n_203),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_178),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_178),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_203),
.B(n_157),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_139),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_291),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_248),
.A2(n_172),
.B1(n_162),
.B2(n_133),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_301),
.A2(n_310),
.B1(n_314),
.B2(n_340),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_302),
.A2(n_290),
.B(n_294),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_140),
.B1(n_193),
.B2(n_176),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_309),
.A2(n_335),
.B1(n_339),
.B2(n_192),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_226),
.A2(n_193),
.B1(n_165),
.B2(n_139),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_227),
.A2(n_165),
.B1(n_163),
.B2(n_177),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_268),
.A2(n_177),
.B1(n_163),
.B2(n_159),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_318),
.A2(n_333),
.B1(n_239),
.B2(n_266),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_215),
.B(n_129),
.C(n_138),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_327),
.C(n_338),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_264),
.B(n_244),
.C(n_257),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_268),
.A2(n_159),
.B1(n_138),
.B2(n_195),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_271),
.A2(n_129),
.B1(n_135),
.B2(n_159),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_249),
.B(n_207),
.C(n_195),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_280),
.A2(n_135),
.B1(n_192),
.B2(n_180),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_241),
.A2(n_281),
.B1(n_270),
.B2(n_263),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_235),
.B(n_207),
.C(n_180),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_243),
.C(n_218),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_221),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_343),
.B(n_344),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_217),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_320),
.A2(n_284),
.B1(n_255),
.B2(n_251),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_345),
.A2(n_348),
.B1(n_352),
.B2(n_357),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_346),
.A2(n_349),
.B1(n_351),
.B2(n_368),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_222),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_370),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_309),
.A2(n_275),
.B1(n_273),
.B2(n_225),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_310),
.A2(n_314),
.B1(n_340),
.B2(n_301),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_233),
.B1(n_242),
.B2(n_229),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_232),
.C(n_220),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_372),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_302),
.A2(n_283),
.B(n_282),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_306),
.A2(n_148),
.B1(n_245),
.B2(n_234),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_286),
.B(n_213),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_356),
.B(n_365),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_285),
.B1(n_231),
.B2(n_224),
.Y(n_357)
);

AO21x1_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_256),
.B(n_260),
.Y(n_358)
);

AO22x1_ASAP7_75t_L g409 ( 
.A1(n_358),
.A2(n_332),
.B1(n_300),
.B2(n_323),
.Y(n_409)
);

A2O1A1O1Ixp25_ASAP7_75t_L g359 ( 
.A1(n_322),
.A2(n_254),
.B(n_262),
.C(n_261),
.D(n_205),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_359),
.A2(n_369),
.B(n_376),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_326),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_366),
.Y(n_402)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_286),
.B(n_274),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_315),
.B(n_262),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_322),
.A2(n_278),
.B1(n_219),
.B2(n_228),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_315),
.A2(n_290),
.B1(n_316),
.B2(n_338),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_272),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_230),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_377),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_290),
.A2(n_308),
.B1(n_336),
.B2(n_316),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_374),
.A2(n_334),
.B1(n_305),
.B2(n_329),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_311),
.Y(n_375)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_341),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_303),
.C(n_328),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_384),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_303),
.B(n_298),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_380),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_293),
.B(n_328),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_293),
.B(n_317),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_381),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_334),
.A2(n_317),
.B1(n_298),
.B2(n_295),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_382),
.A2(n_364),
.B1(n_352),
.B2(n_357),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_304),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_383),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_295),
.B(n_292),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_292),
.B(n_330),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_296),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_325),
.B1(n_324),
.B2(n_289),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_394),
.A2(n_383),
.B1(n_367),
.B2(n_289),
.Y(n_444)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_385),
.Y(n_396)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_349),
.A2(n_324),
.B1(n_325),
.B2(n_329),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_398),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_350),
.A2(n_332),
.B1(n_305),
.B2(n_307),
.Y(n_398)
);

NOR4xp25_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_304),
.C(n_331),
.D(n_296),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_403),
.B(n_380),
.Y(n_429)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_407),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_386),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_409),
.A2(n_414),
.B(n_346),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_350),
.A2(n_313),
.B1(n_337),
.B2(n_300),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_419),
.Y(n_431)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_347),
.A2(n_313),
.B1(n_337),
.B2(n_323),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_288),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_354),
.B(n_331),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_376),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_423),
.A2(n_433),
.B(n_436),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_402),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_425),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_414),
.A2(n_369),
.B1(n_373),
.B2(n_351),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_426),
.A2(n_447),
.B1(n_398),
.B2(n_397),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_427),
.B(n_409),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_429),
.Y(n_468)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_417),
.B(n_356),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_432),
.B(n_411),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_395),
.A2(n_366),
.B(n_355),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_371),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_439),
.C(n_440),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_395),
.A2(n_372),
.B(n_358),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_419),
.A2(n_348),
.B(n_358),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_438),
.A2(n_451),
.B(n_453),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_371),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_371),
.C(n_353),
.Y(n_440)
);

AO32x1_ASAP7_75t_L g442 ( 
.A1(n_422),
.A2(n_359),
.A3(n_379),
.B1(n_374),
.B2(n_378),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_442),
.A2(n_406),
.B(n_409),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_370),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_445),
.C(n_446),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_444),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_372),
.C(n_345),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_400),
.B(n_365),
.C(n_381),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_399),
.A2(n_368),
.B1(n_361),
.B2(n_343),
.Y(n_447)
);

OAI32xp33_ASAP7_75t_L g448 ( 
.A1(n_396),
.A2(n_344),
.A3(n_359),
.B1(n_288),
.B2(n_299),
.Y(n_448)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_360),
.C(n_299),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_450),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_388),
.A2(n_367),
.B(n_412),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_408),
.C(n_388),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_422),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_412),
.A2(n_418),
.B1(n_389),
.B2(n_387),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_417),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_415),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_453),
.A2(n_399),
.B1(n_410),
.B2(n_407),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_472),
.B1(n_438),
.B2(n_437),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_431),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_456),
.B(n_459),
.Y(n_502)
);

XOR2x2_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_408),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_462),
.A2(n_474),
.B1(n_441),
.B2(n_435),
.Y(n_507)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_428),
.Y(n_464)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_467),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_420),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_471),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_393),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_424),
.A2(n_387),
.B1(n_393),
.B2(n_422),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_413),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_476),
.C(n_479),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_426),
.A2(n_422),
.B1(n_406),
.B2(n_415),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_431),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_475),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_477),
.A2(n_481),
.B(n_429),
.Y(n_506)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_428),
.Y(n_478)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_390),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_423),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_423),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_465),
.B(n_425),
.Y(n_484)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_484),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_493),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_490),
.A2(n_506),
.B(n_507),
.Y(n_528)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_442),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_492),
.B(n_457),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_455),
.A2(n_447),
.B1(n_438),
.B2(n_442),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_463),
.A2(n_438),
.B1(n_454),
.B2(n_437),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_494),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_445),
.C(n_449),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_500),
.C(n_508),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_463),
.A2(n_472),
.B1(n_468),
.B2(n_473),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_499),
.Y(n_518)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_464),
.Y(n_498)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_498),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_435),
.B1(n_441),
.B2(n_446),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_461),
.B(n_436),
.C(n_450),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_465),
.B(n_432),
.Y(n_501)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_501),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_466),
.B(n_448),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_503),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_427),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_504),
.A2(n_493),
.B(n_503),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_471),
.B(n_451),
.C(n_433),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_390),
.C(n_392),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_457),
.C(n_481),
.Y(n_516)
);

AOI321xp33_ASAP7_75t_L g511 ( 
.A1(n_502),
.A2(n_459),
.A3(n_483),
.B1(n_479),
.B2(n_477),
.C(n_460),
.Y(n_511)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_511),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_469),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_513),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_505),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_480),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_529),
.C(n_492),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_516),
.B(n_524),
.Y(n_542)
);

INVx13_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_523),
.A2(n_487),
.B1(n_489),
.B2(n_501),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_460),
.C(n_482),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_526),
.A2(n_508),
.B(n_507),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_482),
.C(n_462),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_527),
.B(n_530),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_500),
.B(n_392),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g530 ( 
.A(n_489),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_517),
.A2(n_504),
.B(n_506),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_532),
.A2(n_535),
.B(n_526),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_L g533 ( 
.A1(n_522),
.A2(n_490),
.B(n_498),
.C(n_497),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_533),
.B(n_538),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_534),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_513),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_499),
.C(n_496),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_539),
.B(n_516),
.Y(n_553)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_521),
.Y(n_541)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_541),
.Y(n_559)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_525),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_543),
.B(n_544),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_518),
.A2(n_494),
.B1(n_488),
.B2(n_470),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_515),
.B(n_497),
.C(n_486),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_529),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_540),
.B(n_520),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_548),
.A2(n_552),
.B(n_560),
.Y(n_561)
);

OAI21xp33_ASAP7_75t_SL g549 ( 
.A1(n_532),
.A2(n_525),
.B(n_486),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_549),
.B(n_551),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_546),
.B(n_491),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_531),
.A2(n_524),
.B(n_510),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_553),
.B(n_555),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_554),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_535),
.A2(n_510),
.B1(n_528),
.B2(n_527),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_531),
.A2(n_528),
.B1(n_470),
.B2(n_487),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_557),
.B(n_558),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_560),
.A2(n_542),
.B(n_545),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_SL g579 ( 
.A(n_562),
.B(n_523),
.C(n_458),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_538),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_566),
.A2(n_567),
.B(n_569),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_537),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_552),
.A2(n_533),
.B(n_539),
.Y(n_568)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_568),
.A2(n_556),
.B(n_511),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_555),
.B(n_537),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_514),
.C(n_512),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_571),
.B(n_536),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_563),
.A2(n_548),
.B(n_557),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_572),
.B(n_573),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_578),
.C(n_579),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_561),
.A2(n_553),
.B(n_559),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_576),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_570),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_577),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_564),
.A2(n_458),
.B1(n_405),
.B2(n_416),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_571),
.C(n_561),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_584),
.A2(n_565),
.B(n_568),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_580),
.Y(n_585)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_585),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_586),
.A2(n_587),
.B(n_404),
.Y(n_588)
);

NAND4xp25_ASAP7_75t_L g587 ( 
.A(n_581),
.B(n_574),
.C(n_583),
.D(n_582),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_588),
.B(n_589),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_430),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_430),
.Y(n_592)
);


endmodule