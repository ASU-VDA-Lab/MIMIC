module fake_jpeg_28840_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_68),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_43),
.C(n_49),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_3),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_48),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_50),
.Y(n_97)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_60),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_88),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_58),
.B1(n_47),
.B2(n_59),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_97),
.B(n_7),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_25),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_26),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_7),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_83),
.B(n_5),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_105),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_4),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_121),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_5),
.C(n_6),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_29),
.B(n_42),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_109),
.B(n_113),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_28),
.B(n_41),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_116),
.B(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_23),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_8),
.C(n_10),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_14),
.B(n_18),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_12),
.C(n_13),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_106),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_130),
.A2(n_132),
.B(n_38),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_36),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_112),
.C(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_135),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_128),
.C(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_128),
.C(n_141),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_126),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_123),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_133),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_138),
.Y(n_148)
);


endmodule