module real_aes_8994_n_254 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_254);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_254;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_666;
wire n_320;
wire n_551;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_397;
wire n_663;
wire n_385;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_283;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_0), .A2(n_234), .B1(n_561), .B2(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_1), .A2(n_236), .B1(n_404), .B2(n_407), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_2), .A2(n_29), .B1(n_522), .B2(n_582), .C(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_3), .B(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_SL g727 ( .A1(n_4), .A2(n_52), .B1(n_534), .B2(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_5), .A2(n_14), .B1(n_350), .B2(n_526), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_6), .B(n_505), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_7), .A2(n_251), .B1(n_505), .B2(n_537), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_8), .A2(n_114), .B1(n_468), .B2(n_537), .Y(n_536) );
XOR2x2_ASAP7_75t_L g574 ( .A(n_9), .B(n_575), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_10), .A2(n_172), .B1(n_358), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_11), .A2(n_130), .B1(n_603), .B2(n_605), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_12), .A2(n_211), .B1(n_587), .B2(n_610), .C(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_13), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_15), .A2(n_23), .B1(n_318), .B2(n_407), .Y(n_555) );
INVx1_ASAP7_75t_L g510 ( .A(n_16), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_17), .A2(n_244), .B1(n_407), .B2(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_18), .A2(n_166), .B1(n_394), .B2(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_19), .Y(n_436) );
AO22x2_ASAP7_75t_L g283 ( .A1(n_20), .A2(n_78), .B1(n_284), .B2(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g743 ( .A(n_20), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_21), .Y(n_361) );
AOI22xp5_ASAP7_75t_SL g726 ( .A1(n_22), .A2(n_249), .B1(n_445), .B2(n_561), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_24), .A2(n_57), .B1(n_623), .B2(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_25), .B(n_549), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_26), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_27), .A2(n_134), .B1(n_387), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_28), .A2(n_184), .B1(n_345), .B2(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_30), .A2(n_156), .B1(n_392), .B2(n_527), .Y(n_802) );
AOI22xp5_ASAP7_75t_SL g722 ( .A1(n_31), .A2(n_149), .B1(n_368), .B2(n_560), .Y(n_722) );
AO22x1_ASAP7_75t_L g629 ( .A1(n_32), .A2(n_630), .B1(n_662), .B2(n_663), .Y(n_629) );
INVx1_ASAP7_75t_L g662 ( .A(n_32), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_33), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_34), .A2(n_48), .B1(n_309), .B2(n_316), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_35), .A2(n_213), .B1(n_340), .B2(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_36), .A2(n_242), .B1(n_449), .B2(n_685), .Y(n_684) );
AOI222xp33_ASAP7_75t_L g709 ( .A1(n_37), .A2(n_116), .B1(n_187), .B2(n_309), .C1(n_316), .C2(n_414), .Y(n_709) );
AO22x2_ASAP7_75t_L g287 ( .A1(n_38), .A2(n_79), .B1(n_284), .B2(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g744 ( .A(n_38), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_39), .Y(n_415) );
INVx1_ASAP7_75t_L g784 ( .A(n_40), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_41), .A2(n_59), .B1(n_407), .B2(n_507), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_42), .A2(n_192), .B1(n_408), .B2(n_507), .Y(n_678) );
AOI222xp33_ASAP7_75t_L g540 ( .A1(n_43), .A2(n_148), .B1(n_204), .B2(n_302), .C1(n_500), .C2(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_44), .Y(n_307) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_45), .A2(n_73), .B1(n_612), .B2(n_613), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_46), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_47), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_49), .A2(n_224), .B1(n_368), .B2(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_50), .A2(n_596), .B1(n_597), .B2(n_626), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_50), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_51), .A2(n_238), .B1(n_653), .B2(n_654), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_53), .A2(n_131), .B1(n_405), .B2(n_407), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_54), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_55), .A2(n_189), .B1(n_394), .B2(n_396), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_56), .A2(n_227), .B1(n_449), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_58), .A2(n_119), .B1(n_336), .B2(n_368), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_60), .A2(n_180), .B1(n_395), .B2(n_478), .Y(n_477) );
AOI222xp33_ASAP7_75t_L g765 ( .A1(n_61), .A2(n_82), .B1(n_142), .B2(n_603), .C1(n_644), .C2(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_62), .B(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_63), .A2(n_104), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_64), .A2(n_138), .B1(n_404), .B2(n_411), .Y(n_551) );
INVx1_ASAP7_75t_L g591 ( .A(n_65), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_66), .A2(n_120), .B1(n_485), .B2(n_683), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_67), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_68), .A2(n_117), .B1(n_447), .B2(n_753), .C(n_754), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_69), .A2(n_235), .B1(n_509), .B2(n_589), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_70), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_71), .A2(n_239), .B1(n_319), .B2(n_593), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_72), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_74), .A2(n_202), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_75), .A2(n_137), .B1(n_386), .B2(n_388), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_76), .A2(n_199), .B1(n_408), .B2(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_77), .A2(n_115), .B1(n_392), .B2(n_447), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_80), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_81), .B(n_610), .Y(n_719) );
INVx1_ASAP7_75t_L g262 ( .A(n_83), .Y(n_262) );
AOI211xp5_ASAP7_75t_L g254 ( .A1(n_84), .A2(n_255), .B(n_263), .C(n_745), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_85), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_86), .A2(n_146), .B1(n_445), .B2(n_533), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_87), .A2(n_127), .B1(n_310), .B2(n_318), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_88), .A2(n_178), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_89), .A2(n_101), .B1(n_340), .B2(n_524), .Y(n_697) );
INVx1_ASAP7_75t_L g258 ( .A(n_90), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_91), .A2(n_100), .B1(n_392), .B2(n_442), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_92), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_93), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_94), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_95), .A2(n_111), .B1(n_524), .B2(n_530), .Y(n_661) );
OA22x2_ASAP7_75t_L g423 ( .A1(n_96), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_96), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_97), .A2(n_132), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_98), .A2(n_99), .B1(n_388), .B2(n_619), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_102), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_103), .A2(n_203), .B1(n_336), .B2(n_340), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_105), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_106), .A2(n_113), .B1(n_522), .B2(n_524), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_107), .A2(n_161), .B1(n_318), .B2(n_603), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_108), .A2(n_152), .B1(n_683), .B2(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_109), .Y(n_498) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_110), .A2(n_206), .B1(n_346), .B2(n_360), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_112), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_118), .A2(n_250), .B1(n_624), .B2(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_121), .Y(n_763) );
XNOR2x2_ASAP7_75t_L g518 ( .A(n_122), .B(n_519), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_123), .A2(n_147), .B1(n_534), .B2(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_124), .A2(n_165), .B1(n_340), .B2(n_391), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_125), .Y(n_495) );
AND2x2_ASAP7_75t_L g261 ( .A(n_126), .B(n_262), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_128), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_129), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_133), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_135), .A2(n_205), .B1(n_392), .B2(n_485), .Y(n_484) );
OA22x2_ASAP7_75t_L g543 ( .A1(n_136), .A2(n_544), .B1(n_545), .B2(n_566), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_136), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_139), .B(n_302), .Y(n_434) );
INVx1_ASAP7_75t_L g790 ( .A(n_140), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_141), .B(n_472), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_143), .A2(n_248), .B1(n_345), .B2(n_350), .Y(n_344) );
AND2x6_ASAP7_75t_L g257 ( .A(n_144), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_144), .Y(n_737) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_145), .A2(n_216), .B1(n_284), .B2(n_288), .Y(n_293) );
INVx1_ASAP7_75t_L g792 ( .A(n_150), .Y(n_792) );
AOI22xp5_ASAP7_75t_SL g723 ( .A1(n_151), .A2(n_215), .B1(n_442), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g444 ( .A1(n_153), .A2(n_223), .B1(n_445), .B2(n_447), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_154), .Y(n_675) );
INVx1_ASAP7_75t_L g778 ( .A(n_155), .Y(n_778) );
OA22x2_ASAP7_75t_L g779 ( .A1(n_155), .A2(n_778), .B1(n_780), .B2(n_781), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_157), .A2(n_233), .B1(n_507), .B2(n_509), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_158), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_159), .A2(n_201), .B1(n_311), .B2(n_405), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_160), .B(n_610), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_162), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_163), .A2(n_229), .B1(n_351), .B2(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_164), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_167), .A2(n_175), .B1(n_396), .B2(n_449), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_168), .A2(n_253), .B1(n_586), .B2(n_587), .Y(n_585) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_169), .A2(n_226), .B1(n_284), .B2(n_285), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_170), .A2(n_200), .B1(n_407), .B2(n_465), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_171), .A2(n_212), .B1(n_478), .B2(n_560), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_173), .A2(n_377), .B1(n_420), .B2(n_421), .Y(n_376) );
INVx1_ASAP7_75t_L g420 ( .A(n_173), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_174), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_176), .A2(n_198), .B1(n_310), .B2(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_177), .A2(n_237), .B1(n_387), .B2(n_442), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_179), .B(n_608), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_181), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_182), .A2(n_208), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_183), .A2(n_207), .B1(n_533), .B2(n_534), .Y(n_532) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_185), .A2(n_195), .B1(n_541), .B2(n_644), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_186), .Y(n_701) );
INVx1_ASAP7_75t_L g729 ( .A(n_188), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_190), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_191), .A2(n_243), .B1(n_388), .B2(n_526), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_193), .A2(n_194), .B1(n_449), .B2(n_534), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_196), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_197), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_209), .Y(n_370) );
OA22x2_ASAP7_75t_L g669 ( .A1(n_210), .A2(n_670), .B1(n_671), .B2(n_692), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_210), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_214), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_216), .B(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_217), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_218), .Y(n_384) );
INVx1_ASAP7_75t_L g787 ( .A(n_219), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_220), .A2(n_252), .B1(n_342), .B2(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_221), .Y(n_645) );
INVx1_ASAP7_75t_L g785 ( .A(n_222), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_225), .Y(n_462) );
INVx1_ASAP7_75t_L g740 ( .A(n_226), .Y(n_740) );
OA22x2_ASAP7_75t_L g271 ( .A1(n_228), .A2(n_272), .B1(n_273), .B2(n_274), .Y(n_271) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_228), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_230), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_231), .B(n_610), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_232), .Y(n_356) );
INVx1_ASAP7_75t_L g284 ( .A(n_240), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_240), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_241), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_245), .B(n_549), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_246), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_247), .A2(n_747), .B1(n_767), .B2(n_768), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_247), .Y(n_767) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_258), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_259), .A2(n_735), .B(n_777), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_260), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_666), .B1(n_667), .B2(n_731), .C(n_732), .Y(n_263) );
INVx1_ASAP7_75t_L g731 ( .A(n_264), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B1(n_514), .B2(n_665), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
XNOR2xp5_ASAP7_75t_SL g267 ( .A(n_268), .B(n_422), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B1(n_374), .B2(n_375), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_333), .Y(n_274) );
NOR3xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_300), .C(n_321), .Y(n_275) );
OAI22xp5_ASAP7_75t_SL g276 ( .A1(n_277), .A2(n_294), .B1(n_295), .B2(n_299), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI221xp5_ASAP7_75t_SL g398 ( .A1(n_279), .A2(n_399), .B1(n_400), .B2(n_402), .C(n_403), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_279), .A2(n_295), .B1(n_784), .B2(n_785), .Y(n_783) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx3_ASAP7_75t_L g430 ( .A(n_280), .Y(n_430) );
INVx2_ASAP7_75t_L g635 ( .A(n_280), .Y(n_635) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_289), .Y(n_280) );
INVx2_ASAP7_75t_L g343 ( .A(n_281), .Y(n_343) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_287), .Y(n_281) );
AND2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_287), .Y(n_298) );
AND2x2_ASAP7_75t_L g339 ( .A(n_282), .B(n_314), .Y(n_339) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g304 ( .A(n_283), .B(n_287), .Y(n_304) );
AND2x2_ASAP7_75t_L g315 ( .A(n_283), .B(n_293), .Y(n_315) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g288 ( .A(n_286), .Y(n_288) );
INVx2_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
INVx1_ASAP7_75t_L g353 ( .A(n_287), .Y(n_353) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_290), .B(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_L g369 ( .A(n_290), .B(n_339), .Y(n_369) );
AND2x4_ASAP7_75t_L g470 ( .A(n_290), .B(n_343), .Y(n_470) );
AND2x6_ASAP7_75t_L g472 ( .A(n_290), .B(n_298), .Y(n_472) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g306 ( .A(n_291), .Y(n_306) );
INVx1_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
INVx1_ASAP7_75t_L g331 ( .A(n_291), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_291), .B(n_293), .Y(n_354) );
AND2x2_ASAP7_75t_L g305 ( .A(n_292), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g349 ( .A(n_293), .B(n_331), .Y(n_349) );
BUFx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g401 ( .A(n_296), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_296), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_428) );
BUFx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g638 ( .A(n_297), .Y(n_638) );
AND2x2_ASAP7_75t_L g348 ( .A(n_298), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g360 ( .A(n_298), .B(n_305), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_298), .B(n_349), .Y(n_757) );
OAI21xp33_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_307), .B(n_308), .Y(n_300) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_301), .A2(n_591), .B(n_592), .Y(n_590) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_303), .Y(n_414) );
INVx4_ASAP7_75t_L g463 ( .A(n_303), .Y(n_463) );
INVx2_ASAP7_75t_L g674 ( .A(n_303), .Y(n_674) );
AND2x6_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g328 ( .A(n_304), .Y(n_328) );
AND2x4_ASAP7_75t_L g408 ( .A(n_304), .B(n_330), .Y(n_408) );
AND2x2_ASAP7_75t_L g338 ( .A(n_305), .B(n_339), .Y(n_338) );
AND2x6_ASAP7_75t_L g342 ( .A(n_305), .B(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx4_ASAP7_75t_L g604 ( .A(n_310), .Y(n_604) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_311), .Y(n_411) );
BUFx2_ASAP7_75t_L g541 ( .A(n_311), .Y(n_541) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_311), .Y(n_593) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g320 ( .A(n_313), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_314), .Y(n_323) );
AND2x4_ASAP7_75t_L g319 ( .A(n_315), .B(n_320), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_315), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g405 ( .A(n_315), .B(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx4f_ASAP7_75t_SL g500 ( .A(n_318), .Y(n_500) );
BUFx12f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_319), .Y(n_418) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_319), .Y(n_465) );
OAI22xp33_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_324), .B1(n_325), .B2(n_332), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_322), .A2(n_327), .B1(n_436), .B2(n_437), .Y(n_435) );
BUFx3_ASAP7_75t_L g648 ( .A(n_322), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_322), .A2(n_790), .B1(n_791), .B2(n_792), .Y(n_789) );
AND2x2_ASAP7_75t_L g459 ( .A(n_323), .B(n_373), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_325), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_646) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g764 ( .A(n_326), .Y(n_764) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_327), .Y(n_326) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_355), .C(n_365), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_344), .Y(n_334) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g699 ( .A(n_337), .Y(n_699) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_338), .Y(n_395) );
BUFx2_ASAP7_75t_SL g560 ( .A(n_338), .Y(n_560) );
BUFx2_ASAP7_75t_SL g582 ( .A(n_338), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_339), .B(n_349), .Y(n_364) );
AND2x4_ASAP7_75t_L g372 ( .A(n_339), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g446 ( .A(n_339), .B(n_349), .Y(n_446) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_341), .A2(n_359), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx4_ASAP7_75t_L g533 ( .A(n_341), .Y(n_533) );
INVx5_ASAP7_75t_SL g796 ( .A(n_341), .Y(n_796) );
INVx11_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx11_ASAP7_75t_L g450 ( .A(n_342), .Y(n_450) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g488 ( .A(n_346), .Y(n_488) );
BUFx2_ASAP7_75t_L g724 ( .A(n_346), .Y(n_724) );
INVx4_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
INVx5_ASAP7_75t_L g441 ( .A(n_347), .Y(n_441) );
INVx3_ASAP7_75t_L g526 ( .A(n_347), .Y(n_526) );
INVx1_ASAP7_75t_L g564 ( .A(n_347), .Y(n_564) );
BUFx3_ASAP7_75t_L g620 ( .A(n_347), .Y(n_620) );
INVx8_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g442 ( .A(n_351), .Y(n_442) );
BUFx4f_ASAP7_75t_SL g657 ( .A(n_351), .Y(n_657) );
INVx6_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g388 ( .A(n_352), .Y(n_388) );
INVx1_ASAP7_75t_L g527 ( .A(n_352), .Y(n_527) );
OR2x6_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g406 ( .A(n_353), .Y(n_406) );
INVx1_ASAP7_75t_L g373 ( .A(n_354), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_361), .B2(n_362), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_357), .A2(n_380), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g534 ( .A(n_359), .Y(n_534) );
INVx2_ASAP7_75t_L g660 ( .A(n_359), .Y(n_660) );
INVx3_ASAP7_75t_L g707 ( .A(n_359), .Y(n_707) );
INVx6_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g396 ( .A(n_360), .Y(n_396) );
BUFx3_ASAP7_75t_L g685 ( .A(n_360), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_362), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_370), .B2(n_371), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g392 ( .A(n_369), .Y(n_392) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_369), .Y(n_458) );
INVx2_ASAP7_75t_L g655 ( .A(n_369), .Y(n_655) );
BUFx3_ASAP7_75t_L g690 ( .A(n_369), .Y(n_690) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_372), .Y(n_383) );
BUFx3_ASAP7_75t_L g447 ( .A(n_372), .Y(n_447) );
BUFx3_ASAP7_75t_L g478 ( .A(n_372), .Y(n_478) );
BUFx2_ASAP7_75t_SL g485 ( .A(n_372), .Y(n_485) );
BUFx3_ASAP7_75t_L g524 ( .A(n_372), .Y(n_524) );
BUFx2_ASAP7_75t_L g561 ( .A(n_372), .Y(n_561) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g421 ( .A(n_377), .Y(n_421) );
AND2x2_ASAP7_75t_SL g377 ( .A(n_378), .B(n_397), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_389), .Y(n_378) );
OAI221xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_381), .B1(n_382), .B2(n_384), .C(n_385), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .Y(n_389) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g494 ( .A(n_395), .Y(n_494) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_395), .Y(n_623) );
BUFx3_ASAP7_75t_L g653 ( .A(n_395), .Y(n_653) );
NOR2xp33_ASAP7_75t_SL g397 ( .A(n_398), .B(n_409), .Y(n_397) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g508 ( .A(n_405), .Y(n_508) );
BUFx3_ASAP7_75t_L g589 ( .A(n_405), .Y(n_589) );
INVx1_ASAP7_75t_SL g614 ( .A(n_407), .Y(n_614) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_SL g509 ( .A(n_408), .Y(n_509) );
OAI222xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_413), .B2(n_415), .C1(n_416), .C2(n_419), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
OAI222xp33_ASAP7_75t_L g639 ( .A1(n_413), .A2(n_640), .B1(n_641), .B2(n_642), .C1(n_643), .C2(n_645), .Y(n_639) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_413), .A2(n_787), .B(n_788), .Y(n_786) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g600 ( .A(n_414), .Y(n_600) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g644 ( .A(n_418), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_451), .B1(n_512), .B2(n_513), .Y(n_422) );
INVx2_ASAP7_75t_SL g512 ( .A(n_423), .Y(n_512) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND3x1_ASAP7_75t_L g426 ( .A(n_427), .B(n_438), .C(n_443), .Y(n_426) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .C(n_435), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_448), .Y(n_443) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g476 ( .A(n_446), .Y(n_476) );
BUFx3_ASAP7_75t_L g578 ( .A(n_446), .Y(n_578) );
BUFx3_ASAP7_75t_L g683 ( .A(n_446), .Y(n_683) );
INVx4_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g728 ( .A(n_450), .Y(n_728) );
INVx3_ASAP7_75t_L g753 ( .A(n_450), .Y(n_753) );
INVx1_ASAP7_75t_L g513 ( .A(n_451), .Y(n_513) );
OA22x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_480), .B2(n_511), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
XOR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_479), .Y(n_453) );
NAND3x1_ASAP7_75t_SL g454 ( .A(n_455), .B(n_460), .C(n_474), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVx4_ASAP7_75t_L g523 ( .A(n_458), .Y(n_523) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_466), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_464), .Y(n_461) );
OAI21xp5_ASAP7_75t_SL g497 ( .A1(n_463), .A2(n_498), .B(n_499), .Y(n_497) );
BUFx2_ASAP7_75t_L g553 ( .A(n_463), .Y(n_553) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_463), .A2(n_715), .B(n_716), .Y(n_714) );
INVx4_ASAP7_75t_L g766 ( .A(n_463), .Y(n_766) );
BUFx4f_ASAP7_75t_L g605 ( .A(n_465), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .C(n_473), .Y(n_466) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_468), .Y(n_610) );
INVx5_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g505 ( .A(n_469), .Y(n_505) );
INVx2_ASAP7_75t_L g586 ( .A(n_469), .Y(n_586) );
INVx4_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g503 ( .A(n_472), .Y(n_503) );
INVx1_ASAP7_75t_SL g538 ( .A(n_472), .Y(n_538) );
BUFx4f_ASAP7_75t_L g587 ( .A(n_472), .Y(n_587) );
BUFx2_ASAP7_75t_L g608 ( .A(n_472), .Y(n_608) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g531 ( .A(n_476), .Y(n_531) );
BUFx4f_ASAP7_75t_SL g624 ( .A(n_476), .Y(n_624) );
INVx1_ASAP7_75t_L g511 ( .A(n_480), .Y(n_511) );
XOR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_510), .Y(n_480) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_482), .B(n_496), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .C(n_492), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g688 ( .A(n_494), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .C(n_506), .Y(n_501) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g612 ( .A(n_508), .Y(n_612) );
INVx1_ASAP7_75t_L g665 ( .A(n_514), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_568), .B2(n_664), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_518), .B1(n_542), .B2(n_567), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND4xp75_ASAP7_75t_L g519 ( .A(n_520), .B(n_528), .C(n_535), .D(n_540), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g617 ( .A(n_523), .Y(n_617) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_SL g535 ( .A(n_536), .B(n_539), .Y(n_535) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_SL g549 ( .A(n_538), .Y(n_549) );
INVx1_ASAP7_75t_L g640 ( .A(n_541), .Y(n_640) );
INVx1_ASAP7_75t_L g567 ( .A(n_542), .Y(n_567) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_SL g566 ( .A(n_545), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_546), .B(n_556), .Y(n_545) );
NOR2xp67_ASAP7_75t_SL g546 ( .A(n_547), .B(n_552), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .C(n_551), .Y(n_547) );
OAI21xp5_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_554), .B(n_555), .Y(n_552) );
NOR2x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g664 ( .A(n_568), .Y(n_664) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_628), .B2(n_629), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AO22x1_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_594), .B1(n_595), .B2(n_627), .Y(n_573) );
INVx1_ASAP7_75t_SL g627 ( .A(n_574), .Y(n_627) );
NOR4xp75_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .C(n_584), .D(n_590), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_581), .B(n_583), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g791 ( .A(n_593), .Y(n_791) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g626 ( .A(n_597), .Y(n_626) );
NAND3x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_615), .C(n_621), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_606), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_601), .B(n_602), .Y(n_599) );
INVx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .C(n_611), .Y(n_606) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .Y(n_621) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g663 ( .A(n_630), .Y(n_663) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_650), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_639), .C(n_646), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_636), .B2(n_637), .Y(n_632) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g702 ( .A(n_638), .Y(n_702) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_648), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_658), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_656), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_657), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_693), .B2(n_730), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g692 ( .A(n_671), .Y(n_692) );
NAND2x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_680), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_677), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_675), .B(n_676), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_686), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx3_ASAP7_75t_L g801 ( .A(n_685), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_691), .Y(n_686) );
BUFx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g730 ( .A(n_693), .Y(n_730) );
XNOR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_711), .Y(n_693) );
XOR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_710), .Y(n_694) );
NAND4xp75_ASAP7_75t_L g695 ( .A(n_696), .B(n_700), .C(n_705), .D(n_709), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
OA211x2_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_703), .C(n_704), .Y(n_700) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
XOR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_729), .Y(n_711) );
NAND3x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_721), .C(n_725), .Y(n_712) );
NOR2x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .C(n_720), .Y(n_717) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_738), .Y(n_733) );
OR2x2_ASAP7_75t_SL g805 ( .A(n_734), .B(n_739), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_735), .Y(n_770) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_736), .B(n_774), .Y(n_777) );
CKINVDCx16_ASAP7_75t_R g774 ( .A(n_737), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
OAI322xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_769), .A3(n_771), .B1(n_775), .B2(n_778), .C1(n_779), .C2(n_803), .Y(n_745) );
INVx1_ASAP7_75t_L g768 ( .A(n_747), .Y(n_768) );
AND4x1_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .C(n_760), .D(n_765), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_754) );
BUFx2_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_793), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_786), .C(n_789), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_798), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .Y(n_798) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
endmodule