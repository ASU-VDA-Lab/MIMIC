module fake_jpeg_32121_n_293 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_17),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_32),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_9),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_55),
.Y(n_60)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_0),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_35),
.B1(n_26),
.B2(n_33),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_19),
.B1(n_28),
.B2(n_30),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_59),
.A2(n_71),
.B1(n_89),
.B2(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_26),
.B1(n_33),
.B2(n_20),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_92)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_84),
.Y(n_111)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_19),
.B1(n_28),
.B2(n_30),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_20),
.B1(n_28),
.B2(n_30),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_20),
.B1(n_25),
.B2(n_21),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_25),
.B1(n_21),
.B2(n_38),
.Y(n_74)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OA22x2_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_32),
.B1(n_37),
.B2(n_1),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_46),
.B1(n_53),
.B2(n_32),
.Y(n_98)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_31),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_24),
.B1(n_22),
.B2(n_38),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_102),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_53),
.B1(n_54),
.B2(n_43),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_97),
.A2(n_109),
.B1(n_114),
.B2(n_119),
.Y(n_146)
);

OR2x2_ASAP7_75t_SL g147 ( 
.A(n_98),
.B(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_100),
.B(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_60),
.B(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_46),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_45),
.B1(n_32),
.B2(n_3),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_80),
.B(n_58),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_54),
.B1(n_43),
.B2(n_0),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_124),
.B1(n_83),
.B2(n_76),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_59),
.B(n_2),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_116),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_113),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_5),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_121),
.CI(n_123),
.CON(n_137),
.SN(n_137)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_68),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_67),
.C(n_64),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_5),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_7),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_76),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_63),
.B(n_7),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_8),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_75),
.B(n_77),
.C(n_91),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_139),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_91),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_112),
.B(n_121),
.C(n_123),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_108),
.B1(n_114),
.B2(n_106),
.Y(n_169)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_149),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_122),
.B1(n_104),
.B2(n_99),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_10),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_70),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_112),
.B1(n_124),
.B2(n_119),
.Y(n_162)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_58),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

AO21x2_ASAP7_75t_L g156 ( 
.A1(n_98),
.A2(n_92),
.B(n_105),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_98),
.B1(n_120),
.B2(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_118),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_162),
.A2(n_167),
.B(n_172),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_179),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_112),
.B(n_93),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_173),
.B1(n_182),
.B2(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_98),
.B(n_125),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_184),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_104),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_137),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_134),
.B1(n_129),
.B2(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_107),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_132),
.C(n_137),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_122),
.B1(n_107),
.B2(n_94),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_94),
.B(n_127),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_176),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_204),
.B1(n_169),
.B2(n_184),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_156),
.B(n_152),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_201),
.B(n_185),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_199),
.C(n_203),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_161),
.B1(n_171),
.B2(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_156),
.B(n_136),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_156),
.C(n_151),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_156),
.B1(n_155),
.B2(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_135),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_135),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_211),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_208),
.A2(n_211),
.B(n_163),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_141),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_164),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_140),
.B(n_142),
.Y(n_211)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_171),
.B(n_142),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_198),
.B1(n_209),
.B2(n_208),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_173),
.A3(n_158),
.B1(n_163),
.B2(n_160),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_218),
.B(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_160),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_221),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_223),
.B1(n_226),
.B2(n_190),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_210),
.B(n_10),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_161),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_144),
.B1(n_185),
.B2(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_11),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_191),
.B(n_11),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_230),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_240),
.B1(n_238),
.B2(n_236),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_199),
.C(n_203),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_217),
.C(n_224),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_196),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_198),
.B1(n_204),
.B2(n_193),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_198),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_189),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_SL g245 ( 
.A(n_217),
.B(n_193),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_247),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_221),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_197),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_216),
.C(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_250),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_216),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_255),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_222),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_223),
.C(n_214),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_260),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_222),
.B1(n_231),
.B2(n_232),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_240),
.B1(n_231),
.B2(n_232),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_227),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_245),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_256),
.B1(n_252),
.B2(n_248),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_252),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_257),
.A2(n_238),
.B(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_267),
.A2(n_229),
.B1(n_12),
.B2(n_14),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_249),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_274),
.B1(n_267),
.B2(n_268),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_227),
.B1(n_230),
.B2(n_188),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_11),
.C(n_14),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_277),
.A2(n_264),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_261),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_273),
.B1(n_261),
.B2(n_275),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_281),
.B1(n_282),
.B2(n_15),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_17),
.B(n_15),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_279),
.B1(n_16),
.B2(n_15),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

OAI31xp33_ASAP7_75t_SL g291 ( 
.A1(n_290),
.A2(n_289),
.A3(n_287),
.B(n_285),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_288),
.B(n_286),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_292),
.Y(n_293)
);


endmodule