module real_jpeg_30840_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_650;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_0),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g390 ( 
.A(n_0),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_0),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_0),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_2),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_2),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_2),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_2),
.B(n_175),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_2),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_2),
.B(n_299),
.Y(n_298)
);

NAND2x1_ASAP7_75t_L g387 ( 
.A(n_2),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_3),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_3),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_3),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_3),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_3),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_3),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_3),
.B(n_437),
.Y(n_436)
);

AND2x4_ASAP7_75t_SL g207 ( 
.A(n_4),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_4),
.B(n_76),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_4),
.B(n_211),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g444 ( 
.A(n_4),
.B(n_445),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_4),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_4),
.B(n_277),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_4),
.B(n_373),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_4),
.B(n_580),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_5),
.B(n_238),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_5),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_5),
.B(n_419),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_5),
.B(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_5),
.B(n_529),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_5),
.B(n_546),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_5),
.B(n_553),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_R g90 ( 
.A(n_6),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_6),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_6),
.B(n_186),
.Y(n_185)
);

NAND2x1p5_ASAP7_75t_L g198 ( 
.A(n_6),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_7),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_9),
.Y(n_425)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_10),
.Y(n_454)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_11),
.Y(n_271)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_11),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_12),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_12),
.B(n_114),
.Y(n_225)
);

AND2x4_ASAP7_75t_SL g243 ( 
.A(n_12),
.B(n_244),
.Y(n_243)
);

AND2x4_ASAP7_75t_SL g272 ( 
.A(n_12),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_12),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_12),
.B(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_12),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_12),
.B(n_373),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_13),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_13),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_13),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_13),
.B(n_238),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_13),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_13),
.B(n_526),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_13),
.B(n_369),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_14),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_14),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_14),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_14),
.B(n_117),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_14),
.B(n_427),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_14),
.B(n_494),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_14),
.B(n_505),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_14),
.B(n_538),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B(n_650),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_15),
.B(n_651),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_16),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_16),
.B(n_38),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_16),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_16),
.B(n_432),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_16),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_16),
.B(n_576),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_17),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_17),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_17),
.Y(n_400)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_18),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_18),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_18),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_19),
.B(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_19),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_19),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_19),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_19),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_99),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_98),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_83),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_83),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_68),
.B(n_82),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_26),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_49),
.C(n_61),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_27),
.B(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_43),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_36),
.B2(n_42),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_42),
.C(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_29),
.A2(n_30),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_35),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_37),
.A2(n_52),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_37),
.Y(n_134)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_40),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_41),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_41),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_41),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_51),
.C(n_56),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_47),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_48),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_50),
.B(n_61),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_52),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_52),
.A2(n_133),
.B1(n_144),
.B2(n_313),
.Y(n_327)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2x2_ASAP7_75t_L g131 ( 
.A(n_56),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_60),
.Y(n_284)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_66),
.Y(n_395)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_85),
.C(n_86),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_88),
.B(n_96),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_155),
.B(n_649),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_153),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_102),
.B(n_153),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_148),
.C(n_150),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_104),
.B(n_344),
.Y(n_343)
);

MAJx2_ASAP7_75t_R g104 ( 
.A(n_105),
.B(n_131),
.C(n_135),
.Y(n_104)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_105),
.B(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_120),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_121),
.C(n_126),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.C(n_116),
.Y(n_106)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_107),
.B(n_116),
.Y(n_336)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_112),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_112),
.Y(n_420)
);

XOR2x1_ASAP7_75t_L g335 ( 
.A(n_113),
.B(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_130),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_131),
.B(n_352),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_136),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.C(n_144),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_138),
.B(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_144),
.A2(n_198),
.B1(n_202),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_144),
.Y(n_313)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_147),
.Y(n_549)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_149),
.B(n_151),
.Y(n_344)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21x1_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_358),
.B(n_643),
.Y(n_155)
);

NOR2xp67_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_342),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_314),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_158),
.B(n_314),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_229),
.C(n_285),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_160),
.A2(n_161),
.B1(n_286),
.B2(n_623),
.Y(n_622)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_203),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_162),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_178),
.C(n_192),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_164),
.B(n_627),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_166),
.B(n_173),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_166),
.B(n_173),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_169),
.Y(n_416)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_169),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_169),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_172),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_176),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_177),
.Y(n_429)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_178),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.C(n_188),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_185),
.Y(n_252)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_182),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_183),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_185),
.B1(n_198),
.B2(n_202),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_194),
.C(n_198),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_185),
.B(n_194),
.C(n_198),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_186),
.Y(n_554)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g258 ( 
.A1(n_188),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_258)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_192),
.B(n_626),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g439 ( 
.A(n_201),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_202),
.B(n_307),
.C(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_217),
.C(n_219),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_213),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_206),
.B(n_210),
.C(n_213),
.Y(n_262)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_214),
.Y(n_234)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_210),
.B(n_234),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g338 ( 
.A(n_219),
.B(n_339),
.C(n_340),
.Y(n_338)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_221),
.Y(n_580)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g386 ( 
.A(n_222),
.Y(n_386)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

XOR2x1_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_225),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_227),
.Y(n_317)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_230),
.B(n_622),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_259),
.C(n_263),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_232),
.B(n_632),
.Y(n_631)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_235),
.B1(n_255),
.B2(n_258),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_250),
.C(n_253),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_242),
.C(n_246),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_237),
.A2(n_242),
.B1(n_243),
.B2(n_257),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_247),
.C(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_246),
.B(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_252),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g601 ( 
.A(n_256),
.B(n_258),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_259),
.B(n_264),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.C(n_274),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22x1_ASAP7_75t_L g608 ( 
.A1(n_266),
.A2(n_272),
.B1(n_609),
.B2(n_610),
.Y(n_608)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_266),
.Y(n_610)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_271),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_272),
.Y(n_609)
);

XNOR2x1_ASAP7_75t_L g607 ( 
.A(n_274),
.B(n_608),
.Y(n_607)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.C(n_283),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_590)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_282),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_283),
.B(n_590),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_286),
.Y(n_623)
);

XOR2x1_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_305),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B(n_291),
.Y(n_288)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_292),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_324),
.C(n_325),
.Y(n_323)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_330),
.C(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_330),
.C(n_331),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_320),
.C(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.C(n_318),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_328),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_323),
.C(n_326),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_328),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_332),
.B1(n_333),
.B2(n_341),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_338),
.C(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_345),
.B(n_353),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_343),
.B(n_345),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_343),
.B(n_345),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.C(n_349),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_357),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_350),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI21x1_ASAP7_75t_L g644 ( 
.A1(n_353),
.A2(n_645),
.B(n_646),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_354),
.B(n_356),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_619),
.B(n_640),
.Y(n_358)
);

AOI21x1_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_566),
.B(n_617),
.Y(n_359)
);

OAI21x1_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_481),
.B(n_564),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_462),
.C(n_465),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_363),
.B(n_463),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_407),
.Y(n_363)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_364),
.B(n_615),
.C(n_616),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_381),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_365),
.B(n_382),
.C(n_392),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_374),
.C(n_379),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_366),
.B(n_480),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_367),
.A2(n_368),
.B1(n_371),
.B2(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_374),
.A2(n_375),
.B1(n_379),
.B2(n_380),
.Y(n_480)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_392),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_387),
.B(n_391),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_387),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx8_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_391),
.A2(n_592),
.B1(n_593),
.B2(n_594),
.Y(n_591)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_391),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_SL g603 ( 
.A(n_391),
.B(n_589),
.C(n_593),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_394),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_401),
.B1(n_405),
.B2(n_406),
.Y(n_396)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_397),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_397),
.B(n_405),
.C(n_573),
.Y(n_572)
);

INVx3_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_400),
.Y(n_491)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_401),
.Y(n_405)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_404),
.Y(n_578)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_408),
.B(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_441),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_409),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_417),
.C(n_430),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_410),
.B(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g459 ( 
.A(n_411),
.B(n_413),
.C(n_414),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_430),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.C(n_426),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_418),
.B(n_421),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_426),
.Y(n_518)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_435),
.B1(n_436),
.B2(n_440),
.Y(n_430)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_431),
.Y(n_440)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_441),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_457),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g569 ( 
.A(n_442),
.B(n_458),
.C(n_461),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_448),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_444),
.B(n_450),
.C(n_455),
.Y(n_592)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_455),
.B2(n_456),
.Y(n_448)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_449),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_450),
.Y(n_456)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_458),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_459),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_465),
.B(n_565),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_468),
.C(n_478),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_466),
.B(n_562),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_468),
.B(n_479),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.C(n_473),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_469),
.B(n_470),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_510),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.Y(n_473)
);

AO22x1_ASAP7_75t_SL g507 ( 
.A1(n_474),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_507)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_559),
.B(n_563),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_520),
.B(n_558),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_508),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_508),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_502),
.C(n_507),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_485),
.A2(n_486),
.B1(n_531),
.B2(n_533),
.Y(n_530)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_492),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_514),
.C(n_515),
.Y(n_513)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.Y(n_492)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_493),
.Y(n_515)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_497),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_499),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_502),
.A2(n_503),
.B1(n_507),
.B2(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_506),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_506),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_507),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_511),
.B1(n_512),
.B2(n_519),
.Y(n_508)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_513),
.B(n_516),
.C(n_519),
.Y(n_560)
);

XOR2x1_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

AOI21x1_ASAP7_75t_SL g520 ( 
.A1(n_521),
.A2(n_534),
.B(n_557),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_530),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_SL g557 ( 
.A(n_522),
.B(n_530),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_524),
.C(n_527),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_523),
.B(n_542),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_524),
.A2(n_525),
.B1(n_527),
.B2(n_528),
.Y(n_542)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_531),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_535),
.A2(n_543),
.B(n_556),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_541),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_536),
.B(n_541),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_537),
.B(n_540),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_540),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_540),
.B(n_552),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_544),
.A2(n_551),
.B(n_555),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_550),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_550),
.Y(n_555)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_560),
.B(n_561),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_560),
.B(n_561),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_567),
.A2(n_595),
.B(n_611),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_567),
.B(n_595),
.C(n_618),
.Y(n_617)
);

MAJx2_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_585),
.C(n_587),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_568),
.B(n_613),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_569),
.B(n_570),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_569),
.B(n_571),
.C(n_597),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_583),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_574),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_572),
.A2(n_579),
.B(n_582),
.C(n_606),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_575),
.A2(n_579),
.B1(n_581),
.B2(n_582),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_575),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_575),
.B(n_581),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_577),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_579),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_583),
.Y(n_597)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_586),
.B(n_588),
.Y(n_613)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_591),
.Y(n_588)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_592),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_598),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_596),
.B(n_635),
.C(n_636),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_602),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_599),
.Y(n_636)
);

XNOR2x1_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_601),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_602),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_604),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_R g628 ( 
.A(n_603),
.B(n_629),
.C(n_630),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_603),
.B(n_629),
.C(n_630),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_607),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_605),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_607),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_612),
.B(n_614),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_612),
.B(n_614),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_620),
.B(n_633),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_620),
.A2(n_641),
.B(n_642),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_621),
.B(n_624),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_621),
.B(n_624),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_625),
.B(n_628),
.C(n_631),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_625),
.B(n_639),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_631),
.B(n_638),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_634),
.B(n_637),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_634),
.B(n_637),
.Y(n_641)
);

OAI21x1_ASAP7_75t_SL g643 ( 
.A1(n_644),
.A2(n_647),
.B(n_648),
.Y(n_643)
);


endmodule