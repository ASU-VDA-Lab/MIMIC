module real_jpeg_15370_n_13 (n_5, n_4, n_8, n_0, n_12, n_427, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_427;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_0),
.A2(n_14),
.B(n_424),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_0),
.B(n_425),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_1),
.Y(n_425)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_2),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_3),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_3),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_3),
.Y(n_263)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_4),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_4),
.Y(n_309)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_5),
.Y(n_121)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_5),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_5),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_48),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_6),
.A2(n_40),
.B1(n_72),
.B2(n_74),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_6),
.A2(n_40),
.B1(n_311),
.B2(n_314),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_6),
.A2(n_40),
.B1(n_335),
.B2(n_338),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_7),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_8),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_56),
.B1(n_98),
.B2(n_102),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_8),
.A2(n_56),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_8),
.A2(n_56),
.B1(n_321),
.B2(n_325),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

BUFx4f_ASAP7_75t_L g313 ( 
.A(n_10),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_11),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_11),
.B(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_63),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_11),
.A2(n_63),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_11),
.B(n_153),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_11),
.B(n_261),
.C(n_264),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_134),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_133),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_57),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_18),
.B(n_57),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_21),
.B1(n_38),
.B2(n_52),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_19),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_21),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_24),
.Y(n_206)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_29),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_34),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_39),
.A2(n_62),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_46),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_127),
.C(n_131),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_59),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_69),
.C(n_104),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_138),
.C(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_60),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_60),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_60),
.B(n_104),
.C(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_60),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_60),
.A2(n_328),
.B1(n_341),
.B2(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_60),
.A2(n_143),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_60),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_61),
.B(n_165),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_61),
.B(n_165),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_61),
.B(n_165),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_61),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_61),
.B(n_211),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_67),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_63),
.A2(n_147),
.B(n_149),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_63),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_63),
.B(n_107),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_63),
.B(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_66),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_69),
.A2(n_104),
.B1(n_105),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_78),
.B1(n_88),
.B2(n_97),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_71),
.A2(n_79),
.B1(n_146),
.B2(n_153),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_97),
.B(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_79),
.A2(n_146),
.B(n_153),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_101),
.Y(n_228)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_104),
.A2(n_105),
.B1(n_145),
.B2(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_122),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_106),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_107),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_107)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_108),
.Y(n_264)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_108),
.Y(n_305)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_108),
.Y(n_315)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_115),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_118),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_122),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_360)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_157),
.B(n_422),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_154),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_137),
.B(n_154),
.Y(n_423)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_143),
.A2(n_341),
.B1(n_410),
.B2(n_427),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_144),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_145),
.Y(n_406)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_227),
.A3(n_229),
.B1(n_232),
.B2(n_238),
.Y(n_226)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_398),
.B(n_419),
.Y(n_157)
);

AO221x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_293),
.B1(n_390),
.B2(n_396),
.C(n_397),
.Y(n_158)
);

AO21x2_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_243),
.B(n_292),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_219),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_161),
.B(n_219),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_209),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_184),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_163),
.B(n_184),
.C(n_209),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_164),
.A2(n_211),
.B1(n_217),
.B2(n_218),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_164),
.A2(n_217),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_164),
.A2(n_218),
.B(n_248),
.C(n_250),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_164),
.A2(n_360),
.B(n_361),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_164),
.B(n_360),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_165),
.B(n_211),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_168),
.B1(n_185),
.B2(n_208),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_167),
.B(n_226),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_167),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_167),
.B(n_218),
.C(n_257),
.Y(n_287)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_168),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_168),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_168),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_168),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_168),
.B(n_185),
.Y(n_371)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_179),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_170),
.A2(n_302),
.B1(n_310),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_177),
.Y(n_277)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_179),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_181),
.Y(n_318)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_181),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_183),
.Y(n_281)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_191),
.B(n_199),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_202),
.B(n_207),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_210),
.A2(n_248),
.B1(n_249),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_218),
.B1(n_224),
.B2(n_225),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_218),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_211),
.A2(n_218),
.B1(n_259),
.B2(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_211),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_211),
.B(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_211),
.A2(n_218),
.B1(n_301),
.B2(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_211),
.A2(n_218),
.B1(n_345),
.B2(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_212),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.C(n_242),
.Y(n_219)
);

XOR2x2_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

OAI21x1_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_251),
.B(n_291),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AND3x1_ASAP7_75t_L g383 ( 
.A(n_250),
.B(n_349),
.C(n_384),
.Y(n_383)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_286),
.B(n_290),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_267),
.B(n_285),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_258),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_282),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_288),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_374),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_362),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_295),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_350),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_296),
.B(n_350),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_327),
.C(n_342),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_297),
.B(n_327),
.Y(n_373)
);

OAI22x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_326),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_298),
.B(n_371),
.Y(n_377)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_299),
.A2(n_344),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_300),
.A2(n_343),
.B(n_347),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_310),
.B1(n_316),
.B2(n_319),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_330),
.B1(n_331),
.B2(n_341),
.Y(n_327)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_328),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_R g355 ( 
.A(n_328),
.B(n_331),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_373),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B(n_347),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_343),
.A2(n_347),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_358),
.B2(n_359),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_354),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_413),
.C(n_414),
.Y(n_412)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_361),
.A2(n_402),
.B1(n_403),
.B2(n_407),
.Y(n_401)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_372),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_372),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.C(n_370),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_368),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_386),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_385),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_385),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_380),
.C(n_382),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_388),
.Y(n_393)
);

A2O1A1Ixp33_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_393),
.B(n_394),
.C(n_395),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_415),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_412),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_412),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_408),
.B1(n_409),
.B2(n_411),
.Y(n_400)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_401),
.Y(n_411)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_407),
.C(n_408),
.Y(n_418)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_415),
.A2(n_420),
.B(n_421),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_418),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);


endmodule