module fake_jpeg_23455_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_43),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_45),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_7),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_51),
.A2(n_53),
.B1(n_59),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_20),
.B1(n_27),
.B2(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_27),
.B1(n_33),
.B2(n_26),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_41),
.B1(n_43),
.B2(n_38),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_33),
.B1(n_26),
.B2(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_33),
.B1(n_26),
.B2(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_32),
.B1(n_17),
.B2(n_28),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_28),
.B1(n_24),
.B2(n_17),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_34),
.B1(n_22),
.B2(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_43),
.B1(n_31),
.B2(n_35),
.Y(n_79)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_30),
.B1(n_16),
.B2(n_23),
.Y(n_128)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_85),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_35),
.B1(n_30),
.B2(n_19),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_19),
.B(n_30),
.C(n_44),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_35),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_37),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_104),
.Y(n_124)
);

NAND2x1p5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_37),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_60),
.B(n_16),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_90),
.B(n_107),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_16),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_102),
.Y(n_142)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_37),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_109),
.B1(n_60),
.B2(n_66),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_35),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_74),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_0),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_12),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_121),
.Y(n_161)
);

XOR2x2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_62),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_99),
.C(n_77),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_123),
.B1(n_102),
.B2(n_105),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_15),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_49),
.B1(n_44),
.B2(n_19),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_128),
.B1(n_92),
.B2(n_93),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_30),
.B1(n_23),
.B2(n_16),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_130),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_60),
.B1(n_40),
.B2(n_56),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_137),
.B(n_81),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_66),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_16),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_88),
.Y(n_152)
);

BUFx8_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_141),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_146),
.Y(n_179)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_153),
.B(n_138),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_164),
.B1(n_122),
.B2(n_128),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_159),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_154),
.B(n_155),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_158),
.B1(n_167),
.B2(n_175),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_165),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_76),
.B1(n_96),
.B2(n_110),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_112),
.C(n_111),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_137),
.C(n_132),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_126),
.B1(n_117),
.B2(n_120),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_168),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_76),
.B1(n_96),
.B2(n_97),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_130),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_11),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_12),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_125),
.B(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_119),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_200),
.C(n_146),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_116),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_208),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_118),
.B1(n_121),
.B2(n_124),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_198),
.B1(n_13),
.B2(n_15),
.Y(n_234)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_151),
.A2(n_124),
.B1(n_138),
.B2(n_115),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_159),
.C(n_157),
.Y(n_200)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_154),
.B1(n_166),
.B2(n_161),
.C(n_162),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_115),
.B(n_2),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_1),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_140),
.B(n_139),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_140),
.B(n_139),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_210),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_156),
.B(n_169),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_212),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_168),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_174),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_226),
.C(n_235),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_217),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_144),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_220),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_189),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_209),
.Y(n_220)
);

AO22x1_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_172),
.B1(n_161),
.B2(n_145),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_221),
.A2(n_227),
.B(n_1),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_173),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_222),
.B(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_230),
.B(n_236),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_176),
.C(n_131),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_131),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_237),
.B1(n_199),
.B2(n_180),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_182),
.B1(n_197),
.B2(n_195),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_95),
.C(n_108),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_185),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_245),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_185),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_257),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_192),
.B1(n_190),
.B2(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_202),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_201),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_255),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_186),
.B1(n_193),
.B2(n_178),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_196),
.C(n_95),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_223),
.B(n_188),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_229),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_232),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_238),
.B1(n_230),
.B2(n_236),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_268),
.A2(n_277),
.B1(n_244),
.B2(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_231),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_269),
.B(n_271),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_278),
.Y(n_294)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_228),
.B(n_238),
.C(n_220),
.D(n_216),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_241),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_218),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_213),
.B1(n_214),
.B2(n_226),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_242),
.B(n_222),
.Y(n_278)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_292),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_240),
.C(n_255),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_286),
.C(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_259),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_240),
.C(n_250),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_234),
.B1(n_227),
.B2(n_239),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_273),
.B1(n_263),
.B2(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_264),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_290),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_246),
.Y(n_292)
);

OAI21x1_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_283),
.B(n_281),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_296),
.A2(n_302),
.B1(n_243),
.B2(n_14),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_284),
.C(n_286),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_265),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_268),
.B(n_280),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_290),
.B(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_282),
.B(n_251),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_232),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_5),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_309),
.A2(n_314),
.B1(n_315),
.B2(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_316),
.C(n_301),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_287),
.B1(n_265),
.B2(n_292),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_2),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_324),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_305),
.B(n_302),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_298),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_299),
.C(n_304),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_316),
.B(n_315),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_320),
.B(n_4),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_3),
.A3(n_4),
.B1(n_308),
.B2(n_318),
.C1(n_325),
.C2(n_321),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_322),
.B(n_4),
.C(n_3),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_330),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_331),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_329),
.C(n_327),
.Y(n_334)
);


endmodule