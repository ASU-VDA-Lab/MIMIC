module fake_ariane_722_n_7869 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_7869);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_7869;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_7805;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_6293;
wire n_2482;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_4260;
wire n_903;
wire n_7626;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_7368;
wire n_1690;
wire n_2807;
wire n_6664;
wire n_7562;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_6891;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_6539;
wire n_4824;
wire n_7467;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_7526;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_786;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_863;
wire n_6992;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_6681;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_7507;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_2382;
wire n_1213;
wire n_7379;
wire n_7441;
wire n_780;
wire n_5292;
wire n_1918;
wire n_7438;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_5843;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_1386;
wire n_6236;
wire n_7104;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_5984;
wire n_5204;
wire n_6705;
wire n_6724;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_7840;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6261;
wire n_6659;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3891;
wire n_3372;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_7583;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_2954;
wire n_4438;
wire n_6538;
wire n_974;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_5708;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_3147;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_1247;
wire n_6860;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_6382;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_6615;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_720;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_5149;
wire n_5280;
wire n_3054;
wire n_4970;
wire n_1163;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_5985;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_7868;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_7176;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_1104;
wire n_986;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1498;
wire n_1188;
wire n_7527;
wire n_4856;
wire n_2618;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_6482;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_951;
wire n_7546;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_7481;
wire n_1714;
wire n_4429;
wire n_1044;
wire n_5435;
wire n_6484;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_7605;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_6639;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_6204;
wire n_906;
wire n_1330;
wire n_2295;
wire n_5225;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_7600;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_6946;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_7660;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_6840;
wire n_6645;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_7455;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_7509;
wire n_6205;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_7497;
wire n_7315;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_6706;
wire n_7431;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_1291;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_7505;
wire n_3921;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_775;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_7573;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_7498;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6395;
wire n_3497;
wire n_6403;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_7240;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_1056;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_6541;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_4733;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_7382;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_6744;
wire n_3645;
wire n_793;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_6116;
wire n_3550;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_7671;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7821;
wire n_7620;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_1775;
wire n_908;
wire n_1036;
wire n_7109;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_6716;
wire n_3565;
wire n_6905;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_7817;
wire n_6413;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_1261;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_857;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_2324;
wire n_840;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_7140;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_3303;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_6668;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_7698;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_7650;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_4548;
wire n_7819;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_3707;
wire n_3895;
wire n_768;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6963;
wire n_6951;
wire n_1581;
wire n_946;
wire n_3058;
wire n_757;
wire n_2047;
wire n_5355;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_5915;
wire n_7276;
wire n_6379;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_4716;
wire n_3722;
wire n_1001;
wire n_1313;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_803;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5966;
wire n_4591;
wire n_5569;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_7160;
wire n_7324;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_6055;
wire n_7161;
wire n_1808;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_7837;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_7676;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_7644;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_6607;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_829;
wire n_4814;
wire n_6178;
wire n_6677;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_7550;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_7804;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_1276;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_7826;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_3728;
wire n_2722;
wire n_6596;
wire n_5107;
wire n_7165;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_772;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_3234;
wire n_1351;
wire n_2216;
wire n_2426;
wire n_6947;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7675;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_7774;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_2224;
wire n_1226;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_3046;
wire n_2293;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_3014;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_7764;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_7520;
wire n_5314;
wire n_7616;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_6572;
wire n_3981;
wire n_7271;
wire n_2681;
wire n_7222;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_6387;
wire n_4201;
wire n_6470;
wire n_7206;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_7854;
wire n_926;
wire n_2296;
wire n_5735;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_3377;
wire n_6722;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_7436;
wire n_7020;
wire n_5935;
wire n_6696;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_5488;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1614;
wire n_1377;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_7465;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_729;
wire n_6222;
wire n_2218;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_6587;
wire n_6688;
wire n_6505;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_7449;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_3216;
wire n_3568;
wire n_2555;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_7479;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_6547;
wire n_7177;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_6478;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_7818;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_3459;
wire n_2576;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_7862;
wire n_3735;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_6999;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_6440;
wire n_4977;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_3408;
wire n_2884;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_6464;
wire n_5129;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_6850;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_7743;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_6972;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_3317;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_4251;
wire n_2393;
wire n_5266;
wire n_2143;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_7035;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_6258;
wire n_1288;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_7699;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_5911;
wire n_7340;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_914;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_7207;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_7633;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_2592;
wire n_3490;
wire n_7280;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_4241;
wire n_1622;
wire n_3113;
wire n_2751;
wire n_4183;
wire n_7768;
wire n_1968;
wire n_918;
wire n_5645;
wire n_5020;
wire n_6455;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_2150;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_1262;
wire n_792;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_7101;
wire n_1204;
wire n_7843;
wire n_2428;
wire n_994;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_6993;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7310;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_6105;
wire n_826;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_7609;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_7282;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_6331;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_7820;
wire n_816;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_1629;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_6450;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_1236;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_7723;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_4258;
wire n_5756;
wire n_7693;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_7682;
wire n_7300;
wire n_939;
wire n_1410;
wire n_2297;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_7798;
wire n_4767;
wire n_4569;
wire n_948;
wire n_6528;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_5039;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_4265;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_1583;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_1264;
wire n_6530;
wire n_6602;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_1752;
wire n_2361;
wire n_3030;
wire n_4538;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_7336;
wire n_5932;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_7493;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_5823;
wire n_2423;
wire n_2208;
wire n_1421;
wire n_5422;
wire n_5944;
wire n_6989;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_1069;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_7273;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_6758;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_7601;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_5294;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1187;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_7617;
wire n_4575;
wire n_945;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_7700;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_4968;
wire n_7801;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_5290;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_4176;
wire n_7556;
wire n_4124;
wire n_4431;
wire n_3347;
wire n_1404;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_6691;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5718;
wire n_1461;
wire n_5503;
wire n_7208;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_5610;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_1253;
wire n_1468;
wire n_762;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_6533;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_7483;
wire n_5710;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_5333;
wire n_1083;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_5109;
wire n_1071;
wire n_712;
wire n_909;
wire n_6713;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_5862;
wire n_7477;
wire n_1914;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_7714;
wire n_6415;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6513;
wire n_6392;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_7710;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_5132;
wire n_3498;
wire n_1173;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_4728;
wire n_7171;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_7501;
wire n_6432;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_3983;
wire n_703;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_6957;
wire n_5074;
wire n_3939;
wire n_3788;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_6694;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_3139;
wire n_5681;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_7621;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_7572;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_6662;
wire n_7494;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_6200;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_5657;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_6956;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_6701;
wire n_2594;
wire n_5298;
wire n_1239;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_6362;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_7126;
wire n_5867;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_4436;
wire n_5822;
wire n_5786;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_4385;
wire n_7779;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_1786;
wire n_6309;
wire n_3732;
wire n_1804;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_1318;
wire n_1769;
wire n_1632;
wire n_7349;
wire n_1929;
wire n_4319;
wire n_6585;
wire n_7786;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_7579;
wire n_7122;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_7624;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_5475;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_5315;
wire n_3708;
wire n_2633;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_6685;
wire n_3390;
wire n_756;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_3140;
wire n_2320;
wire n_4082;
wire n_979;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_897;
wire n_7347;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_885;
wire n_3955;
wire n_1659;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_3336;
wire n_7739;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_6549;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_7456;
wire n_7369;
wire n_1472;
wire n_1050;
wire n_7548;
wire n_2578;
wire n_1201;
wire n_7598;
wire n_2475;
wire n_1185;
wire n_7250;
wire n_7823;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_6923;
wire n_7649;
wire n_843;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_7844;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_7371;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_7463;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5755;
wire n_5700;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_6184;
wire n_1767;
wire n_4138;
wire n_3131;
wire n_1040;
wire n_7083;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_7683;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_7330;
wire n_6007;
wire n_6734;
wire n_6535;
wire n_1772;
wire n_6879;
wire n_3106;
wire n_1311;
wire n_6208;
wire n_7190;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_7042;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_3178;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7787;
wire n_7836;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_6764;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_969;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_6569;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_7103;
wire n_6605;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_6832;
wire n_5980;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_7771;
wire n_4255;
wire n_2758;
wire n_6544;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_6289;
wire n_6651;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_7706;
wire n_7813;
wire n_2420;
wire n_7643;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_835;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_839;
wire n_1754;
wire n_7236;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_6786;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7519;
wire n_7802;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_2933;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_6945;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_977;
wire n_2339;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_6175;
wire n_6445;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_6499;
wire n_1982;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_3504;
wire n_2587;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_3112;
wire n_954;
wire n_2562;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_7646;
wire n_3779;
wire n_6982;
wire n_1063;
wire n_7291;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_7017;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_7861;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_7554;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_4014;
wire n_3547;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_6851;
wire n_6621;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_7420;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_7244;
wire n_1463;
wire n_4626;
wire n_7625;
wire n_4997;
wire n_5065;
wire n_6806;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_7154;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_7068;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_4549;
wire n_1073;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_4734;
wire n_6675;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_7384;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_1544;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_7559;
wire n_7576;
wire n_6988;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_6280;
wire n_3280;
wire n_1590;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_7264;
wire n_7842;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_7492;
wire n_804;
wire n_6649;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_6431;
wire n_4223;
wire n_3250;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_824;
wire n_5659;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_7793;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_7746;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_6473;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_836;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_7703;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_7665;
wire n_5262;
wire n_7677;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_3699;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_7203;
wire n_7797;
wire n_1826;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_7111;
wire n_2801;
wire n_4334;
wire n_1177;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_6617;
wire n_7725;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_6217;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_6777;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_6370;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_3009;
wire n_777;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_7530;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_6465;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_1222;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_4463;
wire n_5357;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_7591;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_3953;
wire n_4400;
wire n_7502;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_7065;
wire n_1466;
wire n_6177;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_7367;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1037;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_4035;
wire n_6952;
wire n_1480;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_5577;
wire n_876;
wire n_5872;
wire n_6692;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_3694;
wire n_6854;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_7728;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_7181;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_748;
wire n_7089;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_5868;
wire n_6417;
wire n_7145;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_7803;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_7622;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_6831;
wire n_1773;
wire n_4544;
wire n_3175;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_7564;
wire n_5863;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_6152;
wire n_5734;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_7262;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_763;
wire n_6301;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_6282;
wire n_4934;
wire n_7686;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_6737;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_6448;
wire n_5186;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_7077;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_7663;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_7214;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_3989;
wire n_7652;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_7086;
wire n_5689;
wire n_7732;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_7038;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_7593;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_7757;
wire n_1093;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_6601;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_7439;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_7744;
wire n_3898;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_4168;
wire n_1369;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_7480;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_7380;
wire n_2839;
wire n_3237;
wire n_7708;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_7376;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_6409;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_7657;
wire n_6388;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_6679;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_937;
wire n_1631;
wire n_7602;
wire n_6566;
wire n_1794;
wire n_5696;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_7582;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_7555;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

INVx2_ASAP7_75t_L g700 ( 
.A(n_437),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_404),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_209),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_491),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_157),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_145),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_536),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_144),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_636),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_695),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_18),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_674),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_463),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_468),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_253),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_606),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_630),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_169),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_473),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_255),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_338),
.Y(n_720)
);

BUFx10_ASAP7_75t_L g721 ( 
.A(n_459),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_17),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_272),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_376),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_482),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_214),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_435),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_97),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_214),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_381),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_169),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_432),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_183),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_436),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_454),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_471),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_649),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_372),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_436),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_699),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_219),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_131),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_528),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_65),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_698),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_100),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_289),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_185),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_261),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_566),
.Y(n_750)
);

CKINVDCx14_ASAP7_75t_R g751 ( 
.A(n_303),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_397),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_124),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_648),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_524),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_244),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_572),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_6),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_389),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_391),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_307),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_3),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_177),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_546),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_59),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_189),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_321),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_293),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_447),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_424),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_45),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_505),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_522),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_592),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_362),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_244),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_130),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_683),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_520),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_123),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_178),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_525),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_690),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_470),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_572),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_555),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_10),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_554),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_531),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_114),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_490),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_538),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_43),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_363),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_232),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_77),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_207),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_93),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_1),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_502),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_225),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_383),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_362),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_318),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_171),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_599),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_646),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_14),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_219),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_452),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_130),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_201),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_43),
.Y(n_813)
);

INVxp33_ASAP7_75t_L g814 ( 
.A(n_359),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_263),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_69),
.Y(n_816)
);

CKINVDCx16_ASAP7_75t_R g817 ( 
.A(n_198),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_587),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_157),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_25),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_227),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_685),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_496),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_613),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_536),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_577),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_611),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_42),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_116),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_649),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_321),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_129),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_256),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_225),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_58),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_481),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_311),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_615),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_349),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_506),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_554),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_66),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_182),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_43),
.Y(n_844)
);

INVxp33_ASAP7_75t_R g845 ( 
.A(n_117),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_93),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_662),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_152),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_136),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_122),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_28),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_142),
.Y(n_852)
);

BUFx10_ASAP7_75t_L g853 ( 
.A(n_605),
.Y(n_853)
);

CKINVDCx16_ASAP7_75t_R g854 ( 
.A(n_36),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_496),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_278),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_468),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_279),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_79),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_121),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_314),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_617),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_524),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_41),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_46),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_566),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_469),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_287),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_240),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_249),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_340),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_163),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_414),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_279),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_197),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_173),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_82),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_291),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_659),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_89),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_137),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_50),
.Y(n_882)
);

BUFx10_ASAP7_75t_L g883 ( 
.A(n_251),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_114),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_553),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_477),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_315),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_328),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_413),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_418),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_641),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_304),
.Y(n_892)
);

CKINVDCx16_ASAP7_75t_R g893 ( 
.A(n_95),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_323),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_83),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_124),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_316),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_377),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_491),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_331),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_323),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_109),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_542),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_26),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_343),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_293),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_503),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_226),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_5),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_50),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_480),
.Y(n_911)
);

CKINVDCx14_ASAP7_75t_R g912 ( 
.A(n_307),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_104),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_334),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_595),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_192),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_495),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_328),
.Y(n_918)
);

BUFx10_ASAP7_75t_L g919 ( 
.A(n_665),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_666),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_358),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_590),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_91),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_402),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_77),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_232),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_87),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_281),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_343),
.Y(n_929)
);

BUFx5_ASAP7_75t_L g930 ( 
.A(n_607),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_189),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_23),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_440),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_680),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_622),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_659),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_634),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_25),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_51),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_617),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_503),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_234),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_2),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_132),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_247),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_547),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_74),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_325),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_211),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_257),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_68),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_1),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_650),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_32),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_52),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_118),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_634),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_458),
.Y(n_958)
);

BUFx8_ASAP7_75t_SL g959 ( 
.A(n_633),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_228),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_567),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_430),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_145),
.Y(n_963)
);

CKINVDCx16_ASAP7_75t_R g964 ( 
.A(n_467),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_273),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_324),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_563),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_411),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_680),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_74),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_416),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_74),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_332),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_106),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_180),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_181),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_266),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_466),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_457),
.Y(n_979)
);

CKINVDCx14_ASAP7_75t_R g980 ( 
.A(n_687),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_287),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_515),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_608),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_305),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_10),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_691),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_693),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_230),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_151),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_520),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_562),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_661),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_588),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_563),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_191),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_208),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_585),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_448),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_208),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_384),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_688),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_466),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_619),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_592),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_446),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_247),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_187),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_429),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_669),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_387),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_206),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_616),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_565),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_319),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_155),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_693),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_682),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_670),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_573),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_327),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_559),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_523),
.Y(n_1022)
);

BUFx5_ASAP7_75t_L g1023 ( 
.A(n_47),
.Y(n_1023)
);

CKINVDCx16_ASAP7_75t_R g1024 ( 
.A(n_233),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_696),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_256),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_694),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_697),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_300),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_286),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_630),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_129),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_365),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_64),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_61),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_591),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_151),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_47),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_533),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_176),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_75),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_517),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_292),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_477),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_472),
.Y(n_1046)
);

CKINVDCx16_ASAP7_75t_R g1047 ( 
.A(n_637),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_376),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_340),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_254),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_262),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_694),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_582),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_216),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_3),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_488),
.Y(n_1056)
);

BUFx10_ASAP7_75t_L g1057 ( 
.A(n_148),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_211),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_570),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_416),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_268),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_277),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_227),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_613),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_689),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_40),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_167),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_124),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_346),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_78),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_506),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_502),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_238),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_457),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_155),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_158),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_254),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_186),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_257),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_622),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_370),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_146),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_699),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_108),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_361),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_558),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_308),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_89),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_548),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_368),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_499),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_69),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_623),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_460),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_460),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_68),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_290),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_534),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_414),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_152),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_253),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_107),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_96),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_681),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_61),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_295),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_276),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_697),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_652),
.Y(n_1109)
);

CKINVDCx14_ASAP7_75t_R g1110 ( 
.A(n_115),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_223),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_493),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_672),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_676),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_437),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_198),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_170),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_200),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_549),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_108),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_51),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_653),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_117),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_633),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_367),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_188),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_522),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_103),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_403),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_448),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_243),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_428),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_65),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_369),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_281),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_581),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_36),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_240),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_615),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_40),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_170),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_299),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_361),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_678),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_367),
.Y(n_1145)
);

BUFx8_ASAP7_75t_SL g1146 ( 
.A(n_378),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_194),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_631),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_586),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_517),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_640),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_11),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_45),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_408),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_216),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_2),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_178),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_262),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_669),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_29),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_654),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_310),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_684),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_148),
.Y(n_1164)
);

CKINVDCx16_ASAP7_75t_R g1165 ( 
.A(n_87),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_97),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_213),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_346),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_338),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_569),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_44),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_653),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_298),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_162),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_684),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_350),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_310),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_201),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_92),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_382),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_392),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_429),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_316),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_476),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_306),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_623),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_692),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_228),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_272),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_260),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_492),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_251),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_96),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_210),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_618),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_204),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_501),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_386),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_467),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_546),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_176),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_543),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_175),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_422),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_329),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_103),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_73),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_161),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_81),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_8),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_19),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_70),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_664),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_463),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_95),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_543),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_397),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_442),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_41),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_675),
.Y(n_1220)
);

BUFx5_ASAP7_75t_L g1221 ( 
.A(n_261),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_686),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_415),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_604),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_347),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_60),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_561),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_420),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_465),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_33),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_352),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_424),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_504),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_435),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_428),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_681),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_620),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_548),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_660),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_117),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_159),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_65),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1023),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1023),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_751),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_751),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_912),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1023),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1023),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1023),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1023),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1023),
.Y(n_1252)
);

CKINVDCx16_ASAP7_75t_R g1253 ( 
.A(n_1110),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_912),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_980),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_864),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_864),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_715),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_980),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_864),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_927),
.Y(n_1261)
);

INVxp33_ASAP7_75t_SL g1262 ( 
.A(n_821),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_927),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_927),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1156),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1156),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_959),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_790),
.B(n_0),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_811),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1156),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1219),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1023),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_1219),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1219),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_713),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_713),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_713),
.Y(n_1277)
);

INVxp33_ASAP7_75t_L g1278 ( 
.A(n_821),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_959),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_791),
.Y(n_1280)
);

CKINVDCx14_ASAP7_75t_R g1281 ( 
.A(n_1110),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_767),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_767),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1146),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_767),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_778),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_778),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_1146),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_778),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1023),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_819),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1023),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1023),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_791),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_819),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_819),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_930),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_930),
.B(n_0),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_817),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_817),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_930),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_930),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_930),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_823),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_930),
.Y(n_1305)
);

NOR2xp67_ASAP7_75t_L g1306 ( 
.A(n_790),
.B(n_0),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_930),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_823),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_930),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_964),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_930),
.Y(n_1311)
);

INVxp33_ASAP7_75t_L g1312 ( 
.A(n_982),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_930),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_930),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_715),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_709),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1221),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1221),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1221),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1221),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_882),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_709),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1221),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_964),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1221),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1221),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1024),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1221),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_727),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1221),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1024),
.Y(n_1331)
);

INVx4_ASAP7_75t_R g1332 ( 
.A(n_746),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1221),
.Y(n_1333)
);

INVxp33_ASAP7_75t_L g1334 ( 
.A(n_982),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_882),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_715),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1047),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_746),
.Y(n_1338)
);

INVxp33_ASAP7_75t_SL g1339 ( 
.A(n_1170),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_882),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_882),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_870),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1047),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_811),
.Y(n_1344)
);

CKINVDCx14_ASAP7_75t_R g1345 ( 
.A(n_799),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_882),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_882),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_882),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_814),
.B(n_2),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1093),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1207),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1207),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_1207),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1207),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1207),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_811),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1207),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1207),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_854),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1093),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1033),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1033),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1033),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1153),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1153),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1153),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1210),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1216),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1210),
.Y(n_1369)
);

INVxp33_ASAP7_75t_L g1370 ( 
.A(n_1170),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1210),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_791),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_700),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_791),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_727),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_700),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1216),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_700),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_717),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_717),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_717),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_779),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_791),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_854),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_791),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1068),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_779),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_779),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_870),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_804),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_804),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_893),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_804),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_809),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_809),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_809),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_891),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_891),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_791),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1068),
.B(n_3),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_870),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_891),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_940),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_940),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_940),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_958),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_701),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_825),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_958),
.Y(n_1409)
);

INVxp33_ASAP7_75t_L g1410 ( 
.A(n_1164),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_704),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_958),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_893),
.Y(n_1413)
);

CKINVDCx16_ASAP7_75t_R g1414 ( 
.A(n_1165),
.Y(n_1414)
);

CKINVDCx14_ASAP7_75t_R g1415 ( 
.A(n_799),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_960),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_810),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_825),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_825),
.Y(n_1419)
);

INVxp67_ASAP7_75t_L g1420 ( 
.A(n_1031),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_810),
.Y(n_1421)
);

NOR2xp67_ASAP7_75t_L g1422 ( 
.A(n_790),
.B(n_4),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1038),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_810),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1068),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1038),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1038),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_706),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_708),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_711),
.Y(n_1430)
);

CKINVDCx14_ASAP7_75t_R g1431 ( 
.A(n_799),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_810),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_810),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_810),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_712),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_865),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_716),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1052),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1052),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1052),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1178),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1178),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1178),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1184),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1184),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1184),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_718),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1217),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_810),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1217),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1217),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_740),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1220),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1220),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_841),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1220),
.Y(n_1456)
);

INVxp67_ASAP7_75t_SL g1457 ( 
.A(n_865),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1233),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_740),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1233),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1233),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_865),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_841),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_723),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_960),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1031),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_729),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_932),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_747),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_841),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_939),
.Y(n_1471)
);

INVxp33_ASAP7_75t_SL g1472 ( 
.A(n_1164),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_939),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_939),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1120),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1120),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1120),
.Y(n_1477)
);

CKINVDCx16_ASAP7_75t_R g1478 ( 
.A(n_1165),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1140),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1140),
.Y(n_1480)
);

CKINVDCx16_ASAP7_75t_R g1481 ( 
.A(n_799),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1140),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1031),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1056),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_841),
.Y(n_1485)
);

CKINVDCx16_ASAP7_75t_R g1486 ( 
.A(n_799),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1056),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_841),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1103),
.B(n_4),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1056),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1060),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1060),
.Y(n_1492)
);

BUFx5_ASAP7_75t_L g1493 ( 
.A(n_728),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1060),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_747),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_730),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1122),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_841),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_841),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1122),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_750),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_750),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1122),
.Y(n_1503)
);

CKINVDCx16_ASAP7_75t_R g1504 ( 
.A(n_1057),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1169),
.Y(n_1505)
);

INVxp33_ASAP7_75t_SL g1506 ( 
.A(n_1169),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_862),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_862),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_728),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1169),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_731),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1057),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_732),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1103),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1103),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_734),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_741),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_753),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_733),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_752),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_862),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_745),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_748),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_733),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_733),
.Y(n_1525)
);

INVxp67_ASAP7_75t_SL g1526 ( 
.A(n_744),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_759),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_784),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_752),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_784),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_862),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_784),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_753),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_863),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_863),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_863),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_760),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_771),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1049),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1049),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_761),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1049),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_862),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1104),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1104),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1104),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1118),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1118),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1118),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_862),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_763),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1134),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1134),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1134),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1190),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_744),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_862),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1190),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1190),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1200),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1200),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_764),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1200),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_787),
.B(n_4),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_787),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_808),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_771),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_808),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_820),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_769),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_820),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_828),
.Y(n_1572)
);

CKINVDCx16_ASAP7_75t_R g1573 ( 
.A(n_1057),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_776),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_995),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_828),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_776),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_832),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_814),
.B(n_5),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_832),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_813),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_849),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_849),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_851),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_772),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_851),
.Y(n_1586)
);

CKINVDCx16_ASAP7_75t_R g1587 ( 
.A(n_1057),
.Y(n_1587)
);

XOR2xp5_ASAP7_75t_L g1588 ( 
.A(n_707),
.B(n_5),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_860),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_995),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_860),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_781),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_909),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_909),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_774),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_782),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_910),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_813),
.Y(n_1598)
);

CKINVDCx14_ASAP7_75t_R g1599 ( 
.A(n_1057),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_910),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_913),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_913),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_947),
.Y(n_1603)
);

CKINVDCx16_ASAP7_75t_R g1604 ( 
.A(n_721),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_781),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_947),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_995),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_951),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_951),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_952),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_995),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_952),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_783),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_807),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_920),
.B(n_6),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_785),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_956),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_995),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_956),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_L g1620 ( 
.A(n_920),
.B(n_6),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_963),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_788),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_963),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_807),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_985),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_985),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1029),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1029),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1042),
.Y(n_1629)
);

BUFx2_ASAP7_75t_SL g1630 ( 
.A(n_721),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_789),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_960),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_795),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_968),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_826),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_968),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_968),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1003),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_995),
.Y(n_1639)
);

CKINVDCx16_ASAP7_75t_R g1640 ( 
.A(n_721),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_995),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1003),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1003),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1009),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_816),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1009),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_816),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_801),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1009),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1130),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1130),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1130),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1186),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1030),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_805),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_812),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1186),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1186),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1030),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1205),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1205),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_835),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1205),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1030),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_848),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1208),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1208),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_855),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1208),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_856),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1237),
.Y(n_1671)
);

INVxp33_ASAP7_75t_L g1672 ( 
.A(n_702),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1237),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1237),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1030),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1054),
.B(n_7),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1042),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1088),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_857),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1088),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_826),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1096),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1096),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_835),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_858),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1105),
.B(n_7),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_932),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1436),
.B(n_1030),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1321),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1408),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1338),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1345),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1415),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1408),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1512),
.B(n_721),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1462),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1468),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1687),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1630),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1316),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1322),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1431),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1599),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1353),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1471),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1512),
.B(n_721),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1473),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1474),
.Y(n_1708)
);

CKINVDCx16_ASAP7_75t_R g1709 ( 
.A(n_1481),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1329),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1384),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1475),
.Y(n_1712)
);

NOR2xp67_ASAP7_75t_L g1713 ( 
.A(n_1533),
.B(n_1054),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1476),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1477),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1375),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1355),
.Y(n_1717)
);

CKINVDCx20_ASAP7_75t_R g1718 ( 
.A(n_1452),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1354),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1480),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1482),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1519),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1269),
.B(n_955),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1414),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1457),
.B(n_1030),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1355),
.Y(n_1726)
);

INVxp33_ASAP7_75t_SL g1727 ( 
.A(n_1279),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1459),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1524),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1479),
.B(n_1256),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1525),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1478),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1528),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1530),
.Y(n_1734)
);

INVxp33_ASAP7_75t_SL g1735 ( 
.A(n_1279),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1532),
.Y(n_1736)
);

CKINVDCx20_ASAP7_75t_R g1737 ( 
.A(n_1469),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1354),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1267),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1288),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1372),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1269),
.B(n_1344),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1534),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1535),
.Y(n_1744)
);

NOR2xp67_ASAP7_75t_L g1745 ( 
.A(n_1598),
.B(n_1086),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1630),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1536),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1538),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1495),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1501),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1246),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1246),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1297),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1299),
.Y(n_1754)
);

CKINVDCx16_ASAP7_75t_R g1755 ( 
.A(n_1486),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1372),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1539),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1538),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1540),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1299),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1542),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1544),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1545),
.Y(n_1763)
);

CKINVDCx16_ASAP7_75t_R g1764 ( 
.A(n_1504),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1247),
.Y(n_1765)
);

XNOR2x2_ASAP7_75t_R g1766 ( 
.A(n_1588),
.B(n_845),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1374),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1247),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1255),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1502),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1546),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1547),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1520),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1255),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1548),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1259),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1493),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1374),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1493),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1300),
.Y(n_1780)
);

CKINVDCx16_ASAP7_75t_R g1781 ( 
.A(n_1573),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1297),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1280),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1493),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1493),
.Y(n_1785)
);

CKINVDCx16_ASAP7_75t_R g1786 ( 
.A(n_1587),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1493),
.Y(n_1787)
);

INVxp33_ASAP7_75t_SL g1788 ( 
.A(n_1259),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1549),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1552),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1553),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_R g1792 ( 
.A(n_1281),
.B(n_861),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1554),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1506),
.B(n_794),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1407),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1407),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1506),
.B(n_794),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1555),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1558),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1411),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1559),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1560),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1319),
.Y(n_1803)
);

INVxp33_ASAP7_75t_SL g1804 ( 
.A(n_1284),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1411),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1428),
.Y(n_1806)
);

CKINVDCx20_ASAP7_75t_R g1807 ( 
.A(n_1529),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1300),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1561),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1428),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_1574),
.Y(n_1811)
);

NOR2xp67_ASAP7_75t_L g1812 ( 
.A(n_1645),
.B(n_1647),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1563),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1275),
.Y(n_1814)
);

CKINVDCx16_ASAP7_75t_R g1815 ( 
.A(n_1604),
.Y(n_1815)
);

CKINVDCx20_ASAP7_75t_R g1816 ( 
.A(n_1577),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1276),
.Y(n_1817)
);

NOR2xp67_ASAP7_75t_L g1818 ( 
.A(n_1429),
.B(n_1086),
.Y(n_1818)
);

CKINVDCx20_ASAP7_75t_R g1819 ( 
.A(n_1592),
.Y(n_1819)
);

CKINVDCx20_ASAP7_75t_R g1820 ( 
.A(n_1605),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1277),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1282),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1283),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1429),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1285),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1385),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1319),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1430),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1286),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1287),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1289),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1291),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1581),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1304),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1430),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1295),
.Y(n_1836)
);

CKINVDCx16_ASAP7_75t_R g1837 ( 
.A(n_1640),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1385),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1296),
.Y(n_1839)
);

INVxp67_ASAP7_75t_SL g1840 ( 
.A(n_1498),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1418),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1419),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1498),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1521),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1423),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1435),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1435),
.Y(n_1847)
);

NOR2xp67_ASAP7_75t_L g1848 ( 
.A(n_1437),
.B(n_866),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1426),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1427),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1304),
.Y(n_1851)
);

CKINVDCx16_ASAP7_75t_R g1852 ( 
.A(n_1253),
.Y(n_1852)
);

CKINVDCx20_ASAP7_75t_R g1853 ( 
.A(n_1614),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1437),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1447),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1521),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1438),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1447),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1273),
.B(n_794),
.Y(n_1859)
);

INVxp33_ASAP7_75t_SL g1860 ( 
.A(n_1464),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1464),
.Y(n_1861)
);

CKINVDCx20_ASAP7_75t_R g1862 ( 
.A(n_1624),
.Y(n_1862)
);

INVxp33_ASAP7_75t_SL g1863 ( 
.A(n_1467),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1308),
.Y(n_1864)
);

BUFx3_ASAP7_75t_L g1865 ( 
.A(n_1557),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1557),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_1635),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1467),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1496),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1496),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1439),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1245),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1440),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1511),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1441),
.Y(n_1875)
);

INVxp33_ASAP7_75t_SL g1876 ( 
.A(n_1511),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1442),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1513),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_SL g1879 ( 
.A(n_1483),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1443),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1513),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1308),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1444),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1516),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1516),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1445),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1446),
.Y(n_1887)
);

INVxp33_ASAP7_75t_SL g1888 ( 
.A(n_1517),
.Y(n_1888)
);

INVxp67_ASAP7_75t_SL g1889 ( 
.A(n_1448),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1517),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1450),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1257),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1522),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1522),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1451),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_1681),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1399),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1453),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1454),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1523),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1456),
.Y(n_1901)
);

CKINVDCx20_ASAP7_75t_R g1902 ( 
.A(n_1254),
.Y(n_1902)
);

INVxp33_ASAP7_75t_SL g1903 ( 
.A(n_1523),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1458),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1527),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1527),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1399),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1537),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1537),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1460),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1260),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1541),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_1310),
.Y(n_1913)
);

CKINVDCx16_ASAP7_75t_R g1914 ( 
.A(n_1359),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_1310),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1461),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1509),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1258),
.B(n_794),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1526),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1493),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1541),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1493),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1581),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1493),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1261),
.B(n_1030),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1324),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1324),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1551),
.Y(n_1928)
);

NOR2xp67_ASAP7_75t_L g1929 ( 
.A(n_1551),
.B(n_867),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1562),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1556),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1600),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1327),
.Y(n_1933)
);

CKINVDCx20_ASAP7_75t_R g1934 ( 
.A(n_1327),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1562),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1331),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1263),
.Y(n_1937)
);

INVxp33_ASAP7_75t_SL g1938 ( 
.A(n_1570),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1684),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1570),
.Y(n_1940)
);

NOR2xp67_ASAP7_75t_L g1941 ( 
.A(n_1585),
.B(n_868),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1315),
.B(n_794),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1585),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1264),
.Y(n_1944)
);

INVxp67_ASAP7_75t_SL g1945 ( 
.A(n_1265),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1595),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1595),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_1331),
.Y(n_1948)
);

CKINVDCx20_ASAP7_75t_R g1949 ( 
.A(n_1337),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1266),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1596),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1596),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1336),
.B(n_833),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1613),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1337),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_1343),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1270),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1271),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1274),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1684),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1613),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1298),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1343),
.Y(n_1963)
);

CKINVDCx20_ASAP7_75t_R g1964 ( 
.A(n_1350),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1350),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1360),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1565),
.B(n_1041),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1566),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1616),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1568),
.B(n_1041),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1360),
.Y(n_1971)
);

CKINVDCx20_ASAP7_75t_R g1972 ( 
.A(n_1368),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1392),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1569),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1417),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1342),
.B(n_833),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1571),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_1368),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1616),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1389),
.B(n_833),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1622),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1572),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_1377),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1576),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1622),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1578),
.Y(n_1986)
);

NOR2xp67_ASAP7_75t_L g1987 ( 
.A(n_1631),
.B(n_1633),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1580),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1401),
.B(n_833),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1582),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1377),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1583),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1631),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1420),
.B(n_833),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1413),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_1633),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1648),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1584),
.Y(n_1998)
);

CKINVDCx14_ASAP7_75t_R g1999 ( 
.A(n_1344),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_R g2000 ( 
.A(n_1648),
.B(n_872),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1466),
.B(n_1492),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1655),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1655),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1301),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1656),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1656),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1301),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1665),
.Y(n_2008)
);

INVxp67_ASAP7_75t_L g2009 ( 
.A(n_1518),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1586),
.Y(n_2010)
);

INVxp33_ASAP7_75t_L g2011 ( 
.A(n_1410),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1589),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_SL g2013 ( 
.A(n_1484),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1591),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1593),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1594),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1665),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1597),
.Y(n_2018)
);

INVxp67_ASAP7_75t_L g2019 ( 
.A(n_1567),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1668),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1601),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1602),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1668),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1670),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1603),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1606),
.B(n_1041),
.Y(n_2026)
);

CKINVDCx20_ASAP7_75t_R g2027 ( 
.A(n_1670),
.Y(n_2027)
);

NOR2xp67_ASAP7_75t_L g2028 ( 
.A(n_1679),
.B(n_873),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1608),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_1679),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_1685),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_1685),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1609),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1610),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1612),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1617),
.Y(n_2036)
);

CKINVDCx16_ASAP7_75t_R g2037 ( 
.A(n_1662),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1262),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1262),
.Y(n_2039)
);

INVxp33_ASAP7_75t_SL g2040 ( 
.A(n_1349),
.Y(n_2040)
);

CKINVDCx16_ASAP7_75t_R g2041 ( 
.A(n_1356),
.Y(n_2041)
);

CKINVDCx20_ASAP7_75t_R g2042 ( 
.A(n_1356),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1619),
.B(n_1041),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1621),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1623),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1625),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1339),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_1386),
.Y(n_2048)
);

INVxp67_ASAP7_75t_SL g2049 ( 
.A(n_1268),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1302),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1339),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2011),
.B(n_1672),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1741),
.Y(n_2053)
);

OA21x2_ASAP7_75t_L g2054 ( 
.A1(n_1925),
.A2(n_1244),
.B(n_1243),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1741),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_2049),
.B(n_1892),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_1697),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2040),
.A2(n_1472),
.B1(n_1579),
.B2(n_1676),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1699),
.B(n_1472),
.Y(n_2059)
);

INVx6_ASAP7_75t_L g2060 ( 
.A(n_1782),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1756),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1967),
.Y(n_2062)
);

BUFx6f_ASAP7_75t_L g2063 ( 
.A(n_1782),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1756),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1767),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1692),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1970),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1962),
.B(n_1695),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2026),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2043),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1692),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1719),
.Y(n_2072)
);

BUFx6f_ASAP7_75t_L g2073 ( 
.A(n_1827),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1693),
.Y(n_2074)
);

INVx3_ASAP7_75t_L g2075 ( 
.A(n_1827),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1892),
.B(n_1278),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1719),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1852),
.B(n_707),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_1865),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1738),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_1911),
.B(n_1400),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1693),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_2040),
.B(n_1312),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1706),
.B(n_1306),
.Y(n_2084)
);

AND2x2_ASAP7_75t_SL g2085 ( 
.A(n_1794),
.B(n_1400),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1767),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1738),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1778),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1778),
.Y(n_2089)
);

CKINVDCx20_ASAP7_75t_R g2090 ( 
.A(n_1700),
.Y(n_2090)
);

CKINVDCx20_ASAP7_75t_R g2091 ( 
.A(n_1701),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_1797),
.A2(n_1489),
.B1(n_1422),
.B2(n_1615),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1702),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1826),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_1865),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_1911),
.B(n_1489),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1826),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1838),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1838),
.Y(n_2099)
);

CKINVDCx20_ASAP7_75t_R g2100 ( 
.A(n_1710),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1897),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1689),
.B(n_1677),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_1866),
.Y(n_2103)
);

INVx2_ASAP7_75t_SL g2104 ( 
.A(n_1691),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1897),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1907),
.Y(n_2106)
);

AOI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1918),
.A2(n_1620),
.B1(n_710),
.B2(n_722),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1907),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_1999),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1866),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1975),
.Y(n_2111)
);

CKINVDCx20_ASAP7_75t_R g2112 ( 
.A(n_1716),
.Y(n_2112)
);

AND2x2_ASAP7_75t_SL g2113 ( 
.A(n_1709),
.B(n_1564),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1975),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2004),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1783),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_1698),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2004),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1944),
.B(n_1514),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2007),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2007),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2050),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2050),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_1944),
.B(n_1515),
.Y(n_2124)
);

CKINVDCx20_ASAP7_75t_R g2125 ( 
.A(n_1718),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1704),
.B(n_1677),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1937),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1730),
.B(n_1678),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1777),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_2001),
.A2(n_742),
.B1(n_758),
.B2(n_705),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1950),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1957),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_1783),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1958),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1746),
.B(n_1334),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1702),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1777),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1779),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1959),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1696),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1783),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1783),
.Y(n_2142)
);

INVx5_ASAP7_75t_L g2143 ( 
.A(n_1783),
.Y(n_2143)
);

CKINVDCx16_ASAP7_75t_R g2144 ( 
.A(n_1755),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1779),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1784),
.Y(n_2146)
);

OAI21x1_ASAP7_75t_L g2147 ( 
.A1(n_1784),
.A2(n_1244),
.B(n_1243),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1705),
.Y(n_2148)
);

INVxp67_ASAP7_75t_L g2149 ( 
.A(n_1711),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1707),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1785),
.Y(n_2151)
);

OA21x2_ASAP7_75t_L g2152 ( 
.A1(n_1688),
.A2(n_1249),
.B(n_1248),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1942),
.A2(n_765),
.B1(n_777),
.B2(n_762),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1708),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1785),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1712),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1859),
.B(n_1678),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1690),
.B(n_1680),
.Y(n_2158)
);

BUFx6f_ASAP7_75t_L g2159 ( 
.A(n_1787),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1787),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1920),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1703),
.Y(n_2162)
);

INVxp67_ASAP7_75t_L g2163 ( 
.A(n_1724),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1714),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1703),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_2042),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1920),
.Y(n_2167)
);

INVxp67_ASAP7_75t_L g2168 ( 
.A(n_1732),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1694),
.B(n_1680),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1945),
.B(n_1682),
.Y(n_2170)
);

AND2x6_ASAP7_75t_L g2171 ( 
.A(n_1917),
.B(n_1105),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1715),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_L g2173 ( 
.A(n_1953),
.B(n_1490),
.C(n_1487),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1922),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1922),
.Y(n_2175)
);

AND2x6_ASAP7_75t_L g2176 ( 
.A(n_1919),
.B(n_1121),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_1889),
.B(n_1491),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_1795),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1720),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1924),
.Y(n_2180)
);

BUFx6f_ASAP7_75t_L g2181 ( 
.A(n_1924),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_1814),
.Y(n_2182)
);

AND2x4_ASAP7_75t_L g2183 ( 
.A(n_1931),
.B(n_1494),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1721),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1817),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_1821),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_1822),
.Y(n_2187)
);

NOR2xp67_ASAP7_75t_L g2188 ( 
.A(n_1751),
.B(n_1497),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1823),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_1932),
.B(n_1500),
.Y(n_2190)
);

INVxp67_ASAP7_75t_L g2191 ( 
.A(n_1955),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1825),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1829),
.Y(n_2193)
);

BUFx3_ASAP7_75t_L g2194 ( 
.A(n_1830),
.Y(n_2194)
);

AND2x2_ASAP7_75t_SL g2195 ( 
.A(n_1764),
.B(n_1564),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1831),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1832),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2041),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1836),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1839),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1841),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1812),
.B(n_1682),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1842),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1845),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_2037),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1849),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1850),
.Y(n_2207)
);

INVxp33_ASAP7_75t_SL g2208 ( 
.A(n_1795),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1857),
.Y(n_2209)
);

OAI21x1_ASAP7_75t_L g2210 ( 
.A1(n_1725),
.A2(n_1249),
.B(n_1248),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1871),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1873),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1875),
.Y(n_2213)
);

INVx3_ASAP7_75t_L g2214 ( 
.A(n_1877),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1880),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1883),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1976),
.B(n_1683),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_1980),
.A2(n_793),
.B1(n_796),
.B2(n_780),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1886),
.Y(n_2219)
);

NOR2x1_ASAP7_75t_L g2220 ( 
.A(n_1987),
.B(n_1503),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1887),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1891),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1989),
.B(n_1994),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1895),
.Y(n_2224)
);

CKINVDCx20_ASAP7_75t_R g2225 ( 
.A(n_1728),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1898),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1899),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_1818),
.B(n_1713),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_1901),
.Y(n_2229)
);

INVx2_ASAP7_75t_SL g2230 ( 
.A(n_1742),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1904),
.Y(n_2231)
);

INVx4_ASAP7_75t_L g2232 ( 
.A(n_1968),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1910),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1753),
.B(n_1683),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1916),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1974),
.Y(n_2236)
);

INVxp67_ASAP7_75t_L g2237 ( 
.A(n_1955),
.Y(n_2237)
);

AND2x6_ASAP7_75t_L g2238 ( 
.A(n_1722),
.B(n_1121),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1977),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1729),
.Y(n_2240)
);

CKINVDCx20_ASAP7_75t_R g2241 ( 
.A(n_1737),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1982),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1984),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1986),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_1731),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_1733),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1988),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1734),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1990),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1992),
.Y(n_2250)
);

OR2x6_ASAP7_75t_L g2251 ( 
.A(n_2020),
.B(n_1686),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1736),
.Y(n_2252)
);

BUFx12f_ASAP7_75t_L g2253 ( 
.A(n_1796),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1743),
.Y(n_2254)
);

OAI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_1748),
.A2(n_844),
.B1(n_846),
.B2(n_842),
.Y(n_2255)
);

INVx3_ASAP7_75t_L g2256 ( 
.A(n_1744),
.Y(n_2256)
);

INVxp67_ASAP7_75t_L g2257 ( 
.A(n_2038),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_1745),
.B(n_1505),
.Y(n_2258)
);

AND2x6_ASAP7_75t_L g2259 ( 
.A(n_1747),
.B(n_1179),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1757),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_1998),
.B(n_1510),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_1796),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2010),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1759),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_1761),
.Y(n_2265)
);

BUFx3_ASAP7_75t_L g2266 ( 
.A(n_2012),
.Y(n_2266)
);

INVx3_ASAP7_75t_L g2267 ( 
.A(n_1762),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2014),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_1800),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2015),
.B(n_1370),
.Y(n_2270)
);

INVx6_ASAP7_75t_L g2271 ( 
.A(n_1781),
.Y(n_2271)
);

NOR2x1_ASAP7_75t_L g2272 ( 
.A(n_1848),
.B(n_1386),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_L g2273 ( 
.A(n_1788),
.B(n_1425),
.Y(n_2273)
);

OAI21x1_ASAP7_75t_L g2274 ( 
.A1(n_2016),
.A2(n_1252),
.B(n_1251),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1763),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_1788),
.B(n_2009),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2018),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2021),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2022),
.B(n_1686),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_2025),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_1995),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2029),
.B(n_1425),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2033),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1771),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2034),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_2035),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_2036),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1772),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1775),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_2019),
.B(n_1626),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1789),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2044),
.B(n_1627),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2045),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1790),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2046),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1791),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_1800),
.Y(n_2297)
);

INVx3_ASAP7_75t_L g2298 ( 
.A(n_1793),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_1973),
.Y(n_2299)
);

CKINVDCx20_ASAP7_75t_R g2300 ( 
.A(n_1749),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_SL g2301 ( 
.A1(n_2048),
.A2(n_1588),
.B1(n_829),
.B2(n_884),
.Y(n_2301)
);

CKINVDCx20_ASAP7_75t_R g2302 ( 
.A(n_1750),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1798),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_1799),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1801),
.Y(n_2305)
);

INVx3_ASAP7_75t_L g2306 ( 
.A(n_1802),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_1809),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1813),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1803),
.B(n_1628),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1717),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1726),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_1805),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_1751),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1840),
.Y(n_2314)
);

AND3x2_ASAP7_75t_L g2315 ( 
.A(n_1754),
.B(n_845),
.C(n_1179),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1843),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1844),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_1805),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1856),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_1806),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1879),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1879),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1879),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1929),
.B(n_853),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2013),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2013),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2013),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_1758),
.B(n_1629),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1941),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2028),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1723),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1723),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1833),
.B(n_1361),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1923),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_1752),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_1939),
.B(n_1671),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1960),
.B(n_1361),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2032),
.B(n_1673),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1860),
.B(n_1362),
.Y(n_2339)
);

CKINVDCx6p67_ASAP7_75t_R g2340 ( 
.A(n_1786),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1742),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_1752),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_1806),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1760),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1780),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_1810),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_1914),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_1808),
.B(n_1209),
.Y(n_2348)
);

INVx3_ASAP7_75t_L g2349 ( 
.A(n_1765),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1765),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1834),
.Y(n_2351)
);

AND3x2_ASAP7_75t_L g2352 ( 
.A(n_1851),
.B(n_1209),
.C(n_703),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_1768),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_1810),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_1864),
.B(n_702),
.Y(n_2355)
);

CKINVDCx8_ASAP7_75t_R g2356 ( 
.A(n_1815),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2000),
.B(n_1373),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_1768),
.Y(n_2358)
);

BUFx3_ASAP7_75t_L g2359 ( 
.A(n_1769),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_1769),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_1774),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1882),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_1774),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1860),
.B(n_1362),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_1824),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_2038),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_1824),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1776),
.Y(n_2368)
);

AND2x4_ASAP7_75t_L g2369 ( 
.A(n_1926),
.B(n_703),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_1828),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2039),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1936),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_2039),
.Y(n_2373)
);

INVx2_ASAP7_75t_SL g2374 ( 
.A(n_1792),
.Y(n_2374)
);

INVx3_ASAP7_75t_L g2375 ( 
.A(n_1776),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1863),
.B(n_1363),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1828),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_1835),
.B(n_1657),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_1863),
.B(n_1363),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1963),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_1835),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_1846),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_1846),
.B(n_1657),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1847),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_L g2385 ( 
.A(n_1847),
.Y(n_2385)
);

CKINVDCx5p33_ASAP7_75t_R g2386 ( 
.A(n_1854),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_1971),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1854),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_1855),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_1876),
.B(n_1364),
.Y(n_2390)
);

NAND2xp33_ASAP7_75t_L g2391 ( 
.A(n_1855),
.B(n_1041),
.Y(n_2391)
);

BUFx3_ASAP7_75t_L g2392 ( 
.A(n_1876),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_1858),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1858),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_1861),
.Y(n_2395)
);

NAND2xp33_ASAP7_75t_R g2396 ( 
.A(n_1861),
.B(n_1332),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_1868),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1868),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1869),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_1869),
.B(n_1660),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_1870),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_1870),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1874),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_1874),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_1878),
.Y(n_2405)
);

OAI22xp5_ASAP7_75t_SL g2406 ( 
.A1(n_2047),
.A2(n_890),
.B1(n_903),
.B2(n_874),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_1878),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_1888),
.B(n_1364),
.Y(n_2408)
);

AND2x4_ASAP7_75t_L g2409 ( 
.A(n_1881),
.B(n_714),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1888),
.B(n_1365),
.Y(n_2410)
);

AND2x6_ASAP7_75t_L g2411 ( 
.A(n_1872),
.B(n_714),
.Y(n_2411)
);

INVx6_ASAP7_75t_L g2412 ( 
.A(n_1837),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_1881),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1884),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1884),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1885),
.Y(n_2416)
);

NOR2x1_ASAP7_75t_L g2417 ( 
.A(n_1996),
.B(n_1661),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_1903),
.B(n_1365),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1903),
.B(n_1366),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1885),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1890),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_1890),
.B(n_1663),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1893),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1893),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_1894),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_1894),
.B(n_719),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_1938),
.B(n_1366),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_1900),
.Y(n_2428)
);

CKINVDCx16_ASAP7_75t_R g2429 ( 
.A(n_2006),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1938),
.B(n_1367),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_1900),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1905),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1905),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1906),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_1906),
.B(n_1908),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_SL g2436 ( 
.A(n_1804),
.B(n_798),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_1908),
.B(n_1367),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2047),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_1909),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_1909),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1912),
.Y(n_2441)
);

NAND2xp33_ASAP7_75t_L g2442 ( 
.A(n_1912),
.B(n_1041),
.Y(n_2442)
);

INVx4_ASAP7_75t_L g2443 ( 
.A(n_1921),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1921),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_1928),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2051),
.A2(n_852),
.B1(n_859),
.B2(n_850),
.Y(n_2446)
);

BUFx2_ASAP7_75t_L g2447 ( 
.A(n_1913),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_1928),
.B(n_1369),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_1930),
.B(n_1671),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1930),
.Y(n_2450)
);

AOI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2051),
.A2(n_877),
.B1(n_881),
.B2(n_880),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_1935),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_1935),
.B(n_1396),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_1940),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_1940),
.B(n_1369),
.Y(n_2455)
);

BUFx3_ASAP7_75t_L g2456 ( 
.A(n_1943),
.Y(n_2456)
);

BUFx2_ASAP7_75t_L g2457 ( 
.A(n_1915),
.Y(n_2457)
);

AND2x4_ASAP7_75t_L g2458 ( 
.A(n_1943),
.B(n_719),
.Y(n_2458)
);

HB1xp67_ASAP7_75t_L g2459 ( 
.A(n_1946),
.Y(n_2459)
);

XNOR2x2_ASAP7_75t_L g2460 ( 
.A(n_1766),
.B(n_955),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_1946),
.Y(n_2461)
);

CKINVDCx20_ASAP7_75t_R g2462 ( 
.A(n_1770),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_1947),
.Y(n_2463)
);

CKINVDCx20_ASAP7_75t_R g2464 ( 
.A(n_1773),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1947),
.B(n_1371),
.Y(n_2465)
);

BUFx2_ASAP7_75t_L g2466 ( 
.A(n_1927),
.Y(n_2466)
);

AND2x2_ASAP7_75t_SL g2467 ( 
.A(n_1766),
.B(n_1041),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_1951),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1951),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_1952),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_1952),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_1954),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_1954),
.B(n_720),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_1961),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_1961),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_1969),
.Y(n_2476)
);

OAI22xp5_ASAP7_75t_SL g2477 ( 
.A1(n_1807),
.A2(n_890),
.B1(n_903),
.B2(n_874),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2118),
.Y(n_2478)
);

INVx1_ASAP7_75t_SL g2479 ( 
.A(n_2057),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2115),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2115),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2121),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2118),
.Y(n_2483)
);

BUFx2_ASAP7_75t_L g2484 ( 
.A(n_2117),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2121),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2052),
.Y(n_2486)
);

INVx3_ASAP7_75t_L g2487 ( 
.A(n_2122),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2052),
.B(n_1969),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_2063),
.Y(n_2489)
);

INVxp67_ASAP7_75t_L g2490 ( 
.A(n_2057),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2120),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2122),
.Y(n_2492)
);

AOI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2085),
.A2(n_2083),
.B1(n_2058),
.B2(n_2092),
.Y(n_2493)
);

INVx1_ASAP7_75t_SL g2494 ( 
.A(n_2117),
.Y(n_2494)
);

CKINVDCx8_ASAP7_75t_R g2495 ( 
.A(n_2144),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2085),
.B(n_1979),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2090),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2120),
.Y(n_2498)
);

CKINVDCx8_ASAP7_75t_R g2499 ( 
.A(n_2144),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2053),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2068),
.B(n_1979),
.Y(n_2501)
);

INVxp67_ASAP7_75t_L g2502 ( 
.A(n_2104),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2063),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2223),
.B(n_2217),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2053),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2055),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2055),
.Y(n_2507)
);

XNOR2xp5_ASAP7_75t_L g2508 ( 
.A(n_2301),
.B(n_1811),
.Y(n_2508)
);

OAI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2085),
.A2(n_1985),
.B1(n_1993),
.B2(n_1981),
.Y(n_2509)
);

INVx3_ASAP7_75t_L g2510 ( 
.A(n_2063),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2123),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2123),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2063),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_2063),
.Y(n_2514)
);

NAND2xp33_ASAP7_75t_L g2515 ( 
.A(n_2146),
.B(n_1981),
.Y(n_2515)
);

OAI22xp5_ASAP7_75t_L g2516 ( 
.A1(n_2084),
.A2(n_1993),
.B1(n_1997),
.B2(n_1985),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2072),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2072),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2077),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2157),
.B(n_1997),
.Y(n_2520)
);

XOR2xp5_ASAP7_75t_L g2521 ( 
.A(n_2091),
.B(n_1816),
.Y(n_2521)
);

HB1xp67_ASAP7_75t_L g2522 ( 
.A(n_2198),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2061),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2061),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2077),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2379),
.B(n_2002),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2080),
.Y(n_2527)
);

BUFx8_ASAP7_75t_L g2528 ( 
.A(n_2166),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2128),
.B(n_2002),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2357),
.B(n_2003),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2080),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2087),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2087),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2064),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2098),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2381),
.B(n_2003),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2098),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2073),
.Y(n_2538)
);

INVxp67_ASAP7_75t_L g2539 ( 
.A(n_2104),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2073),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2064),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2105),
.Y(n_2542)
);

INVx3_ASAP7_75t_L g2543 ( 
.A(n_2073),
.Y(n_2543)
);

BUFx3_ASAP7_75t_L g2544 ( 
.A(n_2271),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_SL g2545 ( 
.A(n_2456),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2105),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2106),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2205),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2073),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2073),
.Y(n_2550)
);

AOI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2171),
.A2(n_2005),
.B1(n_2017),
.B2(n_2008),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_SL g2552 ( 
.A1(n_2406),
.A2(n_1820),
.B1(n_1853),
.B2(n_1819),
.Y(n_2552)
);

BUFx6f_ASAP7_75t_SL g2553 ( 
.A(n_2456),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2065),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_2079),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2065),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2106),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2171),
.A2(n_2008),
.B1(n_2017),
.B2(n_2005),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2381),
.B(n_2023),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2086),
.Y(n_2560)
);

AND3x1_ASAP7_75t_L g2561 ( 
.A(n_2273),
.B(n_724),
.C(n_720),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2111),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2357),
.B(n_2338),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2381),
.B(n_2023),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2086),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2088),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2338),
.B(n_2024),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2088),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2111),
.Y(n_2569)
);

INVx4_ASAP7_75t_L g2570 ( 
.A(n_2060),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2325),
.B(n_2326),
.Y(n_2571)
);

NOR2x1_ASAP7_75t_L g2572 ( 
.A(n_2188),
.B(n_2027),
.Y(n_2572)
);

BUFx6f_ASAP7_75t_SL g2573 ( 
.A(n_2392),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_2079),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2114),
.Y(n_2575)
);

BUFx6f_ASAP7_75t_L g2576 ( 
.A(n_2079),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2089),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2089),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2114),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2094),
.Y(n_2580)
);

BUFx6f_ASAP7_75t_L g2581 ( 
.A(n_2079),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2094),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2097),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2097),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2099),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2099),
.Y(n_2586)
);

BUFx6f_ASAP7_75t_L g2587 ( 
.A(n_2079),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2101),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2101),
.Y(n_2589)
);

AND2x4_ASAP7_75t_L g2590 ( 
.A(n_2325),
.B(n_2024),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_2381),
.B(n_1727),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2108),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2108),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2129),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2135),
.B(n_735),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2129),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2332),
.B(n_2030),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2137),
.Y(n_2598)
);

NAND3xp33_ASAP7_75t_L g2599 ( 
.A(n_2276),
.B(n_2031),
.C(n_1934),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2137),
.Y(n_2600)
);

INVxp67_ASAP7_75t_L g2601 ( 
.A(n_2347),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2138),
.Y(n_2602)
);

OAI22xp5_ASAP7_75t_SL g2603 ( 
.A1(n_2477),
.A2(n_1867),
.B1(n_1896),
.B2(n_1862),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_SL g2604 ( 
.A1(n_2100),
.A2(n_829),
.B1(n_884),
.B2(n_798),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2138),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2145),
.Y(n_2606)
);

OAI22xp5_ASAP7_75t_SL g2607 ( 
.A1(n_2112),
.A2(n_972),
.B1(n_1092),
.B2(n_896),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2145),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2151),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2271),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2151),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2155),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2059),
.B(n_1804),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2155),
.Y(n_2614)
);

NAND2xp33_ASAP7_75t_L g2615 ( 
.A(n_2146),
.B(n_1114),
.Y(n_2615)
);

NAND2xp33_ASAP7_75t_SL g2616 ( 
.A(n_2381),
.B(n_1966),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2160),
.Y(n_2617)
);

INVx4_ASAP7_75t_L g2618 ( 
.A(n_2060),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2332),
.B(n_1373),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2125),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2160),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2167),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2167),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2175),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2175),
.Y(n_2625)
);

BUFx8_ASAP7_75t_L g2626 ( 
.A(n_2166),
.Y(n_2626)
);

INVx3_ASAP7_75t_L g2627 ( 
.A(n_2075),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2180),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2385),
.B(n_1727),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2180),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2062),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2075),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2075),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2309),
.B(n_1043),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2290),
.B(n_1043),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2385),
.B(n_1735),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2328),
.B(n_1376),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2326),
.B(n_1933),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2146),
.Y(n_2639)
);

BUFx2_ASAP7_75t_L g2640 ( 
.A(n_2225),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2062),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2067),
.Y(n_2642)
);

OAI21x1_ASAP7_75t_L g2643 ( 
.A1(n_2147),
.A2(n_1272),
.B(n_1250),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2067),
.Y(n_2644)
);

BUFx6f_ASAP7_75t_L g2645 ( 
.A(n_2146),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2328),
.B(n_1376),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2210),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2069),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2210),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2069),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2174),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2331),
.B(n_1378),
.Y(n_2652)
);

BUFx2_ASAP7_75t_L g2653 ( 
.A(n_2241),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2331),
.B(n_1378),
.Y(n_2654)
);

HB1xp67_ASAP7_75t_L g2655 ( 
.A(n_2109),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_2174),
.Y(n_2656)
);

NAND2xp33_ASAP7_75t_SL g2657 ( 
.A(n_2385),
.B(n_1948),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2140),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2385),
.B(n_1735),
.Y(n_2659)
);

INVx1_ASAP7_75t_SL g2660 ( 
.A(n_2300),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2140),
.Y(n_2661)
);

NAND3xp33_ASAP7_75t_SL g2662 ( 
.A(n_2476),
.B(n_1956),
.C(n_1949),
.Y(n_2662)
);

INVx1_ASAP7_75t_SL g2663 ( 
.A(n_2302),
.Y(n_2663)
);

HB1xp67_ASAP7_75t_L g2664 ( 
.A(n_2281),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2148),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2148),
.Y(n_2666)
);

BUFx6f_ASAP7_75t_L g2667 ( 
.A(n_2146),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2150),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2150),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2154),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2174),
.Y(n_2671)
);

INVx1_ASAP7_75t_SL g2672 ( 
.A(n_2462),
.Y(n_2672)
);

NAND3xp33_ASAP7_75t_L g2673 ( 
.A(n_2153),
.B(n_1965),
.C(n_1964),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2054),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2171),
.B(n_735),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2054),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_SL g2677 ( 
.A(n_2356),
.B(n_1972),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2054),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2464),
.Y(n_2679)
);

BUFx6f_ASAP7_75t_L g2680 ( 
.A(n_2159),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2154),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2156),
.Y(n_2682)
);

INVx3_ASAP7_75t_L g2683 ( 
.A(n_2095),
.Y(n_2683)
);

BUFx6f_ASAP7_75t_L g2684 ( 
.A(n_2159),
.Y(n_2684)
);

INVxp67_ASAP7_75t_L g2685 ( 
.A(n_2299),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2070),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_2396),
.Y(n_2687)
);

INVxp67_ASAP7_75t_L g2688 ( 
.A(n_2436),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2054),
.Y(n_2689)
);

NAND2xp33_ASAP7_75t_R g2690 ( 
.A(n_2066),
.B(n_1739),
.Y(n_2690)
);

INVx3_ASAP7_75t_L g2691 ( 
.A(n_2095),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2095),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2081),
.B(n_1379),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2171),
.A2(n_1983),
.B1(n_1991),
.B2(n_1978),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2152),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2070),
.Y(n_2696)
);

NOR2x1_ASAP7_75t_L g2697 ( 
.A(n_2359),
.B(n_924),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_SL g2698 ( 
.A1(n_2208),
.A2(n_972),
.B1(n_1092),
.B2(n_896),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2187),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2187),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2103),
.Y(n_2701)
);

OAI22xp5_ASAP7_75t_SL g2702 ( 
.A1(n_2208),
.A2(n_1166),
.B1(n_976),
.B2(n_984),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2187),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2171),
.B(n_803),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2230),
.B(n_1739),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2152),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2199),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2152),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2199),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_L g2710 ( 
.A(n_2159),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2081),
.B(n_1379),
.Y(n_2711)
);

OAI22xp5_ASAP7_75t_SL g2712 ( 
.A1(n_2429),
.A2(n_1166),
.B1(n_976),
.B2(n_984),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2152),
.Y(n_2713)
);

BUFx2_ASAP7_75t_L g2714 ( 
.A(n_2251),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2199),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2385),
.B(n_853),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2214),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2214),
.Y(n_2718)
);

NAND2xp33_ASAP7_75t_SL g2719 ( 
.A(n_2393),
.B(n_924),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2274),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2274),
.Y(n_2721)
);

INVx3_ASAP7_75t_L g2722 ( 
.A(n_2103),
.Y(n_2722)
);

CKINVDCx20_ASAP7_75t_R g2723 ( 
.A(n_2429),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2159),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2214),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2159),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2076),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2224),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2161),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2224),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2224),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2127),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2161),
.Y(n_2733)
);

INVx1_ASAP7_75t_SL g2734 ( 
.A(n_2076),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2127),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2131),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2131),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2171),
.B(n_803),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2132),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2271),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2161),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2132),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2134),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2134),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2139),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2139),
.Y(n_2746)
);

BUFx3_ASAP7_75t_SL g2747 ( 
.A(n_2238),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2185),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2185),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2189),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2103),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2189),
.Y(n_2752)
);

AOI22xp5_ASAP7_75t_L g2753 ( 
.A1(n_2171),
.A2(n_1000),
.B1(n_1007),
.B2(n_996),
.Y(n_2753)
);

OAI22xp33_ASAP7_75t_L g2754 ( 
.A1(n_2107),
.A2(n_996),
.B1(n_1007),
.B2(n_1000),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2251),
.Y(n_2755)
);

AND2x4_ASAP7_75t_L g2756 ( 
.A(n_2081),
.B(n_724),
.Y(n_2756)
);

HB1xp67_ASAP7_75t_L g2757 ( 
.A(n_2251),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2161),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2204),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2204),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2176),
.B(n_755),
.Y(n_2761)
);

INVx3_ASAP7_75t_L g2762 ( 
.A(n_2110),
.Y(n_2762)
);

OAI22xp5_ASAP7_75t_SL g2763 ( 
.A1(n_2113),
.A2(n_1051),
.B1(n_1080),
.B2(n_1046),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2161),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_SL g2765 ( 
.A(n_2356),
.B(n_1046),
.Y(n_2765)
);

AOI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2176),
.A2(n_1080),
.B1(n_1081),
.B2(n_1051),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2181),
.Y(n_2767)
);

OAI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2232),
.A2(n_902),
.B1(n_904),
.B2(n_895),
.Y(n_2768)
);

INVxp67_ASAP7_75t_L g2769 ( 
.A(n_2366),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2176),
.B(n_1119),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2181),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2206),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2176),
.B(n_1119),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2181),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2181),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2206),
.Y(n_2776)
);

AOI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2176),
.A2(n_1101),
.B1(n_1141),
.B2(n_1081),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2181),
.Y(n_2778)
);

AND2x4_ASAP7_75t_L g2779 ( 
.A(n_2096),
.B(n_725),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2116),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2209),
.Y(n_2781)
);

HB1xp67_ASAP7_75t_L g2782 ( 
.A(n_2251),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2209),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2211),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2096),
.B(n_1380),
.Y(n_2785)
);

HB1xp67_ASAP7_75t_L g2786 ( 
.A(n_2149),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2250),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2250),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2250),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2232),
.A2(n_925),
.B1(n_938),
.B2(n_923),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2250),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2250),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2211),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2212),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2212),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2213),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2096),
.B(n_1380),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2263),
.Y(n_2798)
);

NAND2xp33_ASAP7_75t_SL g2799 ( 
.A(n_2393),
.B(n_1101),
.Y(n_2799)
);

INVx1_ASAP7_75t_SL g2800 ( 
.A(n_2271),
.Y(n_2800)
);

CKINVDCx5p33_ASAP7_75t_R g2801 ( 
.A(n_2178),
.Y(n_2801)
);

INVxp67_ASAP7_75t_L g2802 ( 
.A(n_2373),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2176),
.B(n_1106),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2176),
.B(n_1106),
.Y(n_2804)
);

INVx3_ASAP7_75t_L g2805 ( 
.A(n_2110),
.Y(n_2805)
);

BUFx6f_ASAP7_75t_L g2806 ( 
.A(n_2116),
.Y(n_2806)
);

INVx3_ASAP7_75t_L g2807 ( 
.A(n_2110),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2213),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2215),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2215),
.Y(n_2810)
);

CKINVDCx16_ASAP7_75t_R g2811 ( 
.A(n_2253),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2378),
.B(n_1381),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2219),
.Y(n_2813)
);

BUFx6f_ASAP7_75t_SL g2814 ( 
.A(n_2392),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2116),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2219),
.Y(n_2816)
);

INVx3_ASAP7_75t_L g2817 ( 
.A(n_2133),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2263),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2263),
.Y(n_2819)
);

INVx3_ASAP7_75t_SL g2820 ( 
.A(n_2340),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2263),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_SL g2822 ( 
.A(n_2393),
.B(n_853),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2393),
.B(n_853),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2263),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2280),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2133),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2156),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2164),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2163),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2164),
.Y(n_2830)
);

NAND2xp33_ASAP7_75t_SL g2831 ( 
.A(n_2393),
.B(n_1141),
.Y(n_2831)
);

NAND2x1_ASAP7_75t_L g2832 ( 
.A(n_2060),
.B(n_1333),
.Y(n_2832)
);

INVx3_ASAP7_75t_L g2833 ( 
.A(n_2133),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2172),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2172),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2378),
.B(n_1381),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2280),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2179),
.Y(n_2838)
);

OAI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2232),
.A2(n_944),
.B1(n_954),
.B2(n_943),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2179),
.Y(n_2840)
);

BUFx8_ASAP7_75t_L g2841 ( 
.A(n_2447),
.Y(n_2841)
);

OAI21x1_ASAP7_75t_L g2842 ( 
.A1(n_2147),
.A2(n_1272),
.B(n_1250),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2102),
.B(n_755),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2116),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_SL g2845 ( 
.A(n_2253),
.B(n_1147),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2240),
.Y(n_2846)
);

AND2x4_ASAP7_75t_L g2847 ( 
.A(n_2056),
.B(n_725),
.Y(n_2847)
);

BUFx6f_ASAP7_75t_SL g2848 ( 
.A(n_2359),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2240),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2280),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2060),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2221),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2221),
.Y(n_2853)
);

OAI21x1_ASAP7_75t_L g2854 ( 
.A1(n_2184),
.A2(n_1292),
.B(n_1290),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2222),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2222),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2226),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2056),
.B(n_726),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2226),
.Y(n_2859)
);

INVx1_ASAP7_75t_SL g2860 ( 
.A(n_2412),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2116),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2126),
.B(n_797),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2227),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_SL g2864 ( 
.A1(n_2113),
.A2(n_1149),
.B1(n_1191),
.B2(n_1147),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2227),
.Y(n_2865)
);

INVx1_ASAP7_75t_SL g2866 ( 
.A(n_2412),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2397),
.B(n_853),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2234),
.B(n_1059),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2397),
.B(n_883),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_2168),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2280),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2141),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_SL g2873 ( 
.A(n_2397),
.B(n_883),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2383),
.B(n_1382),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_2397),
.B(n_883),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2231),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2231),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2383),
.B(n_1059),
.Y(n_2878)
);

INVxp67_ASAP7_75t_L g2879 ( 
.A(n_2438),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2235),
.Y(n_2880)
);

BUFx6f_ASAP7_75t_L g2881 ( 
.A(n_2141),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2182),
.Y(n_2882)
);

AND2x6_ASAP7_75t_L g2883 ( 
.A(n_2321),
.B(n_970),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2280),
.Y(n_2884)
);

HB1xp67_ASAP7_75t_L g2885 ( 
.A(n_2230),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2235),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2400),
.B(n_797),
.Y(n_2887)
);

INVx3_ASAP7_75t_L g2888 ( 
.A(n_2182),
.Y(n_2888)
);

HB1xp67_ASAP7_75t_L g2889 ( 
.A(n_2447),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2236),
.Y(n_2890)
);

AND2x4_ASAP7_75t_L g2891 ( 
.A(n_2056),
.B(n_726),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2286),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2236),
.Y(n_2893)
);

BUFx6f_ASAP7_75t_L g2894 ( 
.A(n_2141),
.Y(n_2894)
);

OAI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2334),
.A2(n_1035),
.B1(n_1036),
.B2(n_974),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2239),
.Y(n_2896)
);

CKINVDCx8_ASAP7_75t_R g2897 ( 
.A(n_2178),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2239),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2242),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2400),
.B(n_934),
.Y(n_2900)
);

OAI22xp5_ASAP7_75t_SL g2901 ( 
.A1(n_2113),
.A2(n_1191),
.B1(n_1229),
.B2(n_1149),
.Y(n_2901)
);

OAI22xp5_ASAP7_75t_SL g2902 ( 
.A1(n_2195),
.A2(n_1235),
.B1(n_1229),
.B2(n_1902),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2412),
.Y(n_2903)
);

AOI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2228),
.A2(n_1235),
.B1(n_934),
.B2(n_818),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2242),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2243),
.Y(n_2906)
);

INVxp67_ASAP7_75t_L g2907 ( 
.A(n_2457),
.Y(n_2907)
);

AOI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2228),
.A2(n_818),
.B1(n_1082),
.B2(n_970),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2243),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2244),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2244),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2247),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2247),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2422),
.B(n_1382),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2182),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2249),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2249),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2422),
.B(n_1371),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2286),
.Y(n_2919)
);

INVx4_ASAP7_75t_SL g2920 ( 
.A(n_2639),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2504),
.B(n_2449),
.Y(n_2921)
);

AOI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2493),
.A2(n_2269),
.B1(n_2297),
.B2(n_2262),
.Y(n_2922)
);

INVxp67_ASAP7_75t_L g2923 ( 
.A(n_2484),
.Y(n_2923)
);

NOR3xp33_ASAP7_75t_L g2924 ( 
.A(n_2509),
.B(n_2371),
.C(n_2257),
.Y(n_2924)
);

AND2x4_ASAP7_75t_L g2925 ( 
.A(n_2544),
.B(n_2463),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2478),
.Y(n_2926)
);

BUFx3_ASAP7_75t_L g2927 ( 
.A(n_2544),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2478),
.Y(n_2928)
);

INVx1_ASAP7_75t_SL g2929 ( 
.A(n_2479),
.Y(n_2929)
);

AND2x2_ASAP7_75t_SL g2930 ( 
.A(n_2496),
.B(n_2467),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2610),
.Y(n_2931)
);

CKINVDCx20_ASAP7_75t_R g2932 ( 
.A(n_2521),
.Y(n_2932)
);

INVx2_ASAP7_75t_SL g2933 ( 
.A(n_2610),
.Y(n_2933)
);

INVx2_ASAP7_75t_SL g2934 ( 
.A(n_2639),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2563),
.B(n_2526),
.Y(n_2935)
);

AND2x6_ASAP7_75t_L g2936 ( 
.A(n_2747),
.B(n_2463),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2483),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2483),
.Y(n_2938)
);

INVxp67_ASAP7_75t_L g2939 ( 
.A(n_2484),
.Y(n_2939)
);

AND2x2_ASAP7_75t_SL g2940 ( 
.A(n_2496),
.B(n_2467),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2598),
.Y(n_2941)
);

AND2x4_ASAP7_75t_L g2942 ( 
.A(n_2740),
.B(n_2463),
.Y(n_2942)
);

NAND2xp33_ASAP7_75t_L g2943 ( 
.A(n_2639),
.B(n_2397),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2501),
.B(n_2520),
.Y(n_2944)
);

AND2x4_ASAP7_75t_L g2945 ( 
.A(n_2800),
.B(n_2463),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2491),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_SL g2947 ( 
.A(n_2801),
.B(n_2262),
.Y(n_2947)
);

INVx2_ASAP7_75t_SL g2948 ( 
.A(n_2639),
.Y(n_2948)
);

AND2x4_ASAP7_75t_L g2949 ( 
.A(n_2860),
.B(n_2463),
.Y(n_2949)
);

AND2x4_ASAP7_75t_L g2950 ( 
.A(n_2866),
.B(n_2401),
.Y(n_2950)
);

AND2x4_ASAP7_75t_L g2951 ( 
.A(n_2903),
.B(n_2401),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2491),
.Y(n_2952)
);

AND2x6_ASAP7_75t_L g2953 ( 
.A(n_2695),
.B(n_2401),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2567),
.B(n_2195),
.Y(n_2954)
);

BUFx3_ASAP7_75t_L g2955 ( 
.A(n_2820),
.Y(n_2955)
);

BUFx2_ASAP7_75t_L g2956 ( 
.A(n_2494),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2529),
.B(n_2449),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2567),
.B(n_2195),
.Y(n_2958)
);

BUFx10_ASAP7_75t_L g2959 ( 
.A(n_2545),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2812),
.B(n_2453),
.Y(n_2960)
);

NOR2xp33_ASAP7_75t_L g2961 ( 
.A(n_2530),
.B(n_2269),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2812),
.B(n_2453),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2490),
.B(n_2297),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2639),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2763),
.A2(n_2411),
.B1(n_2467),
.B2(n_2259),
.Y(n_2965)
);

OAI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2753),
.A2(n_2777),
.B1(n_2766),
.B2(n_2558),
.Y(n_2966)
);

INVxp67_ASAP7_75t_SL g2967 ( 
.A(n_2645),
.Y(n_2967)
);

AND2x4_ASAP7_75t_L g2968 ( 
.A(n_2714),
.B(n_2401),
.Y(n_2968)
);

INVx5_ASAP7_75t_L g2969 ( 
.A(n_2645),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2498),
.Y(n_2970)
);

AOI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2488),
.A2(n_2318),
.B1(n_2320),
.B2(n_2312),
.Y(n_2971)
);

NOR2xp33_ASAP7_75t_L g2972 ( 
.A(n_2613),
.B(n_2312),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2836),
.B(n_2349),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2498),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2598),
.Y(n_2975)
);

BUFx6f_ASAP7_75t_L g2976 ( 
.A(n_2645),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2608),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2608),
.Y(n_2978)
);

INVx1_ASAP7_75t_SL g2979 ( 
.A(n_2497),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2732),
.Y(n_2980)
);

NAND2x1p5_ASAP7_75t_L g2981 ( 
.A(n_2645),
.B(n_2401),
.Y(n_2981)
);

BUFx10_ASAP7_75t_L g2982 ( 
.A(n_2545),
.Y(n_2982)
);

INVx4_ASAP7_75t_L g2983 ( 
.A(n_2645),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2836),
.B(n_2874),
.Y(n_2984)
);

INVx2_ASAP7_75t_SL g2985 ( 
.A(n_2667),
.Y(n_2985)
);

AND2x4_ASAP7_75t_L g2986 ( 
.A(n_2714),
.B(n_2404),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2667),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2611),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2732),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2735),
.Y(n_2990)
);

NAND3x1_ASAP7_75t_L g2991 ( 
.A(n_2904),
.B(n_2363),
.C(n_2349),
.Y(n_2991)
);

BUFx2_ASAP7_75t_L g2992 ( 
.A(n_2640),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2551),
.B(n_2404),
.Y(n_2993)
);

BUFx3_ASAP7_75t_L g2994 ( 
.A(n_2820),
.Y(n_2994)
);

CKINVDCx6p67_ASAP7_75t_R g2995 ( 
.A(n_2573),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2611),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2594),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_SL g2998 ( 
.A(n_2801),
.B(n_2318),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2735),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2736),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2631),
.A2(n_2363),
.B1(n_2375),
.B2(n_2349),
.Y(n_3001)
);

OR2x2_ASAP7_75t_L g3002 ( 
.A(n_2521),
.B(n_2620),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2622),
.Y(n_3003)
);

INVx5_ASAP7_75t_L g3004 ( 
.A(n_2667),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2622),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2864),
.A2(n_2411),
.B1(n_2259),
.B2(n_2238),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2874),
.B(n_2914),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2590),
.B(n_2404),
.Y(n_3008)
);

BUFx3_ASAP7_75t_L g3009 ( 
.A(n_2495),
.Y(n_3009)
);

CKINVDCx5p33_ASAP7_75t_R g3010 ( 
.A(n_2690),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2736),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2737),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_SL g3013 ( 
.A1(n_2698),
.A2(n_2343),
.B1(n_2346),
.B2(n_2320),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2914),
.B(n_2363),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2495),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2693),
.B(n_2279),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_2897),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2693),
.B(n_2279),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2500),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2594),
.Y(n_3020)
);

HB1xp67_ASAP7_75t_L g3021 ( 
.A(n_2664),
.Y(n_3021)
);

BUFx3_ASAP7_75t_L g3022 ( 
.A(n_2499),
.Y(n_3022)
);

BUFx2_ASAP7_75t_L g3023 ( 
.A(n_2640),
.Y(n_3023)
);

HB1xp67_ASAP7_75t_L g3024 ( 
.A(n_2548),
.Y(n_3024)
);

AND2x4_ASAP7_75t_L g3025 ( 
.A(n_2590),
.B(n_2404),
.Y(n_3025)
);

AND2x4_ASAP7_75t_L g3026 ( 
.A(n_2590),
.B(n_2571),
.Y(n_3026)
);

AND2x6_ASAP7_75t_L g3027 ( 
.A(n_2695),
.B(n_2404),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2500),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2596),
.Y(n_3029)
);

INVx4_ASAP7_75t_SL g3030 ( 
.A(n_2667),
.Y(n_3030)
);

INVx6_ASAP7_75t_L g3031 ( 
.A(n_2570),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2596),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2635),
.B(n_2637),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2901),
.A2(n_2754),
.B1(n_2902),
.B2(n_2411),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2600),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2667),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2502),
.B(n_2343),
.Y(n_3037)
);

AND2x4_ASAP7_75t_L g3038 ( 
.A(n_2571),
.B(n_2405),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_2499),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2600),
.Y(n_3040)
);

AND2x6_ASAP7_75t_L g3041 ( 
.A(n_2706),
.B(n_2405),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2602),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2505),
.Y(n_3043)
);

AND2x4_ASAP7_75t_L g3044 ( 
.A(n_2571),
.B(n_2405),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2602),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2711),
.B(n_2279),
.Y(n_3046)
);

BUFx3_ASAP7_75t_L g3047 ( 
.A(n_2528),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2605),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2539),
.B(n_2346),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2528),
.Y(n_3050)
);

INVx1_ASAP7_75t_SL g3051 ( 
.A(n_2660),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2505),
.Y(n_3052)
);

CKINVDCx5p33_ASAP7_75t_R g3053 ( 
.A(n_2897),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2637),
.B(n_2646),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2488),
.B(n_2405),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2769),
.B(n_2405),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2737),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2739),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2802),
.B(n_2354),
.Y(n_3059)
);

AO22x2_ASAP7_75t_L g3060 ( 
.A1(n_2706),
.A2(n_2460),
.B1(n_2473),
.B2(n_2426),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2739),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2742),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2742),
.Y(n_3063)
);

INVxp67_ASAP7_75t_SL g3064 ( 
.A(n_2680),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2743),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_L g3066 ( 
.A(n_2879),
.B(n_2354),
.Y(n_3066)
);

INVx4_ASAP7_75t_L g3067 ( 
.A(n_2680),
.Y(n_3067)
);

NAND2x1p5_ASAP7_75t_L g3068 ( 
.A(n_2680),
.B(n_2431),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2506),
.Y(n_3069)
);

AND2x6_ASAP7_75t_L g3070 ( 
.A(n_2708),
.B(n_2431),
.Y(n_3070)
);

INVxp33_ASAP7_75t_SL g3071 ( 
.A(n_2677),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2506),
.Y(n_3072)
);

AND2x6_ASAP7_75t_L g3073 ( 
.A(n_2708),
.B(n_2431),
.Y(n_3073)
);

AND2x4_ASAP7_75t_L g3074 ( 
.A(n_2711),
.B(n_2431),
.Y(n_3074)
);

OAI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_2631),
.A2(n_2642),
.B1(n_2644),
.B2(n_2641),
.Y(n_3075)
);

OAI22xp5_ASAP7_75t_L g3076 ( 
.A1(n_2641),
.A2(n_2375),
.B1(n_2384),
.B2(n_2377),
.Y(n_3076)
);

BUFx2_ASAP7_75t_L g3077 ( 
.A(n_2653),
.Y(n_3077)
);

BUFx10_ASAP7_75t_L g3078 ( 
.A(n_2545),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2507),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2743),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2507),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2744),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2744),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2745),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2785),
.B(n_2341),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2680),
.Y(n_3086)
);

INVxp67_ASAP7_75t_SL g3087 ( 
.A(n_2680),
.Y(n_3087)
);

AND2x4_ASAP7_75t_L g3088 ( 
.A(n_2785),
.B(n_2431),
.Y(n_3088)
);

INVxp67_ASAP7_75t_SL g3089 ( 
.A(n_2684),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2523),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_SL g3091 ( 
.A(n_2685),
.B(n_2313),
.Y(n_3091)
);

INVx3_ASAP7_75t_L g3092 ( 
.A(n_2684),
.Y(n_3092)
);

INVx4_ASAP7_75t_L g3093 ( 
.A(n_2684),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2745),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_L g3095 ( 
.A(n_2516),
.B(n_2365),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2746),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2684),
.Y(n_3097)
);

BUFx10_ASAP7_75t_L g3098 ( 
.A(n_2553),
.Y(n_3098)
);

CKINVDCx5p33_ASAP7_75t_R g3099 ( 
.A(n_2811),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2746),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2705),
.B(n_2365),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2748),
.Y(n_3102)
);

AOI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_2515),
.A2(n_2370),
.B1(n_2382),
.B2(n_2367),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2523),
.Y(n_3104)
);

OAI221xp5_ASAP7_75t_L g3105 ( 
.A1(n_2561),
.A2(n_2451),
.B1(n_2218),
.B2(n_2191),
.C(n_2237),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2524),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2748),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_2885),
.B(n_2313),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2524),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2534),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_2705),
.B(n_2313),
.Y(n_3111)
);

BUFx6f_ASAP7_75t_L g3112 ( 
.A(n_2684),
.Y(n_3112)
);

BUFx3_ASAP7_75t_L g3113 ( 
.A(n_2528),
.Y(n_3113)
);

INVx4_ASAP7_75t_L g3114 ( 
.A(n_2710),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2534),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_2710),
.Y(n_3116)
);

NOR2xp33_ASAP7_75t_L g3117 ( 
.A(n_2601),
.B(n_2367),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2541),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_2710),
.Y(n_3119)
);

INVx2_ASAP7_75t_SL g3120 ( 
.A(n_2710),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2797),
.B(n_2341),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2541),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2554),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2605),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2646),
.B(n_2375),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_SL g3126 ( 
.A(n_2719),
.B(n_2313),
.Y(n_3126)
);

BUFx2_ASAP7_75t_L g3127 ( 
.A(n_2653),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2710),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2606),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_L g3130 ( 
.A(n_2734),
.B(n_2370),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2606),
.Y(n_3131)
);

INVx3_ASAP7_75t_L g3132 ( 
.A(n_2570),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2609),
.Y(n_3133)
);

INVx1_ASAP7_75t_SL g3134 ( 
.A(n_2663),
.Y(n_3134)
);

BUFx3_ASAP7_75t_L g3135 ( 
.A(n_2626),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2554),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2595),
.B(n_2339),
.Y(n_3137)
);

OR2x2_ASAP7_75t_L g3138 ( 
.A(n_2672),
.B(n_2457),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2786),
.B(n_2382),
.Y(n_3139)
);

BUFx2_ASAP7_75t_L g3140 ( 
.A(n_2889),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2749),
.Y(n_3141)
);

BUFx6f_ASAP7_75t_L g3142 ( 
.A(n_2780),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2749),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_SL g3144 ( 
.A(n_2799),
.B(n_2313),
.Y(n_3144)
);

BUFx2_ASAP7_75t_L g3145 ( 
.A(n_2522),
.Y(n_3145)
);

INVx4_ASAP7_75t_L g3146 ( 
.A(n_2570),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2750),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_2831),
.B(n_2335),
.Y(n_3148)
);

AND2x6_ASAP7_75t_L g3149 ( 
.A(n_2713),
.B(n_2335),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2750),
.Y(n_3150)
);

BUFx3_ASAP7_75t_L g3151 ( 
.A(n_2626),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2752),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2755),
.B(n_2335),
.Y(n_3153)
);

CKINVDCx5p33_ASAP7_75t_R g3154 ( 
.A(n_2573),
.Y(n_3154)
);

CKINVDCx5p33_ASAP7_75t_R g3155 ( 
.A(n_2573),
.Y(n_3155)
);

INVx4_ASAP7_75t_SL g3156 ( 
.A(n_2780),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2556),
.Y(n_3157)
);

OR2x2_ASAP7_75t_L g3158 ( 
.A(n_2597),
.B(n_2466),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2556),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_2757),
.B(n_2335),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2752),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2759),
.Y(n_3162)
);

BUFx6f_ASAP7_75t_L g3163 ( 
.A(n_2780),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2759),
.Y(n_3164)
);

INVx4_ASAP7_75t_L g3165 ( 
.A(n_2618),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2760),
.Y(n_3166)
);

INVx3_ASAP7_75t_L g3167 ( 
.A(n_2618),
.Y(n_3167)
);

NOR2xp33_ASAP7_75t_L g3168 ( 
.A(n_2829),
.B(n_2386),
.Y(n_3168)
);

NAND2x1p5_ASAP7_75t_L g3169 ( 
.A(n_2656),
.B(n_2184),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2760),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2843),
.B(n_2862),
.Y(n_3171)
);

AND2x4_ASAP7_75t_L g3172 ( 
.A(n_2797),
.B(n_2443),
.Y(n_3172)
);

BUFx6f_ASAP7_75t_L g3173 ( 
.A(n_2780),
.Y(n_3173)
);

AOI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_2515),
.A2(n_2407),
.B1(n_2413),
.B2(n_2386),
.Y(n_3174)
);

AND2x6_ASAP7_75t_L g3175 ( 
.A(n_2713),
.B(n_2335),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2560),
.Y(n_3176)
);

BUFx2_ASAP7_75t_L g3177 ( 
.A(n_2679),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2560),
.Y(n_3178)
);

NAND2xp33_ASAP7_75t_L g3179 ( 
.A(n_2651),
.B(n_2342),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_SL g3180 ( 
.A(n_2782),
.B(n_2342),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2772),
.Y(n_3181)
);

INVx5_ASAP7_75t_L g3182 ( 
.A(n_2780),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_2597),
.B(n_2342),
.Y(n_3183)
);

OAI22xp5_ASAP7_75t_L g3184 ( 
.A1(n_2642),
.A2(n_2384),
.B1(n_2389),
.B2(n_2377),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2565),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2772),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2776),
.Y(n_3187)
);

BUFx6f_ASAP7_75t_L g3188 ( 
.A(n_2806),
.Y(n_3188)
);

AOI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_2553),
.A2(n_2413),
.B1(n_2421),
.B2(n_2407),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2918),
.B(n_2364),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2776),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2781),
.Y(n_3192)
);

BUFx3_ASAP7_75t_L g3193 ( 
.A(n_2626),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2847),
.B(n_2270),
.Y(n_3194)
);

AOI22xp5_ASAP7_75t_L g3195 ( 
.A1(n_2553),
.A2(n_2445),
.B1(n_2452),
.B2(n_2421),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2870),
.B(n_2445),
.Y(n_3196)
);

NOR2xp67_ASAP7_75t_L g3197 ( 
.A(n_2687),
.B(n_2374),
.Y(n_3197)
);

OR2x2_ASAP7_75t_L g3198 ( 
.A(n_2878),
.B(n_2466),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2565),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2868),
.B(n_2376),
.Y(n_3200)
);

CKINVDCx5p33_ASAP7_75t_R g3201 ( 
.A(n_2814),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2609),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2634),
.B(n_2390),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2612),
.Y(n_3204)
);

CKINVDCx5p33_ASAP7_75t_R g3205 ( 
.A(n_2814),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2566),
.Y(n_3206)
);

INVx5_ASAP7_75t_L g3207 ( 
.A(n_2806),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2612),
.Y(n_3208)
);

INVx4_ASAP7_75t_SL g3209 ( 
.A(n_2806),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_2907),
.B(n_2452),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2566),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2614),
.Y(n_3212)
);

BUFx6f_ASAP7_75t_L g3213 ( 
.A(n_2806),
.Y(n_3213)
);

INVx1_ASAP7_75t_SL g3214 ( 
.A(n_2655),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2568),
.Y(n_3215)
);

HB1xp67_ASAP7_75t_L g3216 ( 
.A(n_2727),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_L g3217 ( 
.A1(n_2675),
.A2(n_2411),
.B1(n_2259),
.B2(n_2238),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2568),
.Y(n_3218)
);

BUFx10_ASAP7_75t_L g3219 ( 
.A(n_2848),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_2847),
.B(n_2443),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2781),
.B(n_2783),
.Y(n_3221)
);

AND2x4_ASAP7_75t_L g3222 ( 
.A(n_2847),
.B(n_2443),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2806),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_2858),
.B(n_2270),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_2486),
.B(n_2468),
.Y(n_3225)
);

AND2x4_ASAP7_75t_L g3226 ( 
.A(n_2858),
.B(n_2266),
.Y(n_3226)
);

INVx3_ASAP7_75t_L g3227 ( 
.A(n_2618),
.Y(n_3227)
);

AOI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_2848),
.A2(n_2474),
.B1(n_2476),
.B2(n_2468),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2577),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2614),
.Y(n_3230)
);

INVx1_ASAP7_75t_SL g3231 ( 
.A(n_2723),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2577),
.Y(n_3232)
);

INVx4_ASAP7_75t_SL g3233 ( 
.A(n_2815),
.Y(n_3233)
);

BUFx10_ASAP7_75t_L g3234 ( 
.A(n_2848),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2617),
.Y(n_3235)
);

INVx4_ASAP7_75t_L g3236 ( 
.A(n_2489),
.Y(n_3236)
);

CKINVDCx5p33_ASAP7_75t_R g3237 ( 
.A(n_2814),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_2858),
.B(n_2266),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2783),
.B(n_2408),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2617),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_2578),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2784),
.B(n_2410),
.Y(n_3242)
);

INVx2_ASAP7_75t_SL g3243 ( 
.A(n_2656),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_2578),
.Y(n_3244)
);

NAND3xp33_ASAP7_75t_L g3245 ( 
.A(n_2599),
.B(n_2474),
.C(n_2470),
.Y(n_3245)
);

AOI22xp33_ASAP7_75t_L g3246 ( 
.A1(n_2704),
.A2(n_2411),
.B1(n_2259),
.B2(n_2238),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_SL g3247 ( 
.A(n_2656),
.B(n_2342),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2621),
.Y(n_3248)
);

AND2x2_ASAP7_75t_SL g3249 ( 
.A(n_2765),
.B(n_2615),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2580),
.Y(n_3250)
);

BUFx6f_ASAP7_75t_L g3251 ( 
.A(n_2815),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_2580),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_2841),
.Y(n_3253)
);

CKINVDCx16_ASAP7_75t_R g3254 ( 
.A(n_2723),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2784),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_2583),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_2738),
.A2(n_2411),
.B1(n_2259),
.B2(n_2238),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_2688),
.B(n_2388),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2793),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_2891),
.B(n_2336),
.Y(n_3260)
);

INVx5_ASAP7_75t_L g3261 ( 
.A(n_2815),
.Y(n_3261)
);

AND2x2_ASAP7_75t_SL g3262 ( 
.A(n_2615),
.B(n_2342),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2583),
.Y(n_3263)
);

AND2x6_ASAP7_75t_L g3264 ( 
.A(n_2674),
.B(n_2358),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2793),
.B(n_2794),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2584),
.Y(n_3266)
);

BUFx2_ASAP7_75t_L g3267 ( 
.A(n_2841),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_2891),
.B(n_2336),
.Y(n_3268)
);

CKINVDCx5p33_ASAP7_75t_R g3269 ( 
.A(n_2687),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_2891),
.B(n_2177),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_2794),
.B(n_2177),
.Y(n_3271)
);

INVx2_ASAP7_75t_SL g3272 ( 
.A(n_2489),
.Y(n_3272)
);

NOR2xp33_ASAP7_75t_L g3273 ( 
.A(n_2694),
.B(n_2388),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2795),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_2616),
.B(n_2353),
.Y(n_3275)
);

BUFx2_ASAP7_75t_L g3276 ( 
.A(n_2841),
.Y(n_3276)
);

BUFx6f_ASAP7_75t_L g3277 ( 
.A(n_2815),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2584),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2795),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2796),
.B(n_2808),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_SL g3281 ( 
.A(n_2657),
.B(n_2353),
.Y(n_3281)
);

OR2x6_ASAP7_75t_L g3282 ( 
.A(n_2796),
.B(n_2412),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2585),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2808),
.Y(n_3284)
);

AND2x6_ASAP7_75t_L g3285 ( 
.A(n_2674),
.B(n_2353),
.Y(n_3285)
);

INVx5_ASAP7_75t_L g3286 ( 
.A(n_2815),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_2673),
.B(n_2394),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2585),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_2887),
.B(n_2394),
.Y(n_3289)
);

AOI22xp33_ASAP7_75t_L g3290 ( 
.A1(n_2761),
.A2(n_2411),
.B1(n_2259),
.B2(n_2238),
.Y(n_3290)
);

INVx1_ASAP7_75t_SL g3291 ( 
.A(n_2638),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2809),
.Y(n_3292)
);

INVxp67_ASAP7_75t_SL g3293 ( 
.A(n_2489),
.Y(n_3293)
);

BUFx10_ASAP7_75t_L g3294 ( 
.A(n_2638),
.Y(n_3294)
);

INVx4_ASAP7_75t_L g3295 ( 
.A(n_2489),
.Y(n_3295)
);

BUFx6f_ASAP7_75t_L g3296 ( 
.A(n_2844),
.Y(n_3296)
);

HB1xp67_ASAP7_75t_L g3297 ( 
.A(n_2638),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2809),
.Y(n_3298)
);

INVx4_ASAP7_75t_L g3299 ( 
.A(n_2489),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2810),
.Y(n_3300)
);

BUFx6f_ASAP7_75t_L g3301 ( 
.A(n_2844),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_2586),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_2586),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_2900),
.B(n_2353),
.Y(n_3304)
);

INVx2_ASAP7_75t_SL g3305 ( 
.A(n_2503),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2810),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2621),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_2813),
.B(n_2353),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2480),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2813),
.Y(n_3310)
);

AND2x4_ASAP7_75t_L g3311 ( 
.A(n_2658),
.B(n_2358),
.Y(n_3311)
);

AND2x2_ASAP7_75t_SL g3312 ( 
.A(n_2770),
.B(n_2361),
.Y(n_3312)
);

INVxp67_ASAP7_75t_L g3313 ( 
.A(n_2845),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_SL g3314 ( 
.A(n_2816),
.B(n_2358),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2816),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2852),
.Y(n_3316)
);

INVx4_ASAP7_75t_L g3317 ( 
.A(n_2503),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2852),
.Y(n_3318)
);

OR2x2_ASAP7_75t_L g3319 ( 
.A(n_2756),
.B(n_2340),
.Y(n_3319)
);

BUFx3_ASAP7_75t_L g3320 ( 
.A(n_2851),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2853),
.B(n_2418),
.Y(n_3321)
);

BUFx6f_ASAP7_75t_L g3322 ( 
.A(n_2844),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2853),
.B(n_2419),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_2503),
.Y(n_3324)
);

INVx4_ASAP7_75t_L g3325 ( 
.A(n_2503),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2855),
.B(n_2427),
.Y(n_3326)
);

AND2x4_ASAP7_75t_L g3327 ( 
.A(n_2661),
.B(n_2358),
.Y(n_3327)
);

NOR2xp33_ASAP7_75t_L g3328 ( 
.A(n_2536),
.B(n_2399),
.Y(n_3328)
);

INVx1_ASAP7_75t_SL g3329 ( 
.A(n_2508),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_2855),
.B(n_2358),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2856),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_2480),
.Y(n_3332)
);

BUFx3_ASAP7_75t_L g3333 ( 
.A(n_2851),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_SL g3334 ( 
.A(n_2856),
.B(n_2361),
.Y(n_3334)
);

OR2x2_ASAP7_75t_L g3335 ( 
.A(n_2756),
.B(n_2334),
.Y(n_3335)
);

INVx4_ASAP7_75t_L g3336 ( 
.A(n_2503),
.Y(n_3336)
);

INVx6_ASAP7_75t_L g3337 ( 
.A(n_2513),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_2559),
.B(n_2399),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_2857),
.B(n_2361),
.Y(n_3339)
);

BUFx6f_ASAP7_75t_L g3340 ( 
.A(n_2844),
.Y(n_3340)
);

OR2x6_ASAP7_75t_L g3341 ( 
.A(n_2857),
.B(n_2361),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_2481),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2481),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_2482),
.Y(n_3344)
);

INVx6_ASAP7_75t_L g3345 ( 
.A(n_2513),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2859),
.Y(n_3346)
);

BUFx2_ASAP7_75t_L g3347 ( 
.A(n_2756),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_2859),
.B(n_2863),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_L g3349 ( 
.A(n_2564),
.B(n_2403),
.Y(n_3349)
);

AND2x6_ASAP7_75t_L g3350 ( 
.A(n_2676),
.B(n_2361),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_2863),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2865),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_2865),
.B(n_2430),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2876),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_2482),
.Y(n_3355)
);

INVx3_ASAP7_75t_L g3356 ( 
.A(n_2513),
.Y(n_3356)
);

AND2x4_ASAP7_75t_L g3357 ( 
.A(n_2665),
.B(n_2666),
.Y(n_3357)
);

AOI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_2883),
.A2(n_2395),
.B1(n_2398),
.B2(n_2389),
.Y(n_3358)
);

OR2x2_ASAP7_75t_L g3359 ( 
.A(n_2779),
.B(n_2459),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_2876),
.B(n_2395),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2877),
.B(n_2398),
.Y(n_3361)
);

NAND2xp33_ASAP7_75t_L g3362 ( 
.A(n_2651),
.B(n_2402),
.Y(n_3362)
);

AOI22xp33_ASAP7_75t_L g3363 ( 
.A1(n_2773),
.A2(n_2259),
.B1(n_2238),
.B2(n_2426),
.Y(n_3363)
);

INVxp67_ASAP7_75t_SL g3364 ( 
.A(n_2513),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_2877),
.B(n_2402),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_2668),
.B(n_2321),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_2485),
.Y(n_3367)
);

OR2x2_ASAP7_75t_L g3368 ( 
.A(n_2779),
.B(n_2344),
.Y(n_3368)
);

INVx5_ASAP7_75t_L g3369 ( 
.A(n_2844),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_2880),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2485),
.Y(n_3371)
);

INVx3_ASAP7_75t_L g3372 ( 
.A(n_2513),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2492),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_2880),
.B(n_2425),
.Y(n_3374)
);

BUFx6f_ASAP7_75t_L g3375 ( 
.A(n_2861),
.Y(n_3375)
);

INVx5_ASAP7_75t_L g3376 ( 
.A(n_2861),
.Y(n_3376)
);

BUFx3_ASAP7_75t_L g3377 ( 
.A(n_2851),
.Y(n_3377)
);

AND2x6_ASAP7_75t_L g3378 ( 
.A(n_2676),
.B(n_2322),
.Y(n_3378)
);

CKINVDCx20_ASAP7_75t_R g3379 ( 
.A(n_2712),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_2886),
.B(n_2177),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2623),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_2492),
.Y(n_3382)
);

HB1xp67_ASAP7_75t_L g3383 ( 
.A(n_2779),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2623),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_2624),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_3026),
.B(n_2619),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2921),
.B(n_2425),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2941),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_2941),
.Y(n_3389)
);

AOI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_2972),
.A2(n_2702),
.B1(n_2414),
.B2(n_2415),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2935),
.B(n_2428),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3182),
.B(n_2882),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_2975),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_2975),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_2977),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3137),
.B(n_2428),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2962),
.B(n_2434),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3060),
.A2(n_2883),
.B1(n_2604),
.B2(n_2607),
.Y(n_3398)
);

AND2x6_ASAP7_75t_L g3399 ( 
.A(n_3220),
.B(n_3222),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2980),
.Y(n_3400)
);

CKINVDCx5p33_ASAP7_75t_R g3401 ( 
.A(n_3010),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2962),
.B(n_2434),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_2954),
.B(n_2409),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_2977),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_2978),
.Y(n_3405)
);

NAND3xp33_ASAP7_75t_L g3406 ( 
.A(n_3095),
.B(n_2414),
.C(n_2403),
.Y(n_3406)
);

O2A1O1Ixp5_ASAP7_75t_L g3407 ( 
.A1(n_2993),
.A2(n_2822),
.B(n_2823),
.C(n_2716),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_2978),
.Y(n_3408)
);

AOI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_3101),
.A2(n_2416),
.B1(n_2420),
.B2(n_2415),
.Y(n_3409)
);

NOR3xp33_ASAP7_75t_L g3410 ( 
.A(n_3013),
.B(n_2435),
.C(n_2662),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_L g3411 ( 
.A1(n_3060),
.A2(n_2883),
.B1(n_2804),
.B2(n_2803),
.Y(n_3411)
);

INVx2_ASAP7_75t_SL g3412 ( 
.A(n_2955),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3190),
.B(n_2439),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2989),
.Y(n_3414)
);

INVxp67_ASAP7_75t_L g3415 ( 
.A(n_2956),
.Y(n_3415)
);

NOR3xp33_ASAP7_75t_L g3416 ( 
.A(n_2961),
.B(n_3066),
.C(n_3059),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_2990),
.Y(n_3417)
);

OAI22xp5_ASAP7_75t_SL g3418 ( 
.A1(n_2932),
.A2(n_2552),
.B1(n_2603),
.B2(n_2508),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3200),
.B(n_2439),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3203),
.B(n_2440),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3033),
.B(n_2440),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2999),
.Y(n_3422)
);

INVx8_ASAP7_75t_L g3423 ( 
.A(n_3282),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3289),
.B(n_2441),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3271),
.B(n_2441),
.Y(n_3425)
);

NOR2xp33_ASAP7_75t_L g3426 ( 
.A(n_2944),
.B(n_2416),
.Y(n_3426)
);

NOR2xp33_ASAP7_75t_L g3427 ( 
.A(n_2957),
.B(n_2420),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3000),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3271),
.B(n_2444),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3380),
.B(n_2444),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3273),
.B(n_2423),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3060),
.A2(n_2883),
.B1(n_2650),
.B2(n_2644),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_SL g3433 ( 
.A(n_3182),
.B(n_2882),
.Y(n_3433)
);

AOI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3130),
.A2(n_2424),
.B1(n_2432),
.B2(n_2423),
.Y(n_3434)
);

AOI22x1_ASAP7_75t_L g3435 ( 
.A1(n_3169),
.A2(n_2671),
.B1(n_2886),
.B2(n_2475),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3380),
.B(n_2472),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_L g3437 ( 
.A(n_2954),
.B(n_2424),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2988),
.Y(n_3438)
);

INVx2_ASAP7_75t_SL g3439 ( 
.A(n_2955),
.Y(n_3439)
);

O2A1O1Ixp5_ASAP7_75t_L g3440 ( 
.A1(n_3304),
.A2(n_2869),
.B(n_2873),
.C(n_2867),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_SL g3441 ( 
.A(n_3182),
.B(n_3207),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_L g3442 ( 
.A(n_2958),
.B(n_2432),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_2984),
.B(n_2472),
.Y(n_3443)
);

INVx4_ASAP7_75t_L g3444 ( 
.A(n_2994),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_2984),
.B(n_2475),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_SL g3446 ( 
.A(n_3071),
.B(n_1740),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3007),
.B(n_2619),
.Y(n_3447)
);

NAND3xp33_ASAP7_75t_L g3448 ( 
.A(n_2963),
.B(n_2450),
.C(n_2433),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3182),
.B(n_2882),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3007),
.B(n_2433),
.Y(n_3450)
);

HB1xp67_ASAP7_75t_L g3451 ( 
.A(n_2956),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3060),
.A2(n_2966),
.B1(n_3034),
.B2(n_2930),
.Y(n_3452)
);

INVx2_ASAP7_75t_SL g3453 ( 
.A(n_2994),
.Y(n_3453)
);

BUFx6f_ASAP7_75t_SL g3454 ( 
.A(n_3047),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_2988),
.Y(n_3455)
);

AOI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_3179),
.A2(n_2721),
.B(n_2720),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_2960),
.B(n_2450),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3011),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_2958),
.B(n_2409),
.Y(n_3459)
);

INVx4_ASAP7_75t_L g3460 ( 
.A(n_3282),
.Y(n_3460)
);

CKINVDCx5p33_ASAP7_75t_R g3461 ( 
.A(n_3010),
.Y(n_3461)
);

O2A1O1Ixp33_ASAP7_75t_L g3462 ( 
.A1(n_3105),
.A2(n_2461),
.B(n_2469),
.C(n_2454),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3171),
.B(n_2454),
.Y(n_3463)
);

INVx2_ASAP7_75t_SL g3464 ( 
.A(n_2959),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_2996),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3054),
.B(n_2461),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_2996),
.Y(n_3467)
);

BUFx6f_ASAP7_75t_L g3468 ( 
.A(n_3182),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3194),
.B(n_2409),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_SL g3470 ( 
.A(n_3207),
.B(n_2888),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3194),
.B(n_2426),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3012),
.Y(n_3472)
);

NOR2x1p5_ASAP7_75t_L g3473 ( 
.A(n_3047),
.B(n_2066),
.Y(n_3473)
);

AOI22xp5_ASAP7_75t_L g3474 ( 
.A1(n_3117),
.A2(n_2470),
.B1(n_2471),
.B2(n_2469),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3003),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3003),
.Y(n_3476)
);

AOI22xp33_ASAP7_75t_L g3477 ( 
.A1(n_2930),
.A2(n_2940),
.B1(n_2965),
.B2(n_3006),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3016),
.B(n_2471),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_SL g3479 ( 
.A(n_3207),
.B(n_2888),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3005),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3005),
.Y(n_3481)
);

INVx3_ASAP7_75t_L g3482 ( 
.A(n_3146),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3057),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3309),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_3207),
.B(n_2888),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_2923),
.B(n_2350),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_SL g3487 ( 
.A(n_3207),
.B(n_2915),
.Y(n_3487)
);

AOI221xp5_ASAP7_75t_L g3488 ( 
.A1(n_3287),
.A2(n_2130),
.B1(n_2446),
.B2(n_2255),
.C(n_2895),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3016),
.B(n_2652),
.Y(n_3489)
);

NOR2xp33_ASAP7_75t_L g3490 ( 
.A(n_2939),
.B(n_2350),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3018),
.B(n_2652),
.Y(n_3491)
);

BUFx6f_ASAP7_75t_L g3492 ( 
.A(n_3261),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3309),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3058),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_L g3495 ( 
.A(n_2922),
.B(n_2360),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3224),
.B(n_2458),
.Y(n_3496)
);

BUFx6f_ASAP7_75t_L g3497 ( 
.A(n_3261),
.Y(n_3497)
);

NOR2xp67_ASAP7_75t_L g3498 ( 
.A(n_3017),
.B(n_2374),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3018),
.B(n_2654),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3046),
.B(n_2654),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_3261),
.B(n_2915),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_3359),
.B(n_2360),
.Y(n_3502)
);

BUFx3_ASAP7_75t_L g3503 ( 
.A(n_2927),
.Y(n_3503)
);

AO22x1_ASAP7_75t_L g3504 ( 
.A1(n_3071),
.A2(n_1740),
.B1(n_2074),
.B2(n_2071),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3046),
.B(n_2368),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3085),
.B(n_2368),
.Y(n_3506)
);

INVxp67_ASAP7_75t_SL g3507 ( 
.A(n_3142),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3239),
.A2(n_3321),
.B1(n_3323),
.B2(n_3242),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_3326),
.A2(n_2650),
.B1(n_2686),
.B2(n_2648),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_L g3510 ( 
.A1(n_2940),
.A2(n_2883),
.B1(n_2648),
.B2(n_2696),
.Y(n_3510)
);

NAND3xp33_ASAP7_75t_L g3511 ( 
.A(n_3258),
.B(n_2074),
.C(n_2071),
.Y(n_3511)
);

A2O1A1Ixp33_ASAP7_75t_L g3512 ( 
.A1(n_3125),
.A2(n_2696),
.B(n_2686),
.C(n_2511),
.Y(n_3512)
);

INVx8_ASAP7_75t_L g3513 ( 
.A(n_3282),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3085),
.B(n_2437),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3121),
.B(n_2448),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_3261),
.B(n_2915),
.Y(n_3516)
);

NOR2xp33_ASAP7_75t_SL g3517 ( 
.A(n_2947),
.B(n_2082),
.Y(n_3517)
);

BUFx5_ASAP7_75t_L g3518 ( 
.A(n_2953),
.Y(n_3518)
);

AOI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3210),
.A2(n_3139),
.B1(n_3196),
.B2(n_3168),
.Y(n_3519)
);

INVx2_ASAP7_75t_SL g3520 ( 
.A(n_2959),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3121),
.B(n_3353),
.Y(n_3521)
);

INVxp67_ASAP7_75t_L g3522 ( 
.A(n_3145),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3260),
.B(n_2455),
.Y(n_3523)
);

BUFx6f_ASAP7_75t_L g3524 ( 
.A(n_3261),
.Y(n_3524)
);

AOI22xp5_ASAP7_75t_L g3525 ( 
.A1(n_3225),
.A2(n_2082),
.B1(n_2136),
.B2(n_2093),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3061),
.Y(n_3526)
);

CKINVDCx20_ASAP7_75t_R g3527 ( 
.A(n_2932),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_SL g3528 ( 
.A(n_3286),
.B(n_2724),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3260),
.B(n_2465),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_3359),
.B(n_2344),
.Y(n_3530)
);

OAI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3221),
.A2(n_2671),
.B(n_2699),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3198),
.B(n_2345),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3268),
.B(n_2669),
.Y(n_3533)
);

AOI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_2998),
.A2(n_2093),
.B1(n_2162),
.B2(n_2136),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3268),
.B(n_2670),
.Y(n_3535)
);

INVx3_ASAP7_75t_L g3536 ( 
.A(n_3146),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3270),
.B(n_3224),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_3286),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3270),
.B(n_2681),
.Y(n_3539)
);

OAI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_3265),
.A2(n_2512),
.B1(n_2827),
.B2(n_2682),
.Y(n_3540)
);

AO22x1_ASAP7_75t_L g3541 ( 
.A1(n_3099),
.A2(n_2162),
.B1(n_2165),
.B2(n_2572),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3172),
.B(n_2828),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_SL g3543 ( 
.A(n_3099),
.B(n_2165),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3062),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3172),
.B(n_2830),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3172),
.B(n_2834),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3286),
.B(n_2724),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_SL g3548 ( 
.A(n_3286),
.B(n_2726),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_L g3549 ( 
.A1(n_3249),
.A2(n_2883),
.B1(n_2893),
.B2(n_2890),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3179),
.A2(n_2721),
.B(n_2720),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3357),
.B(n_2835),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3347),
.B(n_2458),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3357),
.B(n_2838),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_3286),
.B(n_2726),
.Y(n_3554)
);

HB1xp67_ASAP7_75t_L g3555 ( 
.A(n_3347),
.Y(n_3555)
);

NAND3xp33_ASAP7_75t_L g3556 ( 
.A(n_3037),
.B(n_2173),
.C(n_2272),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_L g3557 ( 
.A1(n_3249),
.A2(n_2883),
.B1(n_2936),
.B2(n_2893),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_3369),
.B(n_2729),
.Y(n_3558)
);

OAI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3280),
.A2(n_2700),
.B(n_2699),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_L g3560 ( 
.A(n_3198),
.B(n_2345),
.Y(n_3560)
);

OAI22xp33_ASAP7_75t_L g3561 ( 
.A1(n_3335),
.A2(n_2908),
.B1(n_2846),
.B2(n_2849),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_SL g3562 ( 
.A(n_3369),
.B(n_2729),
.Y(n_3562)
);

NOR2xp33_ASAP7_75t_L g3563 ( 
.A(n_3158),
.B(n_2351),
.Y(n_3563)
);

AOI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3049),
.A2(n_2078),
.B1(n_2362),
.B2(n_2351),
.Y(n_3564)
);

OR2x2_ASAP7_75t_L g3565 ( 
.A(n_3158),
.B(n_2362),
.Y(n_3565)
);

AND2x4_ASAP7_75t_SL g3566 ( 
.A(n_2959),
.B(n_2228),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_2943),
.A2(n_3362),
.B(n_3075),
.Y(n_3567)
);

A2O1A1Ixp33_ASAP7_75t_L g3568 ( 
.A1(n_2973),
.A2(n_2840),
.B(n_2896),
.C(n_2890),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3357),
.B(n_2202),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3348),
.B(n_2458),
.Y(n_3570)
);

HB1xp67_ASAP7_75t_L g3571 ( 
.A(n_3145),
.Y(n_3571)
);

NOR3xp33_ASAP7_75t_L g3572 ( 
.A(n_3245),
.B(n_2629),
.C(n_2591),
.Y(n_3572)
);

INVxp67_ASAP7_75t_L g3573 ( 
.A(n_2929),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_SL g3574 ( 
.A(n_3017),
.B(n_2315),
.Y(n_3574)
);

HB1xp67_ASAP7_75t_L g3575 ( 
.A(n_3383),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3063),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3065),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_SL g3578 ( 
.A(n_3053),
.B(n_3050),
.Y(n_3578)
);

INVx2_ASAP7_75t_SL g3579 ( 
.A(n_2982),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3332),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3348),
.B(n_2473),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3080),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3082),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_2971),
.B(n_2372),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3083),
.Y(n_3585)
);

NAND2xp33_ASAP7_75t_L g3586 ( 
.A(n_2953),
.B(n_2700),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3014),
.B(n_2473),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3332),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3084),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_SL g3590 ( 
.A(n_3369),
.B(n_2733),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3220),
.B(n_3222),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3220),
.B(n_3222),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3094),
.Y(n_3593)
);

INVxp67_ASAP7_75t_SL g3594 ( 
.A(n_3142),
.Y(n_3594)
);

OAI22x1_ASAP7_75t_SL g3595 ( 
.A1(n_3379),
.A2(n_1055),
.B1(n_1066),
.B2(n_1039),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3074),
.B(n_2170),
.Y(n_3596)
);

NOR2xp33_ASAP7_75t_L g3597 ( 
.A(n_3074),
.B(n_2372),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3074),
.B(n_2119),
.Y(n_3598)
);

INVx2_ASAP7_75t_SL g3599 ( 
.A(n_2982),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3088),
.B(n_2119),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3342),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_3369),
.B(n_2733),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3096),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_3088),
.B(n_2380),
.Y(n_3604)
);

AOI22xp5_ASAP7_75t_L g3605 ( 
.A1(n_3103),
.A2(n_3174),
.B1(n_3088),
.B2(n_3189),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3100),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3335),
.B(n_2380),
.Y(n_3607)
);

INVxp67_ASAP7_75t_L g3608 ( 
.A(n_3024),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3102),
.Y(n_3609)
);

NOR2xp33_ASAP7_75t_R g3610 ( 
.A(n_3053),
.B(n_2322),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3107),
.Y(n_3611)
);

BUFx6f_ASAP7_75t_SL g3612 ( 
.A(n_3050),
.Y(n_3612)
);

INVxp67_ASAP7_75t_L g3613 ( 
.A(n_3021),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_2943),
.A2(n_2649),
.B(n_2647),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3140),
.B(n_2387),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3141),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_3369),
.B(n_2741),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3226),
.B(n_2119),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3143),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3226),
.B(n_2124),
.Y(n_3620)
);

BUFx12f_ASAP7_75t_L g3621 ( 
.A(n_3154),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3147),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3150),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3226),
.B(n_3238),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3376),
.B(n_2741),
.Y(n_3625)
);

INVx2_ASAP7_75t_SL g3626 ( 
.A(n_2982),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3342),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3152),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3238),
.B(n_2124),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3161),
.Y(n_3630)
);

HB1xp67_ASAP7_75t_L g3631 ( 
.A(n_3140),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3162),
.Y(n_3632)
);

NOR2xp67_ASAP7_75t_L g3633 ( 
.A(n_3269),
.B(n_2323),
.Y(n_3633)
);

NOR2xp33_ASAP7_75t_SL g3634 ( 
.A(n_3113),
.B(n_2387),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3164),
.Y(n_3635)
);

AND2x6_ASAP7_75t_SL g3636 ( 
.A(n_3328),
.B(n_2355),
.Y(n_3636)
);

AOI22xp5_ASAP7_75t_L g3637 ( 
.A1(n_3195),
.A2(n_2697),
.B1(n_2417),
.B2(n_2659),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3238),
.B(n_2124),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3368),
.B(n_2282),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_3343),
.Y(n_3640)
);

OR2x2_ASAP7_75t_L g3641 ( 
.A(n_3002),
.B(n_2333),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_SL g3642 ( 
.A(n_3376),
.B(n_2969),
.Y(n_3642)
);

NOR2xp67_ASAP7_75t_L g3643 ( 
.A(n_3269),
.B(n_2323),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3008),
.B(n_2258),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3166),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3368),
.B(n_3319),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3376),
.B(n_2758),
.Y(n_3647)
);

NOR2x1p5_ASAP7_75t_L g3648 ( 
.A(n_3113),
.B(n_2327),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3008),
.B(n_3025),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3170),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3008),
.B(n_2258),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3025),
.B(n_2258),
.Y(n_3652)
);

NOR2xp33_ASAP7_75t_L g3653 ( 
.A(n_3319),
.B(n_2636),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3025),
.B(n_2348),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3343),
.Y(n_3655)
);

INVxp33_ASAP7_75t_SL g3656 ( 
.A(n_3228),
.Y(n_3656)
);

NOR2xp33_ASAP7_75t_R g3657 ( 
.A(n_3154),
.B(n_2327),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_R g3658 ( 
.A(n_3155),
.B(n_2510),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_SL g3659 ( 
.A(n_3376),
.B(n_2758),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3026),
.B(n_2348),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3026),
.B(n_2348),
.Y(n_3661)
);

BUFx3_ASAP7_75t_L g3662 ( 
.A(n_2927),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3361),
.B(n_2292),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3374),
.B(n_2292),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_3376),
.B(n_2764),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_2969),
.B(n_2764),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3344),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_2928),
.B(n_2337),
.Y(n_3668)
);

NOR3xp33_ASAP7_75t_L g3669 ( 
.A(n_2924),
.B(n_3055),
.C(n_3184),
.Y(n_3669)
);

INVx3_ASAP7_75t_L g3670 ( 
.A(n_3146),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3344),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3181),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3186),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3355),
.Y(n_3674)
);

INVx4_ASAP7_75t_L g3675 ( 
.A(n_3282),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_2928),
.B(n_2282),
.Y(n_3676)
);

AOI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_3214),
.A2(n_2355),
.B1(n_2369),
.B2(n_2220),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_2970),
.B(n_2183),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_2970),
.B(n_2183),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3187),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3355),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3191),
.B(n_2183),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3192),
.B(n_2190),
.Y(n_3683)
);

INVx2_ASAP7_75t_SL g3684 ( 
.A(n_3078),
.Y(n_3684)
);

CKINVDCx11_ASAP7_75t_R g3685 ( 
.A(n_3254),
.Y(n_3685)
);

NOR2xp33_ASAP7_75t_L g3686 ( 
.A(n_3216),
.B(n_2329),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3367),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3255),
.B(n_2190),
.Y(n_3688)
);

INVx3_ASAP7_75t_L g3689 ( 
.A(n_3165),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3297),
.B(n_2329),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3367),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_3362),
.A2(n_2649),
.B(n_2647),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_SL g3693 ( 
.A(n_2969),
.B(n_2767),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3259),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3274),
.B(n_2190),
.Y(n_3695)
);

NAND2xp33_ASAP7_75t_L g3696 ( 
.A(n_2953),
.B(n_2703),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3279),
.B(n_2355),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3371),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3284),
.B(n_2369),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_L g3700 ( 
.A(n_3338),
.B(n_2330),
.Y(n_3700)
);

INVxp67_ASAP7_75t_L g3701 ( 
.A(n_3138),
.Y(n_3701)
);

INVx3_ASAP7_75t_L g3702 ( 
.A(n_3165),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3292),
.B(n_2369),
.Y(n_3703)
);

OR2x2_ASAP7_75t_L g3704 ( 
.A(n_3002),
.B(n_2261),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3371),
.Y(n_3705)
);

BUFx2_ASAP7_75t_L g3706 ( 
.A(n_2992),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3298),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_L g3708 ( 
.A(n_3349),
.B(n_2330),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3300),
.B(n_2261),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3306),
.B(n_2261),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3310),
.Y(n_3711)
);

INVx2_ASAP7_75t_SL g3712 ( 
.A(n_3078),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3315),
.Y(n_3713)
);

AND2x4_ASAP7_75t_L g3714 ( 
.A(n_2968),
.B(n_2194),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3316),
.B(n_2896),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3318),
.B(n_2898),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3331),
.B(n_2898),
.Y(n_3717)
);

AND2x4_ASAP7_75t_L g3718 ( 
.A(n_2968),
.B(n_2194),
.Y(n_3718)
);

HB1xp67_ASAP7_75t_L g3719 ( 
.A(n_2992),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_SL g3720 ( 
.A(n_2969),
.B(n_2767),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3346),
.B(n_2899),
.Y(n_3721)
);

AOI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_2968),
.A2(n_2768),
.B1(n_2839),
.B2(n_2790),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3351),
.B(n_3352),
.Y(n_3723)
);

NAND2xp33_ASAP7_75t_L g3724 ( 
.A(n_2953),
.B(n_2703),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3354),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_SL g3726 ( 
.A(n_3135),
.B(n_2787),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3183),
.B(n_2184),
.Y(n_3727)
);

INVx1_ASAP7_75t_SL g3728 ( 
.A(n_2979),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3370),
.B(n_2899),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_L g3730 ( 
.A(n_3291),
.B(n_2245),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3373),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_2986),
.B(n_2905),
.Y(n_3732)
);

INVx3_ASAP7_75t_L g3733 ( 
.A(n_3165),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3111),
.B(n_2245),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_L g3735 ( 
.A(n_2986),
.B(n_2245),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_2986),
.B(n_2905),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_SL g3737 ( 
.A(n_2969),
.B(n_2771),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_2942),
.B(n_2906),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3373),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_SL g3740 ( 
.A(n_3004),
.B(n_2771),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_SL g3741 ( 
.A(n_3004),
.B(n_2774),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_2942),
.B(n_2906),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_2942),
.B(n_2909),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_2926),
.Y(n_3744)
);

O2A1O1Ixp33_ASAP7_75t_L g3745 ( 
.A1(n_3076),
.A2(n_2875),
.B(n_2324),
.C(n_2308),
.Y(n_3745)
);

BUFx6f_ASAP7_75t_L g3746 ( 
.A(n_3142),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_2937),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_2945),
.B(n_2909),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_2945),
.B(n_2910),
.Y(n_3749)
);

A2O1A1Ixp33_ASAP7_75t_L g3750 ( 
.A1(n_3358),
.A2(n_2911),
.B(n_2912),
.C(n_2910),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_2945),
.B(n_2911),
.Y(n_3751)
);

A2O1A1Ixp33_ASAP7_75t_L g3752 ( 
.A1(n_2938),
.A2(n_2952),
.B(n_2974),
.C(n_2946),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_2949),
.B(n_2912),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_2997),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_2997),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_2949),
.B(n_2913),
.Y(n_3756)
);

A2O1A1Ixp33_ASAP7_75t_L g3757 ( 
.A1(n_3020),
.A2(n_2916),
.B(n_2917),
.C(n_2913),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_2949),
.B(n_2916),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3020),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3029),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_SL g3761 ( 
.A(n_3135),
.B(n_2787),
.Y(n_3761)
);

BUFx2_ASAP7_75t_L g3762 ( 
.A(n_3023),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_2950),
.B(n_2917),
.Y(n_3763)
);

OR2x6_ASAP7_75t_L g3764 ( 
.A(n_3151),
.B(n_2788),
.Y(n_3764)
);

NAND2xp33_ASAP7_75t_L g3765 ( 
.A(n_2953),
.B(n_2707),
.Y(n_3765)
);

HB1xp67_ASAP7_75t_L g3766 ( 
.A(n_3023),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3029),
.Y(n_3767)
);

INVx2_ASAP7_75t_SL g3768 ( 
.A(n_3078),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3032),
.Y(n_3769)
);

AOI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_2991),
.A2(n_2709),
.B1(n_2715),
.B2(n_2707),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3382),
.Y(n_3771)
);

BUFx6f_ASAP7_75t_L g3772 ( 
.A(n_3142),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_SL g3773 ( 
.A(n_3004),
.B(n_2774),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_2950),
.B(n_2951),
.Y(n_3774)
);

AOI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_2991),
.A2(n_2715),
.B1(n_2717),
.B2(n_2709),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3382),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_L g3777 ( 
.A(n_3077),
.B(n_2246),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_2950),
.B(n_2246),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_2951),
.B(n_2246),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_2951),
.B(n_2248),
.Y(n_3780)
);

NOR2xp33_ASAP7_75t_L g3781 ( 
.A(n_3077),
.B(n_2248),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3038),
.B(n_2248),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_SL g3783 ( 
.A(n_3004),
.B(n_2775),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3388),
.Y(n_3784)
);

BUFx6f_ASAP7_75t_L g3785 ( 
.A(n_3468),
.Y(n_3785)
);

BUFx6f_ASAP7_75t_L g3786 ( 
.A(n_3468),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3389),
.Y(n_3787)
);

AND2x6_ASAP7_75t_SL g3788 ( 
.A(n_3431),
.B(n_2460),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3400),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3393),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3394),
.Y(n_3791)
);

BUFx8_ASAP7_75t_L g3792 ( 
.A(n_3454),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3431),
.B(n_3313),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3639),
.B(n_3127),
.Y(n_3794)
);

AOI22xp33_ASAP7_75t_L g3795 ( 
.A1(n_3398),
.A2(n_3379),
.B1(n_2936),
.B2(n_3144),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3426),
.B(n_3051),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_SL g3797 ( 
.A(n_3495),
.B(n_3262),
.Y(n_3797)
);

OR2x6_ASAP7_75t_L g3798 ( 
.A(n_3423),
.B(n_3151),
.Y(n_3798)
);

BUFx2_ASAP7_75t_L g3799 ( 
.A(n_3527),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3414),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3426),
.B(n_3134),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3417),
.Y(n_3802)
);

NOR2x1p5_ASAP7_75t_L g3803 ( 
.A(n_3621),
.B(n_3193),
.Y(n_3803)
);

CKINVDCx16_ASAP7_75t_R g3804 ( 
.A(n_3446),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3422),
.Y(n_3805)
);

OAI22xp5_ASAP7_75t_L g3806 ( 
.A1(n_3519),
.A2(n_3341),
.B1(n_3001),
.B2(n_3327),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3563),
.B(n_3038),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3398),
.A2(n_2936),
.B1(n_3148),
.B2(n_3126),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3395),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3428),
.Y(n_3810)
);

INVx3_ASAP7_75t_L g3811 ( 
.A(n_3399),
.Y(n_3811)
);

NOR2x1_ASAP7_75t_R g3812 ( 
.A(n_3685),
.B(n_3193),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3563),
.B(n_3038),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3458),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3530),
.B(n_3044),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3530),
.B(n_3044),
.Y(n_3816)
);

INVx2_ASAP7_75t_SL g3817 ( 
.A(n_3473),
.Y(n_3817)
);

BUFx2_ASAP7_75t_L g3818 ( 
.A(n_3706),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3404),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3532),
.B(n_3044),
.Y(n_3820)
);

INVxp67_ASAP7_75t_L g3821 ( 
.A(n_3451),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3405),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3532),
.B(n_3127),
.Y(n_3823)
);

NOR3xp33_ASAP7_75t_SL g3824 ( 
.A(n_3511),
.B(n_815),
.C(n_754),
.Y(n_3824)
);

AOI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3584),
.A2(n_3177),
.B1(n_3138),
.B2(n_3231),
.Y(n_3825)
);

A2O1A1Ixp33_ASAP7_75t_L g3826 ( 
.A1(n_3495),
.A2(n_3327),
.B(n_3311),
.C(n_3363),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3565),
.B(n_3177),
.Y(n_3827)
);

CKINVDCx5p33_ASAP7_75t_R g3828 ( 
.A(n_3401),
.Y(n_3828)
);

INVx3_ASAP7_75t_L g3829 ( 
.A(n_3399),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_SL g3830 ( 
.A(n_3700),
.B(n_3262),
.Y(n_3830)
);

INVx4_ASAP7_75t_L g3831 ( 
.A(n_3399),
.Y(n_3831)
);

BUFx2_ASAP7_75t_L g3832 ( 
.A(n_3762),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3472),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3483),
.Y(n_3834)
);

OR2x4_ASAP7_75t_L g3835 ( 
.A(n_3584),
.B(n_2304),
.Y(n_3835)
);

INVx4_ASAP7_75t_L g3836 ( 
.A(n_3399),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3560),
.B(n_3366),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3560),
.B(n_3366),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3494),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3526),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3408),
.Y(n_3841)
);

OR2x6_ASAP7_75t_L g3842 ( 
.A(n_3423),
.B(n_3253),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3607),
.B(n_3366),
.Y(n_3843)
);

NOR2xp33_ASAP7_75t_R g3844 ( 
.A(n_3461),
.B(n_3155),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3607),
.B(n_3521),
.Y(n_3845)
);

AOI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_3437),
.A2(n_3442),
.B1(n_3416),
.B2(n_3488),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3427),
.B(n_3009),
.Y(n_3847)
);

AND2x6_ASAP7_75t_L g3848 ( 
.A(n_3468),
.B(n_3032),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3427),
.B(n_3437),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3442),
.B(n_3009),
.Y(n_3850)
);

NAND2x1p5_ASAP7_75t_L g3851 ( 
.A(n_3460),
.B(n_3004),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3463),
.B(n_3015),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3438),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3502),
.B(n_3015),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3455),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3544),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3465),
.Y(n_3857)
);

NAND2x1p5_ASAP7_75t_L g3858 ( 
.A(n_3460),
.B(n_2925),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3467),
.Y(n_3859)
);

O2A1O1Ixp33_ASAP7_75t_L g3860 ( 
.A1(n_3424),
.A2(n_3365),
.B(n_3360),
.C(n_3091),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3475),
.Y(n_3861)
);

NOR2xp33_ASAP7_75t_L g3862 ( 
.A(n_3646),
.B(n_3022),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3576),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3476),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3480),
.Y(n_3865)
);

BUFx3_ASAP7_75t_L g3866 ( 
.A(n_3503),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3481),
.Y(n_3867)
);

AOI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3452),
.A2(n_3561),
.B1(n_3432),
.B2(n_3477),
.Y(n_3868)
);

INVxp67_ASAP7_75t_L g3869 ( 
.A(n_3451),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3484),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3493),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3577),
.Y(n_3872)
);

BUFx2_ASAP7_75t_L g3873 ( 
.A(n_3571),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3580),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3588),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3601),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3627),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3640),
.Y(n_3878)
);

INVxp67_ASAP7_75t_L g3879 ( 
.A(n_3571),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3403),
.B(n_3267),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3582),
.Y(n_3881)
);

INVx3_ASAP7_75t_L g3882 ( 
.A(n_3399),
.Y(n_3882)
);

AND2x4_ASAP7_75t_L g3883 ( 
.A(n_3386),
.B(n_2925),
.Y(n_3883)
);

NOR2xp33_ASAP7_75t_L g3884 ( 
.A(n_3646),
.B(n_3022),
.Y(n_3884)
);

OR2x6_ASAP7_75t_L g3885 ( 
.A(n_3423),
.B(n_3253),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3583),
.Y(n_3886)
);

NOR2xp33_ASAP7_75t_L g3887 ( 
.A(n_3656),
.B(n_3700),
.Y(n_3887)
);

AOI22xp33_ASAP7_75t_L g3888 ( 
.A1(n_3452),
.A2(n_2936),
.B1(n_3246),
.B2(n_3217),
.Y(n_3888)
);

NAND3xp33_ASAP7_75t_L g3889 ( 
.A(n_3406),
.B(n_3281),
.C(n_3275),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3585),
.Y(n_3890)
);

AOI22xp33_ASAP7_75t_L g3891 ( 
.A1(n_3561),
.A2(n_2936),
.B1(n_3290),
.B2(n_3257),
.Y(n_3891)
);

INVx3_ASAP7_75t_L g3892 ( 
.A(n_3675),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3655),
.Y(n_3893)
);

NOR2x1p5_ASAP7_75t_L g3894 ( 
.A(n_3704),
.B(n_2995),
.Y(n_3894)
);

BUFx6f_ASAP7_75t_L g3895 ( 
.A(n_3468),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3502),
.B(n_3039),
.Y(n_3896)
);

INVxp67_ASAP7_75t_L g3897 ( 
.A(n_3631),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3514),
.B(n_3039),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3589),
.Y(n_3899)
);

INVx3_ASAP7_75t_L g3900 ( 
.A(n_3675),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3593),
.Y(n_3901)
);

AOI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3525),
.A2(n_2936),
.B1(n_3327),
.B2(n_3311),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3515),
.B(n_3508),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3603),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3432),
.A2(n_3311),
.B1(n_1160),
.B2(n_1242),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3606),
.Y(n_3906)
);

OAI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3390),
.A2(n_3341),
.B1(n_1082),
.B2(n_1242),
.Y(n_3907)
);

AND2x4_ASAP7_75t_L g3908 ( 
.A(n_3386),
.B(n_2925),
.Y(n_3908)
);

AOI22xp5_ASAP7_75t_L g3909 ( 
.A1(n_3543),
.A2(n_3205),
.B1(n_3237),
.B2(n_3201),
.Y(n_3909)
);

AND2x6_ASAP7_75t_SL g3910 ( 
.A(n_3615),
.B(n_736),
.Y(n_3910)
);

NOR2xp33_ASAP7_75t_L g3911 ( 
.A(n_3708),
.B(n_3056),
.Y(n_3911)
);

AOI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3653),
.A2(n_3201),
.B1(n_3237),
.B2(n_3205),
.Y(n_3912)
);

AOI22xp33_ASAP7_75t_L g3913 ( 
.A1(n_3477),
.A2(n_1160),
.B1(n_3312),
.B2(n_3040),
.Y(n_3913)
);

A2O1A1Ixp33_ASAP7_75t_L g3914 ( 
.A1(n_3708),
.A2(n_3462),
.B(n_3567),
.C(n_3722),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3615),
.B(n_3413),
.Y(n_3915)
);

INVx3_ASAP7_75t_L g3916 ( 
.A(n_3492),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3509),
.B(n_3312),
.Y(n_3917)
);

BUFx3_ASAP7_75t_L g3918 ( 
.A(n_3503),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3609),
.Y(n_3919)
);

AOI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3653),
.A2(n_3341),
.B1(n_3267),
.B2(n_3276),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_SL g3921 ( 
.A(n_3669),
.B(n_3510),
.Y(n_3921)
);

OR2x2_ASAP7_75t_L g3922 ( 
.A(n_3701),
.B(n_3276),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3614),
.A2(n_3341),
.B(n_3247),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3510),
.B(n_2981),
.Y(n_3924)
);

BUFx6f_ASAP7_75t_L g3925 ( 
.A(n_3492),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3396),
.B(n_3329),
.Y(n_3926)
);

INVx3_ASAP7_75t_L g3927 ( 
.A(n_3492),
.Y(n_3927)
);

CKINVDCx5p33_ASAP7_75t_R g3928 ( 
.A(n_3454),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_SL g3929 ( 
.A(n_3518),
.B(n_2981),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_3456),
.A2(n_3064),
.B(n_2967),
.Y(n_3930)
);

OAI22xp5_ASAP7_75t_L g3931 ( 
.A1(n_3409),
.A2(n_3068),
.B1(n_2981),
.B2(n_3108),
.Y(n_3931)
);

INVx2_ASAP7_75t_SL g3932 ( 
.A(n_3648),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3611),
.Y(n_3933)
);

AND2x4_ASAP7_75t_L g3934 ( 
.A(n_3714),
.B(n_2931),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3419),
.B(n_3294),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3616),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3667),
.Y(n_3937)
);

NOR2xp33_ASAP7_75t_L g3938 ( 
.A(n_3591),
.B(n_3294),
.Y(n_3938)
);

INVxp67_ASAP7_75t_SL g3939 ( 
.A(n_3586),
.Y(n_3939)
);

INVx1_ASAP7_75t_SL g3940 ( 
.A(n_3728),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3420),
.B(n_3294),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3619),
.Y(n_3942)
);

HB1xp67_ASAP7_75t_L g3943 ( 
.A(n_3555),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3671),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3391),
.B(n_3197),
.Y(n_3945)
);

HB1xp67_ASAP7_75t_L g3946 ( 
.A(n_3555),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3506),
.B(n_2995),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3387),
.B(n_3035),
.Y(n_3948)
);

INVxp67_ASAP7_75t_L g3949 ( 
.A(n_3631),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3676),
.B(n_3035),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3674),
.Y(n_3951)
);

INVx5_ASAP7_75t_L g3952 ( 
.A(n_3513),
.Y(n_3952)
);

INVx3_ASAP7_75t_L g3953 ( 
.A(n_3492),
.Y(n_3953)
);

BUFx6f_ASAP7_75t_L g3954 ( 
.A(n_3497),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3447),
.B(n_3042),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3681),
.Y(n_3956)
);

INVx1_ASAP7_75t_SL g3957 ( 
.A(n_3719),
.Y(n_3957)
);

OR2x6_ASAP7_75t_L g3958 ( 
.A(n_3513),
.B(n_2931),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3459),
.A2(n_3411),
.B1(n_3418),
.B2(n_3557),
.Y(n_3959)
);

OR2x6_ASAP7_75t_L g3960 ( 
.A(n_3513),
.B(n_2933),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3622),
.Y(n_3961)
);

AND2x4_ASAP7_75t_L g3962 ( 
.A(n_3714),
.B(n_2933),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3623),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3628),
.Y(n_3964)
);

BUFx3_ASAP7_75t_L g3965 ( 
.A(n_3662),
.Y(n_3965)
);

OR2x2_ASAP7_75t_L g3966 ( 
.A(n_3641),
.B(n_2268),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3630),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3632),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3687),
.Y(n_3969)
);

NOR2xp33_ASAP7_75t_L g3970 ( 
.A(n_3592),
.B(n_3243),
.Y(n_3970)
);

NOR2xp33_ASAP7_75t_L g3971 ( 
.A(n_3660),
.B(n_3243),
.Y(n_3971)
);

OR2x2_ASAP7_75t_L g3972 ( 
.A(n_3719),
.B(n_2268),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3489),
.B(n_3040),
.Y(n_3973)
);

INVx4_ASAP7_75t_L g3974 ( 
.A(n_3444),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3635),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3491),
.B(n_3042),
.Y(n_3976)
);

CKINVDCx5p33_ASAP7_75t_R g3977 ( 
.A(n_3612),
.Y(n_3977)
);

NAND2x1p5_ASAP7_75t_L g3978 ( 
.A(n_3662),
.B(n_2983),
.Y(n_3978)
);

NOR2xp33_ASAP7_75t_L g3979 ( 
.A(n_3661),
.B(n_3153),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3411),
.A2(n_3557),
.B1(n_3549),
.B2(n_3552),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3645),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3691),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_SL g3983 ( 
.A(n_3518),
.B(n_3068),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3650),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3672),
.Y(n_3985)
);

NOR2xp33_ASAP7_75t_SL g3986 ( 
.A(n_3517),
.B(n_3098),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3673),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3499),
.B(n_3045),
.Y(n_3988)
);

BUFx6f_ASAP7_75t_SL g3989 ( 
.A(n_3444),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3698),
.Y(n_3990)
);

A2O1A1Ixp33_ASAP7_75t_L g3991 ( 
.A1(n_3512),
.A2(n_3048),
.B(n_3124),
.C(n_3045),
.Y(n_3991)
);

AOI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3634),
.A2(n_3180),
.B1(n_3160),
.B2(n_3027),
.Y(n_3992)
);

INVx1_ASAP7_75t_SL g3993 ( 
.A(n_3766),
.Y(n_3993)
);

INVx2_ASAP7_75t_SL g3994 ( 
.A(n_3766),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3469),
.B(n_883),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3680),
.Y(n_3996)
);

INVx3_ASAP7_75t_L g3997 ( 
.A(n_3497),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3705),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3731),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3500),
.B(n_3048),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3694),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3549),
.A2(n_3129),
.B1(n_3131),
.B2(n_3124),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3739),
.Y(n_4003)
);

NOR2xp33_ASAP7_75t_L g4004 ( 
.A(n_3537),
.B(n_3169),
.Y(n_4004)
);

AOI22xp33_ASAP7_75t_L g4005 ( 
.A1(n_3570),
.A2(n_3131),
.B1(n_3133),
.B2(n_3129),
.Y(n_4005)
);

AND2x4_ASAP7_75t_L g4006 ( 
.A(n_3718),
.B(n_2920),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3771),
.Y(n_4007)
);

AOI22xp5_ASAP7_75t_L g4008 ( 
.A1(n_3534),
.A2(n_3027),
.B1(n_3041),
.B2(n_2953),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3466),
.B(n_3133),
.Y(n_4009)
);

BUFx8_ASAP7_75t_L g4010 ( 
.A(n_3612),
.Y(n_4010)
);

INVx2_ASAP7_75t_L g4011 ( 
.A(n_3776),
.Y(n_4011)
);

AOI22xp5_ASAP7_75t_L g4012 ( 
.A1(n_3597),
.A2(n_3041),
.B1(n_3070),
.B2(n_3027),
.Y(n_4012)
);

CKINVDCx5p33_ASAP7_75t_R g4013 ( 
.A(n_3504),
.Y(n_4013)
);

INVx2_ASAP7_75t_SL g4014 ( 
.A(n_3412),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_SL g4015 ( 
.A(n_3518),
.B(n_3068),
.Y(n_4015)
);

BUFx12f_ASAP7_75t_L g4016 ( 
.A(n_3439),
.Y(n_4016)
);

NAND2x1p5_ASAP7_75t_L g4017 ( 
.A(n_3497),
.B(n_2983),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_SL g4018 ( 
.A(n_3518),
.B(n_2964),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3707),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3711),
.Y(n_4020)
);

AND2x2_ASAP7_75t_SL g4021 ( 
.A(n_3696),
.B(n_2983),
.Y(n_4021)
);

NOR2xp33_ASAP7_75t_L g4022 ( 
.A(n_3523),
.B(n_3169),
.Y(n_4022)
);

BUFx6f_ASAP7_75t_L g4023 ( 
.A(n_3497),
.Y(n_4023)
);

INVx2_ASAP7_75t_SL g4024 ( 
.A(n_3453),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3713),
.Y(n_4025)
);

INVx2_ASAP7_75t_SL g4026 ( 
.A(n_3658),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3725),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3744),
.Y(n_4028)
);

NAND2xp33_ASAP7_75t_L g4029 ( 
.A(n_3518),
.B(n_3027),
.Y(n_4029)
);

OR2x2_ASAP7_75t_SL g4030 ( 
.A(n_3448),
.B(n_3556),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3478),
.B(n_3202),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3529),
.B(n_3202),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_SL g4033 ( 
.A(n_3518),
.B(n_2964),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3450),
.B(n_3204),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_SL g4035 ( 
.A(n_3605),
.B(n_2964),
.Y(n_4035)
);

AND2x4_ASAP7_75t_L g4036 ( 
.A(n_3718),
.B(n_2920),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_3540),
.B(n_2964),
.Y(n_4037)
);

CKINVDCx5p33_ASAP7_75t_R g4038 ( 
.A(n_3541),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3471),
.B(n_883),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3747),
.Y(n_4040)
);

INVx8_ASAP7_75t_L g4041 ( 
.A(n_3764),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3754),
.Y(n_4042)
);

NOR2xp33_ASAP7_75t_L g4043 ( 
.A(n_3415),
.B(n_3204),
.Y(n_4043)
);

HB1xp67_ASAP7_75t_L g4044 ( 
.A(n_3575),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3496),
.B(n_919),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3755),
.Y(n_4046)
);

NOR2xp33_ASAP7_75t_L g4047 ( 
.A(n_3522),
.B(n_3208),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3759),
.Y(n_4048)
);

NOR2x1p5_ASAP7_75t_L g4049 ( 
.A(n_3618),
.B(n_2256),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3760),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3767),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3769),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3723),
.Y(n_4053)
);

AND2x4_ASAP7_75t_L g4054 ( 
.A(n_3624),
.B(n_2920),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3738),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3457),
.B(n_3208),
.Y(n_4056)
);

INVx5_ASAP7_75t_L g4057 ( 
.A(n_3524),
.Y(n_4057)
);

OR2x2_ASAP7_75t_L g4058 ( 
.A(n_3608),
.B(n_2277),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3421),
.B(n_3212),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3551),
.Y(n_4060)
);

BUFx3_ASAP7_75t_L g4061 ( 
.A(n_3764),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3553),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3597),
.B(n_3212),
.Y(n_4063)
);

OR2x2_ASAP7_75t_L g4064 ( 
.A(n_3613),
.B(n_2277),
.Y(n_4064)
);

AND2x4_ASAP7_75t_SL g4065 ( 
.A(n_3764),
.B(n_3098),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_L g4066 ( 
.A(n_3620),
.B(n_3230),
.Y(n_4066)
);

INVx5_ASAP7_75t_L g4067 ( 
.A(n_3524),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3742),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3443),
.Y(n_4069)
);

AND2x4_ASAP7_75t_L g4070 ( 
.A(n_3629),
.B(n_2920),
.Y(n_4070)
);

NOR2xp33_ASAP7_75t_R g4071 ( 
.A(n_3578),
.B(n_3098),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3604),
.B(n_3230),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3445),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3743),
.Y(n_4074)
);

INVx5_ASAP7_75t_L g4075 ( 
.A(n_3524),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3604),
.B(n_3235),
.Y(n_4076)
);

INVx4_ASAP7_75t_L g4077 ( 
.A(n_3524),
.Y(n_4077)
);

AND2x4_ASAP7_75t_L g4078 ( 
.A(n_3638),
.B(n_3030),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_SL g4079 ( 
.A(n_3559),
.B(n_2964),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3397),
.Y(n_4080)
);

BUFx6f_ASAP7_75t_L g4081 ( 
.A(n_3538),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_3748),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3749),
.Y(n_4083)
);

INVxp67_ASAP7_75t_L g4084 ( 
.A(n_3777),
.Y(n_4084)
);

INVx4_ASAP7_75t_L g4085 ( 
.A(n_3538),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3505),
.B(n_3235),
.Y(n_4086)
);

AND2x4_ASAP7_75t_L g4087 ( 
.A(n_3598),
.B(n_3030),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3402),
.Y(n_4088)
);

BUFx6f_ASAP7_75t_L g4089 ( 
.A(n_3538),
.Y(n_4089)
);

AND2x4_ASAP7_75t_L g4090 ( 
.A(n_3600),
.B(n_3030),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_SL g4091 ( 
.A(n_3512),
.B(n_2976),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3533),
.B(n_3240),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3535),
.B(n_3240),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3715),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3486),
.B(n_3248),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3716),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_3575),
.B(n_919),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3751),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3486),
.B(n_3248),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3490),
.B(n_3307),
.Y(n_4100)
);

CKINVDCx5p33_ASAP7_75t_R g4101 ( 
.A(n_3610),
.Y(n_4101)
);

A2O1A1Ixp33_ASAP7_75t_L g4102 ( 
.A1(n_3568),
.A2(n_3381),
.B(n_3384),
.C(n_3307),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3717),
.Y(n_4103)
);

A2O1A1Ixp33_ASAP7_75t_L g4104 ( 
.A1(n_3568),
.A2(n_3384),
.B(n_3385),
.C(n_3381),
.Y(n_4104)
);

INVx5_ASAP7_75t_L g4105 ( 
.A(n_3538),
.Y(n_4105)
);

BUFx3_ASAP7_75t_L g4106 ( 
.A(n_3566),
.Y(n_4106)
);

BUFx3_ASAP7_75t_L g4107 ( 
.A(n_3746),
.Y(n_4107)
);

INVx3_ASAP7_75t_L g4108 ( 
.A(n_3482),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3721),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3729),
.Y(n_4110)
);

INVx3_ASAP7_75t_L g4111 ( 
.A(n_3482),
.Y(n_4111)
);

NOR2xp33_ASAP7_75t_L g4112 ( 
.A(n_3434),
.B(n_3385),
.Y(n_4112)
);

INVx2_ASAP7_75t_SL g4113 ( 
.A(n_3658),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_3490),
.B(n_2256),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_SL g4115 ( 
.A(n_3770),
.B(n_2976),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3581),
.B(n_2256),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_3775),
.B(n_2976),
.Y(n_4117)
);

A2O1A1Ixp33_ASAP7_75t_L g4118 ( 
.A1(n_3587),
.A2(n_2717),
.B(n_2725),
.C(n_2718),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_3649),
.B(n_3030),
.Y(n_4119)
);

AOI21xp5_ASAP7_75t_L g4120 ( 
.A1(n_3550),
.A2(n_3089),
.B(n_3087),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_3753),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3777),
.B(n_2265),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3724),
.A2(n_3364),
.B(n_3293),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3531),
.B(n_2976),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3781),
.B(n_2265),
.Y(n_4125)
);

INVx3_ASAP7_75t_L g4126 ( 
.A(n_3536),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3781),
.B(n_2265),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3752),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3752),
.Y(n_4129)
);

OR2x2_ASAP7_75t_SL g4130 ( 
.A(n_3595),
.B(n_756),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3425),
.B(n_2267),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_3464),
.B(n_3156),
.Y(n_4132)
);

INVx2_ASAP7_75t_SL g4133 ( 
.A(n_3520),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3429),
.B(n_3430),
.Y(n_4134)
);

AOI22xp33_ASAP7_75t_L g4135 ( 
.A1(n_3436),
.A2(n_2283),
.B1(n_2285),
.B2(n_2278),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_SL g4136 ( 
.A(n_3542),
.B(n_2976),
.Y(n_4136)
);

INVxp67_ASAP7_75t_L g4137 ( 
.A(n_3686),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3668),
.B(n_3663),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3682),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3664),
.B(n_2267),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3539),
.B(n_2267),
.Y(n_4141)
);

NOR2xp33_ASAP7_75t_L g4142 ( 
.A(n_3644),
.B(n_2298),
.Y(n_4142)
);

BUFx2_ASAP7_75t_L g4143 ( 
.A(n_3573),
.Y(n_4143)
);

NOR2xp33_ASAP7_75t_R g4144 ( 
.A(n_3574),
.B(n_3219),
.Y(n_4144)
);

INVx5_ASAP7_75t_L g4145 ( 
.A(n_3746),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3756),
.Y(n_4146)
);

BUFx3_ASAP7_75t_L g4147 ( 
.A(n_3746),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_3564),
.B(n_919),
.Y(n_4148)
);

BUFx2_ASAP7_75t_L g4149 ( 
.A(n_3610),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3683),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3545),
.B(n_2987),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3569),
.B(n_2298),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3688),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3695),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3709),
.Y(n_4155)
);

BUFx6f_ASAP7_75t_L g4156 ( 
.A(n_3746),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_3758),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3710),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_3763),
.Y(n_4159)
);

OAI22xp33_ASAP7_75t_L g4160 ( 
.A1(n_3678),
.A2(n_1084),
.B1(n_1102),
.B2(n_1070),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3887),
.B(n_3686),
.Y(n_4161)
);

NAND2xp33_ASAP7_75t_SL g4162 ( 
.A(n_3849),
.B(n_3546),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3887),
.B(n_3474),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_SL g4164 ( 
.A(n_3846),
.B(n_3726),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_SL g4165 ( 
.A(n_3847),
.B(n_3761),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_SL g4166 ( 
.A(n_3845),
.B(n_3772),
.Y(n_4166)
);

NAND2xp33_ASAP7_75t_SL g4167 ( 
.A(n_3844),
.B(n_4071),
.Y(n_4167)
);

AND2x2_ASAP7_75t_L g4168 ( 
.A(n_3868),
.B(n_3774),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_SL g4169 ( 
.A(n_3915),
.B(n_3772),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_SL g4170 ( 
.A(n_3903),
.B(n_3772),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_SL g4171 ( 
.A(n_3793),
.B(n_3772),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_3850),
.B(n_3410),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3796),
.B(n_3690),
.Y(n_4173)
);

NAND2xp33_ASAP7_75t_SL g4174 ( 
.A(n_3844),
.B(n_3657),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3914),
.B(n_3732),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3914),
.B(n_3736),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_SL g4177 ( 
.A(n_3801),
.B(n_3730),
.Y(n_4177)
);

NAND2xp33_ASAP7_75t_SL g4178 ( 
.A(n_4071),
.B(n_3657),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_SL g4179 ( 
.A(n_3911),
.B(n_3730),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_SL g4180 ( 
.A(n_3911),
.B(n_3498),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_4094),
.B(n_3735),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4096),
.B(n_4103),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_4109),
.B(n_3735),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_SL g4184 ( 
.A(n_4137),
.B(n_3633),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_SL g4185 ( 
.A(n_4137),
.B(n_3852),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_SL g4186 ( 
.A(n_3862),
.B(n_3884),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_SL g4187 ( 
.A(n_3862),
.B(n_3643),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_3868),
.B(n_3757),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_SL g4189 ( 
.A(n_3884),
.B(n_3637),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_SL g4190 ( 
.A(n_3823),
.B(n_3734),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_4112),
.B(n_3734),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_SL g4192 ( 
.A(n_4112),
.B(n_3727),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_SL g4193 ( 
.A(n_3837),
.B(n_3727),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_SL g4194 ( 
.A(n_3838),
.B(n_3572),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4110),
.B(n_3679),
.Y(n_4195)
);

NAND2xp33_ASAP7_75t_SL g4196 ( 
.A(n_3843),
.B(n_3697),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_4053),
.B(n_4060),
.Y(n_4197)
);

OR2x2_ASAP7_75t_L g4198 ( 
.A(n_3943),
.B(n_3654),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_SL g4199 ( 
.A(n_3907),
.B(n_3677),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_SL g4200 ( 
.A(n_3907),
.B(n_3579),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_SL g4201 ( 
.A(n_3854),
.B(n_3896),
.Y(n_4201)
);

NAND2xp33_ASAP7_75t_SL g4202 ( 
.A(n_4026),
.B(n_3699),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_SL g4203 ( 
.A(n_3986),
.B(n_3599),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_SL g4204 ( 
.A(n_3920),
.B(n_3626),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_SL g4205 ( 
.A(n_3820),
.B(n_3684),
.Y(n_4205)
);

NAND2xp33_ASAP7_75t_SL g4206 ( 
.A(n_4113),
.B(n_3703),
.Y(n_4206)
);

AND2x4_ASAP7_75t_L g4207 ( 
.A(n_3831),
.B(n_3156),
.Y(n_4207)
);

NAND2xp33_ASAP7_75t_SL g4208 ( 
.A(n_3974),
.B(n_3536),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_3943),
.B(n_3757),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_SL g4210 ( 
.A(n_3807),
.B(n_3813),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_3946),
.B(n_3507),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_SL g4212 ( 
.A(n_4084),
.B(n_3712),
.Y(n_4212)
);

NAND2xp33_ASAP7_75t_SL g4213 ( 
.A(n_3974),
.B(n_3670),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_SL g4214 ( 
.A(n_4084),
.B(n_3768),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4062),
.B(n_3596),
.Y(n_4215)
);

NAND2xp33_ASAP7_75t_SL g4216 ( 
.A(n_3989),
.B(n_3670),
.Y(n_4216)
);

NAND2xp33_ASAP7_75t_SL g4217 ( 
.A(n_3989),
.B(n_3689),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_SL g4218 ( 
.A(n_4138),
.B(n_3690),
.Y(n_4218)
);

NAND2xp33_ASAP7_75t_SL g4219 ( 
.A(n_3824),
.B(n_3689),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_SL g4220 ( 
.A(n_3825),
.B(n_2987),
.Y(n_4220)
);

AND2x4_ASAP7_75t_L g4221 ( 
.A(n_3831),
.B(n_3156),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_SL g4222 ( 
.A(n_3815),
.B(n_2987),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_3816),
.B(n_2987),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_SL g4224 ( 
.A(n_4095),
.B(n_2987),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_SL g4225 ( 
.A(n_4099),
.B(n_3036),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_4100),
.B(n_3036),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3794),
.B(n_3926),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_SL g4228 ( 
.A(n_3947),
.B(n_3036),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_SL g4229 ( 
.A(n_4114),
.B(n_3036),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_3804),
.B(n_3036),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_SL g4231 ( 
.A(n_3830),
.B(n_3097),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_3830),
.B(n_3097),
.Y(n_4232)
);

NAND2xp33_ASAP7_75t_SL g4233 ( 
.A(n_3824),
.B(n_3702),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_SL g4234 ( 
.A(n_3898),
.B(n_3097),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_SL g4235 ( 
.A(n_3902),
.B(n_3097),
.Y(n_4235)
);

NAND2xp33_ASAP7_75t_SL g4236 ( 
.A(n_3828),
.B(n_3702),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_SL g4237 ( 
.A(n_3935),
.B(n_3097),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_SL g4238 ( 
.A(n_3941),
.B(n_3112),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_SL g4239 ( 
.A(n_4013),
.B(n_3112),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_3827),
.B(n_3636),
.Y(n_4240)
);

AND2x4_ASAP7_75t_L g4241 ( 
.A(n_3836),
.B(n_3156),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_SL g4242 ( 
.A(n_4063),
.B(n_3112),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_SL g4243 ( 
.A(n_4072),
.B(n_3112),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_4076),
.B(n_3112),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_3957),
.B(n_3651),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_SL g4246 ( 
.A(n_4139),
.B(n_3778),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_SL g4247 ( 
.A(n_4150),
.B(n_3779),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_SL g4248 ( 
.A(n_4153),
.B(n_3780),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_SL g4249 ( 
.A(n_4154),
.B(n_3142),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_3993),
.B(n_3652),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_SL g4251 ( 
.A(n_4155),
.B(n_3163),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_4158),
.B(n_3163),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_SL g4253 ( 
.A(n_4021),
.B(n_3992),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_SL g4254 ( 
.A(n_4021),
.B(n_3163),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_SL g4255 ( 
.A(n_4022),
.B(n_3163),
.Y(n_4255)
);

NAND2xp33_ASAP7_75t_SL g4256 ( 
.A(n_4101),
.B(n_3733),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4080),
.B(n_3782),
.Y(n_4257)
);

NAND2xp33_ASAP7_75t_SL g4258 ( 
.A(n_3817),
.B(n_3733),
.Y(n_4258)
);

NAND2xp33_ASAP7_75t_SL g4259 ( 
.A(n_3836),
.B(n_3163),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_SL g4260 ( 
.A(n_4022),
.B(n_3173),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_SL g4261 ( 
.A(n_4122),
.B(n_3173),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_SL g4262 ( 
.A(n_4125),
.B(n_3173),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_SL g4263 ( 
.A(n_4127),
.B(n_3173),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_3946),
.B(n_4046),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_SL g4265 ( 
.A(n_4066),
.B(n_3173),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_SL g4266 ( 
.A(n_4066),
.B(n_3188),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_SL g4267 ( 
.A(n_3806),
.B(n_3188),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_SL g4268 ( 
.A(n_3945),
.B(n_3188),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_SL g4269 ( 
.A(n_4134),
.B(n_3188),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_SL g4270 ( 
.A(n_4142),
.B(n_3188),
.Y(n_4270)
);

AND2x2_ASAP7_75t_L g4271 ( 
.A(n_4042),
.B(n_3594),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_SL g4272 ( 
.A(n_4142),
.B(n_3213),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4088),
.B(n_2278),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_SL g4274 ( 
.A(n_3811),
.B(n_3829),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_SL g4275 ( 
.A(n_3811),
.B(n_3213),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_3829),
.B(n_3213),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_SL g4277 ( 
.A(n_3882),
.B(n_3213),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_3882),
.B(n_3213),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_SL g4279 ( 
.A(n_4038),
.B(n_3223),
.Y(n_4279)
);

NAND2xp33_ASAP7_75t_SL g4280 ( 
.A(n_4144),
.B(n_3223),
.Y(n_4280)
);

NAND2xp33_ASAP7_75t_SL g4281 ( 
.A(n_4144),
.B(n_3223),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_SL g4282 ( 
.A(n_3797),
.B(n_3912),
.Y(n_4282)
);

NAND2xp33_ASAP7_75t_SL g4283 ( 
.A(n_4092),
.B(n_3223),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_4107),
.B(n_4147),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_SL g4285 ( 
.A(n_3797),
.B(n_3223),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_4069),
.B(n_2283),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_SL g4287 ( 
.A(n_4009),
.B(n_3251),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_4073),
.B(n_2285),
.Y(n_4288)
);

NAND2xp33_ASAP7_75t_SL g4289 ( 
.A(n_4093),
.B(n_4149),
.Y(n_4289)
);

NAND2xp33_ASAP7_75t_SL g4290 ( 
.A(n_3994),
.B(n_3251),
.Y(n_4290)
);

NAND2xp33_ASAP7_75t_SL g4291 ( 
.A(n_4031),
.B(n_3251),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_4044),
.B(n_2293),
.Y(n_4292)
);

AND2x4_ASAP7_75t_L g4293 ( 
.A(n_4107),
.B(n_3209),
.Y(n_4293)
);

AND2x4_ASAP7_75t_L g4294 ( 
.A(n_4147),
.B(n_3209),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_SL g4295 ( 
.A(n_4056),
.B(n_3251),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_SL g4296 ( 
.A(n_3892),
.B(n_3251),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_SL g4297 ( 
.A(n_3892),
.B(n_3277),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_SL g4298 ( 
.A(n_3900),
.B(n_3277),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_SL g4299 ( 
.A(n_3900),
.B(n_3277),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_SL g4300 ( 
.A(n_3921),
.B(n_3277),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_SL g4301 ( 
.A(n_3921),
.B(n_3277),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_SL g4302 ( 
.A(n_4032),
.B(n_3296),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_SL g4303 ( 
.A(n_3866),
.B(n_3296),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_SL g4304 ( 
.A(n_3866),
.B(n_3296),
.Y(n_4304)
);

AND2x4_ASAP7_75t_L g4305 ( 
.A(n_4145),
.B(n_3209),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_SL g4306 ( 
.A(n_3918),
.B(n_3296),
.Y(n_4306)
);

NAND2xp33_ASAP7_75t_SL g4307 ( 
.A(n_4034),
.B(n_3296),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_SL g4308 ( 
.A(n_3918),
.B(n_3301),
.Y(n_4308)
);

NAND2xp33_ASAP7_75t_SL g4309 ( 
.A(n_3873),
.B(n_3803),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_SL g4310 ( 
.A(n_3965),
.B(n_3301),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_SL g4311 ( 
.A(n_3965),
.B(n_3301),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4044),
.B(n_2293),
.Y(n_4312)
);

NAND2xp33_ASAP7_75t_SL g4313 ( 
.A(n_4049),
.B(n_3973),
.Y(n_4313)
);

AND2x2_ASAP7_75t_SL g4314 ( 
.A(n_3891),
.B(n_3765),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_SL g4315 ( 
.A(n_4070),
.B(n_3301),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_SL g4316 ( 
.A(n_4070),
.B(n_3301),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4078),
.B(n_3340),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_SL g4318 ( 
.A(n_4078),
.B(n_3340),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_3821),
.B(n_2295),
.Y(n_4319)
);

AND2x2_ASAP7_75t_L g4320 ( 
.A(n_4048),
.B(n_3750),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_SL g4321 ( 
.A(n_4008),
.B(n_3938),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_SL g4322 ( 
.A(n_3938),
.B(n_4057),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_SL g4323 ( 
.A(n_4057),
.B(n_3340),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_SL g4324 ( 
.A(n_4057),
.B(n_3340),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_SL g4325 ( 
.A(n_4057),
.B(n_3340),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_4067),
.B(n_4075),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_SL g4327 ( 
.A(n_4067),
.B(n_3375),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_SL g4328 ( 
.A(n_4067),
.B(n_3375),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_SL g4329 ( 
.A(n_4067),
.B(n_3375),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_SL g4330 ( 
.A(n_4075),
.B(n_3375),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_SL g4331 ( 
.A(n_4075),
.B(n_3375),
.Y(n_4331)
);

AND2x4_ASAP7_75t_L g4332 ( 
.A(n_4145),
.B(n_3209),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_SL g4333 ( 
.A(n_4075),
.B(n_3322),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_SL g4334 ( 
.A(n_4105),
.B(n_3322),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_SL g4335 ( 
.A(n_4105),
.B(n_4087),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_SL g4336 ( 
.A(n_4105),
.B(n_3322),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_SL g4337 ( 
.A(n_4105),
.B(n_3322),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_SL g4338 ( 
.A(n_4087),
.B(n_3322),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_SL g4339 ( 
.A(n_4090),
.B(n_3219),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_4090),
.B(n_3219),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_3821),
.B(n_3869),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_3869),
.B(n_2295),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_SL g4343 ( 
.A(n_3971),
.B(n_4141),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_3879),
.B(n_3378),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_SL g4345 ( 
.A(n_3971),
.B(n_3879),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_SL g4346 ( 
.A(n_3897),
.B(n_3234),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_SL g4347 ( 
.A(n_3897),
.B(n_3234),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_SL g4348 ( 
.A(n_3949),
.B(n_3234),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_SL g4349 ( 
.A(n_3949),
.B(n_3067),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_3940),
.B(n_3378),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_SL g4351 ( 
.A(n_4004),
.B(n_3067),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4055),
.B(n_3378),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4068),
.B(n_3378),
.Y(n_4353)
);

AND2x4_ASAP7_75t_L g4354 ( 
.A(n_4145),
.B(n_3233),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_SL g4355 ( 
.A(n_4004),
.B(n_3067),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_SL g4356 ( 
.A(n_3976),
.B(n_3093),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_SL g4357 ( 
.A(n_3988),
.B(n_3093),
.Y(n_4357)
);

NAND2xp33_ASAP7_75t_SL g4358 ( 
.A(n_4000),
.B(n_3093),
.Y(n_4358)
);

NAND2xp33_ASAP7_75t_SL g4359 ( 
.A(n_3950),
.B(n_3114),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_SL g4360 ( 
.A(n_4152),
.B(n_3114),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_SL g4361 ( 
.A(n_4054),
.B(n_3114),
.Y(n_4361)
);

NAND2xp33_ASAP7_75t_SL g4362 ( 
.A(n_3955),
.B(n_3128),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_SL g4363 ( 
.A(n_4054),
.B(n_3970),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_SL g4364 ( 
.A(n_3970),
.B(n_3128),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_SL g4365 ( 
.A(n_4043),
.B(n_3128),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4074),
.B(n_3378),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_SL g4367 ( 
.A(n_4043),
.B(n_3236),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4050),
.B(n_3750),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_SL g4369 ( 
.A(n_4047),
.B(n_3236),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_SL g4370 ( 
.A(n_4047),
.B(n_3236),
.Y(n_4370)
);

NAND2xp33_ASAP7_75t_SL g4371 ( 
.A(n_3818),
.B(n_3441),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_SL g4372 ( 
.A(n_4145),
.B(n_3295),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_SL g4373 ( 
.A(n_4132),
.B(n_3295),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_SL g4374 ( 
.A(n_4132),
.B(n_3295),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_SL g4375 ( 
.A(n_3934),
.B(n_3299),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_SL g4376 ( 
.A(n_3934),
.B(n_3299),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_4082),
.B(n_3378),
.Y(n_4377)
);

NAND2xp33_ASAP7_75t_SL g4378 ( 
.A(n_3832),
.B(n_3441),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_SL g4379 ( 
.A(n_3962),
.B(n_3299),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_SL g4380 ( 
.A(n_3962),
.B(n_4059),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_SL g4381 ( 
.A(n_3785),
.B(n_3317),
.Y(n_4381)
);

NAND2xp33_ASAP7_75t_SL g4382 ( 
.A(n_4140),
.B(n_3642),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_SL g4383 ( 
.A(n_3785),
.B(n_3317),
.Y(n_4383)
);

NAND2xp33_ASAP7_75t_SL g4384 ( 
.A(n_4116),
.B(n_3642),
.Y(n_4384)
);

NAND2xp33_ASAP7_75t_SL g4385 ( 
.A(n_3799),
.B(n_3308),
.Y(n_4385)
);

AND2x4_ASAP7_75t_L g4386 ( 
.A(n_4006),
.B(n_4036),
.Y(n_4386)
);

NAND2xp33_ASAP7_75t_SL g4387 ( 
.A(n_4108),
.B(n_4111),
.Y(n_4387)
);

NAND2xp33_ASAP7_75t_SL g4388 ( 
.A(n_4108),
.B(n_3314),
.Y(n_4388)
);

AND3x1_ASAP7_75t_L g4389 ( 
.A(n_3909),
.B(n_737),
.C(n_736),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_SL g4390 ( 
.A(n_3785),
.B(n_3317),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_SL g4391 ( 
.A(n_3785),
.B(n_3325),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_SL g4392 ( 
.A(n_3786),
.B(n_3325),
.Y(n_4392)
);

NAND2xp33_ASAP7_75t_SL g4393 ( 
.A(n_4111),
.B(n_3330),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_SL g4394 ( 
.A(n_3786),
.B(n_3325),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_SL g4395 ( 
.A(n_3786),
.B(n_3336),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_SL g4396 ( 
.A(n_3786),
.B(n_3336),
.Y(n_4396)
);

OR2x2_ASAP7_75t_L g4397 ( 
.A(n_3972),
.B(n_3528),
.Y(n_4397)
);

NAND2xp33_ASAP7_75t_SL g4398 ( 
.A(n_4126),
.B(n_3334),
.Y(n_4398)
);

NAND2xp33_ASAP7_75t_SL g4399 ( 
.A(n_4126),
.B(n_3339),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_SL g4400 ( 
.A(n_3895),
.B(n_3336),
.Y(n_4400)
);

NAND2xp33_ASAP7_75t_SL g4401 ( 
.A(n_4133),
.B(n_3894),
.Y(n_4401)
);

AND2x4_ASAP7_75t_L g4402 ( 
.A(n_4006),
.B(n_3233),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4051),
.B(n_3086),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_4083),
.B(n_2678),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4098),
.B(n_4121),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_SL g4406 ( 
.A(n_3895),
.B(n_3925),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_SL g4407 ( 
.A(n_3895),
.B(n_3435),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4146),
.B(n_2678),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4157),
.B(n_2689),
.Y(n_4409)
);

NAND2xp33_ASAP7_75t_SL g4410 ( 
.A(n_3932),
.B(n_2934),
.Y(n_4410)
);

NAND2xp33_ASAP7_75t_SL g4411 ( 
.A(n_3928),
.B(n_2934),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_SL g4412 ( 
.A(n_3895),
.B(n_3233),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_SL g4413 ( 
.A(n_3925),
.B(n_3233),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_4159),
.B(n_2689),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_SL g4415 ( 
.A(n_3925),
.B(n_3086),
.Y(n_4415)
);

NAND2xp33_ASAP7_75t_SL g4416 ( 
.A(n_3977),
.B(n_2948),
.Y(n_4416)
);

AND2x2_ASAP7_75t_L g4417 ( 
.A(n_4052),
.B(n_3086),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_3925),
.B(n_3092),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_SL g4419 ( 
.A(n_3954),
.B(n_3092),
.Y(n_4419)
);

NAND2xp33_ASAP7_75t_SL g4420 ( 
.A(n_4014),
.B(n_4024),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_SL g4421 ( 
.A(n_3954),
.B(n_3092),
.Y(n_4421)
);

NAND2xp33_ASAP7_75t_SL g4422 ( 
.A(n_4156),
.B(n_2948),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_SL g4423 ( 
.A(n_3954),
.B(n_3119),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_SL g4424 ( 
.A(n_3954),
.B(n_3119),
.Y(n_4424)
);

NAND2xp33_ASAP7_75t_SL g4425 ( 
.A(n_4156),
.B(n_2985),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_SL g4426 ( 
.A(n_4023),
.B(n_4081),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4128),
.B(n_4129),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_3948),
.B(n_3027),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_SL g4429 ( 
.A(n_4023),
.B(n_3119),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_SL g4430 ( 
.A(n_4023),
.B(n_3324),
.Y(n_4430)
);

NAND2xp33_ASAP7_75t_SL g4431 ( 
.A(n_4156),
.B(n_2985),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_SL g4432 ( 
.A(n_4023),
.B(n_3324),
.Y(n_4432)
);

NAND2xp33_ASAP7_75t_SL g4433 ( 
.A(n_4156),
.B(n_3116),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_SL g4434 ( 
.A(n_4081),
.B(n_3324),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_SL g4435 ( 
.A(n_4081),
.B(n_3356),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_SL g4436 ( 
.A(n_4081),
.B(n_3356),
.Y(n_4436)
);

NAND2xp33_ASAP7_75t_SL g4437 ( 
.A(n_4005),
.B(n_3116),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_SL g4438 ( 
.A(n_4089),
.B(n_3356),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_SL g4439 ( 
.A(n_4089),
.B(n_3939),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_SL g4440 ( 
.A(n_4089),
.B(n_3372),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4020),
.B(n_3372),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_SL g4442 ( 
.A(n_4089),
.B(n_3372),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_SL g4443 ( 
.A(n_3939),
.B(n_3407),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_SL g4444 ( 
.A(n_4086),
.B(n_3120),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_SL g4445 ( 
.A(n_4012),
.B(n_3120),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4027),
.B(n_3272),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_SL g4447 ( 
.A(n_3979),
.B(n_3392),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4005),
.B(n_3027),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4028),
.B(n_3272),
.Y(n_4449)
);

NAND2xp33_ASAP7_75t_SL g4450 ( 
.A(n_3891),
.B(n_2718),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_SL g4451 ( 
.A(n_3979),
.B(n_4119),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_SL g4452 ( 
.A(n_4119),
.B(n_3392),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_SL g4453 ( 
.A(n_3931),
.B(n_3433),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_SL g4454 ( 
.A(n_3826),
.B(n_3433),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_SL g4455 ( 
.A(n_3826),
.B(n_3449),
.Y(n_4455)
);

OR2x2_ASAP7_75t_L g4456 ( 
.A(n_4035),
.B(n_3789),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_SL g4457 ( 
.A(n_3978),
.B(n_3449),
.Y(n_4457)
);

NAND2xp33_ASAP7_75t_SL g4458 ( 
.A(n_3880),
.B(n_2725),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4035),
.B(n_3041),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_SL g4460 ( 
.A(n_3978),
.B(n_3470),
.Y(n_4460)
);

NAND2xp33_ASAP7_75t_SL g4461 ( 
.A(n_4058),
.B(n_2728),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_SL g4462 ( 
.A(n_3952),
.B(n_3470),
.Y(n_4462)
);

NAND2xp33_ASAP7_75t_SL g4463 ( 
.A(n_4064),
.B(n_2728),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_SL g4464 ( 
.A(n_3952),
.B(n_3479),
.Y(n_4464)
);

NOR2xp33_ASAP7_75t_SL g4465 ( 
.A(n_3952),
.B(n_3041),
.Y(n_4465)
);

NAND2xp33_ASAP7_75t_SL g4466 ( 
.A(n_4148),
.B(n_2730),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_SL g4467 ( 
.A(n_3952),
.B(n_3479),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_SL g4468 ( 
.A(n_3959),
.B(n_3485),
.Y(n_4468)
);

AND2x4_ASAP7_75t_L g4469 ( 
.A(n_4036),
.B(n_3528),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_SL g4470 ( 
.A(n_3959),
.B(n_3922),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_3800),
.B(n_3041),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_SL g4472 ( 
.A(n_3795),
.B(n_3485),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_SL g4473 ( 
.A(n_3795),
.B(n_3487),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_SL g4474 ( 
.A(n_4131),
.B(n_3487),
.Y(n_4474)
);

AND2x4_ASAP7_75t_L g4475 ( 
.A(n_3916),
.B(n_3547),
.Y(n_4475)
);

AND2x4_ASAP7_75t_L g4476 ( 
.A(n_3916),
.B(n_3547),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_SL g4477 ( 
.A(n_3860),
.B(n_3501),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_SL g4478 ( 
.A(n_3860),
.B(n_3501),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_SL g4479 ( 
.A(n_3927),
.B(n_3516),
.Y(n_4479)
);

NAND2xp33_ASAP7_75t_SL g4480 ( 
.A(n_3913),
.B(n_2730),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_SL g4481 ( 
.A(n_3927),
.B(n_3516),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_SL g4482 ( 
.A(n_3953),
.B(n_3773),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_3802),
.B(n_3041),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_SL g4484 ( 
.A(n_3953),
.B(n_3773),
.Y(n_4484)
);

NAND2xp33_ASAP7_75t_SL g4485 ( 
.A(n_3913),
.B(n_2731),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_SL g4486 ( 
.A(n_3997),
.B(n_3783),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_SL g4487 ( 
.A(n_3997),
.B(n_3783),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_SL g4488 ( 
.A(n_3889),
.B(n_3548),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_3805),
.B(n_3070),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_SL g4490 ( 
.A(n_4077),
.B(n_3548),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_SL g4491 ( 
.A(n_4077),
.B(n_3590),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_SL g4492 ( 
.A(n_4085),
.B(n_4002),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_SL g4493 ( 
.A(n_4085),
.B(n_3590),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_SL g4494 ( 
.A(n_4002),
.B(n_3602),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_SL g4495 ( 
.A(n_4160),
.B(n_3602),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_SL g4496 ( 
.A(n_4160),
.B(n_3617),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_SL g4497 ( 
.A(n_3883),
.B(n_3617),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_SL g4498 ( 
.A(n_3883),
.B(n_3908),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_SL g4499 ( 
.A(n_3908),
.B(n_3625),
.Y(n_4499)
);

NAND2xp33_ASAP7_75t_SL g4500 ( 
.A(n_3905),
.B(n_2731),
.Y(n_4500)
);

NAND2xp33_ASAP7_75t_SL g4501 ( 
.A(n_3905),
.B(n_3305),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_3810),
.B(n_3070),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_SL g4503 ( 
.A(n_4143),
.B(n_3647),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_3814),
.B(n_3305),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_3833),
.B(n_3070),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_SL g4506 ( 
.A(n_3858),
.B(n_3659),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_SL g4507 ( 
.A(n_3858),
.B(n_3659),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_SL g4508 ( 
.A(n_3808),
.B(n_3665),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_SL g4509 ( 
.A(n_3808),
.B(n_3665),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_SL g4510 ( 
.A(n_3917),
.B(n_3666),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_SL g4511 ( 
.A(n_3917),
.B(n_3666),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_SL g4512 ( 
.A(n_3995),
.B(n_4039),
.Y(n_4512)
);

NAND2xp33_ASAP7_75t_SL g4513 ( 
.A(n_3966),
.B(n_754),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_SL g4514 ( 
.A(n_4045),
.B(n_3851),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_SL g4515 ( 
.A(n_3851),
.B(n_3693),
.Y(n_4515)
);

NAND2xp33_ASAP7_75t_SL g4516 ( 
.A(n_4037),
.B(n_815),
.Y(n_4516)
);

AND2x2_ASAP7_75t_L g4517 ( 
.A(n_3834),
.B(n_3554),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_SL g4518 ( 
.A(n_4017),
.B(n_3720),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_SL g4519 ( 
.A(n_4017),
.B(n_3720),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_SL g4520 ( 
.A(n_4135),
.B(n_3737),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_SL g4521 ( 
.A(n_4135),
.B(n_3737),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_SL g4522 ( 
.A(n_4115),
.B(n_3740),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_SL g4523 ( 
.A(n_4115),
.B(n_3740),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_3839),
.B(n_3070),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_3840),
.B(n_3070),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_SL g4526 ( 
.A(n_4117),
.B(n_3554),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_SL g4527 ( 
.A(n_4117),
.B(n_3558),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_SL g4528 ( 
.A(n_4106),
.B(n_3558),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_SL g4529 ( 
.A(n_4106),
.B(n_3562),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_SL g4530 ( 
.A(n_4061),
.B(n_3562),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_SL g4531 ( 
.A(n_4061),
.B(n_3991),
.Y(n_4531)
);

NAND2xp33_ASAP7_75t_SL g4532 ( 
.A(n_4037),
.B(n_822),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_SL g4533 ( 
.A(n_3991),
.B(n_3625),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_4136),
.B(n_3647),
.Y(n_4534)
);

NAND2xp5_ASAP7_75t_SL g4535 ( 
.A(n_4136),
.B(n_4151),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_SL g4536 ( 
.A(n_4151),
.B(n_3693),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_3910),
.B(n_2252),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_SL g4538 ( 
.A(n_4102),
.B(n_3741),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_3856),
.B(n_3741),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_3863),
.B(n_2252),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_SL g4541 ( 
.A(n_4102),
.B(n_3440),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_3872),
.B(n_2254),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_SL g4543 ( 
.A(n_4104),
.B(n_3745),
.Y(n_4543)
);

NAND2xp33_ASAP7_75t_SL g4544 ( 
.A(n_3888),
.B(n_822),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_SL g4545 ( 
.A(n_4104),
.B(n_2538),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_3881),
.B(n_2254),
.Y(n_4546)
);

NAND2xp5_ASAP7_75t_SL g4547 ( 
.A(n_4123),
.B(n_3980),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_3886),
.B(n_2260),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_SL g4549 ( 
.A(n_4123),
.B(n_2538),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_3890),
.B(n_2260),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_SL g4551 ( 
.A(n_3980),
.B(n_2538),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_3899),
.B(n_2264),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_SL g4553 ( 
.A(n_4118),
.B(n_2538),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_3901),
.B(n_1387),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_SL g4555 ( 
.A(n_4118),
.B(n_2538),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_SL g4556 ( 
.A(n_4065),
.B(n_2555),
.Y(n_4556)
);

NAND2xp33_ASAP7_75t_SL g4557 ( 
.A(n_3888),
.B(n_824),
.Y(n_4557)
);

NAND2xp33_ASAP7_75t_SL g4558 ( 
.A(n_3812),
.B(n_824),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_SL g4559 ( 
.A(n_4065),
.B(n_2555),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_SL g4560 ( 
.A(n_4016),
.B(n_2555),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_SL g4561 ( 
.A(n_3904),
.B(n_2555),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_SL g4562 ( 
.A(n_3906),
.B(n_2555),
.Y(n_4562)
);

O2A1O1Ixp33_ASAP7_75t_L g4563 ( 
.A1(n_4172),
.A2(n_738),
.B(n_739),
.C(n_737),
.Y(n_4563)
);

BUFx2_ASAP7_75t_L g4564 ( 
.A(n_4309),
.Y(n_4564)
);

BUFx3_ASAP7_75t_L g4565 ( 
.A(n_4386),
.Y(n_4565)
);

OAI22xp5_ASAP7_75t_SL g4566 ( 
.A1(n_4389),
.A2(n_4130),
.B1(n_4030),
.B2(n_3835),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4173),
.B(n_3919),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4264),
.B(n_4019),
.Y(n_4568)
);

A2O1A1Ixp33_ASAP7_75t_SL g4569 ( 
.A1(n_4163),
.A2(n_739),
.B(n_743),
.C(n_738),
.Y(n_4569)
);

HB1xp67_ASAP7_75t_L g4570 ( 
.A(n_4209),
.Y(n_4570)
);

HB1xp67_ASAP7_75t_L g4571 ( 
.A(n_4209),
.Y(n_4571)
);

O2A1O1Ixp33_ASAP7_75t_L g4572 ( 
.A1(n_4164),
.A2(n_749),
.B(n_756),
.C(n_743),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4543),
.A2(n_4029),
.B(n_4314),
.Y(n_4573)
);

CKINVDCx11_ASAP7_75t_R g4574 ( 
.A(n_4284),
.Y(n_4574)
);

AOI21xp5_ASAP7_75t_L g4575 ( 
.A1(n_4314),
.A2(n_4029),
.B(n_4091),
.Y(n_4575)
);

INVxp67_ASAP7_75t_L g4576 ( 
.A(n_4456),
.Y(n_4576)
);

BUFx4_ASAP7_75t_SL g4577 ( 
.A(n_4198),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4264),
.Y(n_4578)
);

INVx2_ASAP7_75t_SL g4579 ( 
.A(n_4386),
.Y(n_4579)
);

AOI222xp33_ASAP7_75t_L g4580 ( 
.A1(n_4199),
.A2(n_768),
.B1(n_757),
.B2(n_770),
.C1(n_766),
.C2(n_749),
.Y(n_4580)
);

NOR2xp33_ASAP7_75t_L g4581 ( 
.A(n_4161),
.B(n_3835),
.Y(n_4581)
);

BUFx3_ASAP7_75t_L g4582 ( 
.A(n_4386),
.Y(n_4582)
);

AND2x2_ASAP7_75t_L g4583 ( 
.A(n_4186),
.B(n_3933),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4227),
.B(n_3936),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4456),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4211),
.B(n_4240),
.Y(n_4586)
);

INVx3_ASAP7_75t_L g4587 ( 
.A(n_4284),
.Y(n_4587)
);

O2A1O1Ixp33_ASAP7_75t_SL g4588 ( 
.A1(n_4191),
.A2(n_4079),
.B(n_4091),
.C(n_4124),
.Y(n_4588)
);

CKINVDCx11_ASAP7_75t_R g4589 ( 
.A(n_4284),
.Y(n_4589)
);

O2A1O1Ixp33_ASAP7_75t_L g4590 ( 
.A1(n_4192),
.A2(n_766),
.B(n_768),
.C(n_757),
.Y(n_4590)
);

NAND2x1p5_ASAP7_75t_L g4591 ( 
.A(n_4305),
.B(n_4332),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4211),
.B(n_3942),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4210),
.B(n_3961),
.Y(n_4593)
);

BUFx2_ASAP7_75t_L g4594 ( 
.A(n_4284),
.Y(n_4594)
);

BUFx4_ASAP7_75t_SL g4595 ( 
.A(n_4198),
.Y(n_4595)
);

A2O1A1Ixp33_ASAP7_75t_L g4596 ( 
.A1(n_4437),
.A2(n_4450),
.B(n_4314),
.C(n_4544),
.Y(n_4596)
);

NAND2xp5_ASAP7_75t_SL g4597 ( 
.A(n_4289),
.B(n_4079),
.Y(n_4597)
);

INVx5_ASAP7_75t_L g4598 ( 
.A(n_4305),
.Y(n_4598)
);

AOI221xp5_ASAP7_75t_L g4599 ( 
.A1(n_4389),
.A2(n_1133),
.B1(n_1137),
.B2(n_1128),
.C(n_1123),
.Y(n_4599)
);

BUFx6f_ASAP7_75t_L g4600 ( 
.A(n_4305),
.Y(n_4600)
);

HB1xp67_ASAP7_75t_L g4601 ( 
.A(n_4341),
.Y(n_4601)
);

NAND3xp33_ASAP7_75t_L g4602 ( 
.A(n_4162),
.B(n_4097),
.C(n_839),
.Y(n_4602)
);

BUFx2_ASAP7_75t_L g4603 ( 
.A(n_4167),
.Y(n_4603)
);

AOI21xp5_ASAP7_75t_L g4604 ( 
.A1(n_4358),
.A2(n_3692),
.B(n_3930),
.Y(n_4604)
);

OR2x2_ASAP7_75t_L g4605 ( 
.A(n_4397),
.B(n_3963),
.Y(n_4605)
);

AOI22xp33_ASAP7_75t_L g4606 ( 
.A1(n_4557),
.A2(n_3788),
.B1(n_773),
.B2(n_775),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4181),
.B(n_4025),
.Y(n_4607)
);

AND2x2_ASAP7_75t_L g4608 ( 
.A(n_4271),
.B(n_3964),
.Y(n_4608)
);

O2A1O1Ixp5_ASAP7_75t_L g4609 ( 
.A1(n_4541),
.A2(n_4124),
.B(n_3923),
.C(n_3924),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4405),
.Y(n_4610)
);

OAI22xp5_ASAP7_75t_L g4611 ( 
.A1(n_4179),
.A2(n_3924),
.B1(n_3968),
.B2(n_3967),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4182),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4182),
.Y(n_4613)
);

BUFx2_ASAP7_75t_L g4614 ( 
.A(n_4236),
.Y(n_4614)
);

CKINVDCx16_ASAP7_75t_R g4615 ( 
.A(n_4174),
.Y(n_4615)
);

BUFx6f_ASAP7_75t_L g4616 ( 
.A(n_4305),
.Y(n_4616)
);

BUFx6f_ASAP7_75t_L g4617 ( 
.A(n_4332),
.Y(n_4617)
);

OAI21x1_ASAP7_75t_SL g4618 ( 
.A1(n_4292),
.A2(n_3923),
.B(n_3975),
.Y(n_4618)
);

INVx3_ASAP7_75t_L g4619 ( 
.A(n_4475),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4181),
.B(n_3996),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4405),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4197),
.Y(n_4622)
);

AOI22xp5_ASAP7_75t_L g4623 ( 
.A1(n_4480),
.A2(n_3848),
.B1(n_3798),
.B2(n_3842),
.Y(n_4623)
);

HB1xp67_ASAP7_75t_L g4624 ( 
.A(n_4320),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_SL g4625 ( 
.A(n_4196),
.B(n_4018),
.Y(n_4625)
);

AOI21xp5_ASAP7_75t_L g4626 ( 
.A1(n_4362),
.A2(n_4120),
.B(n_3930),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4197),
.Y(n_4627)
);

CKINVDCx5p33_ASAP7_75t_R g4628 ( 
.A(n_4420),
.Y(n_4628)
);

AND2x2_ASAP7_75t_L g4629 ( 
.A(n_4271),
.B(n_3981),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4517),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4183),
.B(n_4001),
.Y(n_4631)
);

INVx3_ASAP7_75t_L g4632 ( 
.A(n_4475),
.Y(n_4632)
);

BUFx10_ASAP7_75t_L g4633 ( 
.A(n_4332),
.Y(n_4633)
);

INVx4_ASAP7_75t_L g4634 ( 
.A(n_4332),
.Y(n_4634)
);

BUFx3_ASAP7_75t_L g4635 ( 
.A(n_4386),
.Y(n_4635)
);

AOI211xp5_ASAP7_75t_L g4636 ( 
.A1(n_4282),
.A2(n_773),
.B(n_775),
.C(n_770),
.Y(n_4636)
);

BUFx3_ASAP7_75t_L g4637 ( 
.A(n_4402),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4446),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4517),
.Y(n_4639)
);

BUFx6f_ASAP7_75t_L g4640 ( 
.A(n_4354),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4539),
.Y(n_4641)
);

BUFx6f_ASAP7_75t_L g4642 ( 
.A(n_4354),
.Y(n_4642)
);

AND2x6_ASAP7_75t_L g4643 ( 
.A(n_4207),
.B(n_3848),
.Y(n_4643)
);

OAI22xp5_ASAP7_75t_L g4644 ( 
.A1(n_4537),
.A2(n_3985),
.B1(n_3987),
.B2(n_3984),
.Y(n_4644)
);

BUFx8_ASAP7_75t_SL g4645 ( 
.A(n_4245),
.Y(n_4645)
);

INVx5_ASAP7_75t_L g4646 ( 
.A(n_4354),
.Y(n_4646)
);

NAND2x1p5_ASAP7_75t_L g4647 ( 
.A(n_4354),
.B(n_3929),
.Y(n_4647)
);

NAND2x1_ASAP7_75t_L g4648 ( 
.A(n_4475),
.B(n_3848),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4539),
.Y(n_4649)
);

O2A1O1Ixp33_ASAP7_75t_L g4650 ( 
.A1(n_4194),
.A2(n_792),
.B(n_800),
.C(n_786),
.Y(n_4650)
);

HB1xp67_ASAP7_75t_L g4651 ( 
.A(n_4320),
.Y(n_4651)
);

AOI21xp5_ASAP7_75t_L g4652 ( 
.A1(n_4359),
.A2(n_4120),
.B(n_4018),
.Y(n_4652)
);

BUFx6f_ASAP7_75t_L g4653 ( 
.A(n_4402),
.Y(n_4653)
);

BUFx2_ASAP7_75t_L g4654 ( 
.A(n_4401),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4427),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_4446),
.Y(n_4656)
);

AOI22xp5_ASAP7_75t_L g4657 ( 
.A1(n_4485),
.A2(n_3848),
.B1(n_3798),
.B2(n_3842),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4441),
.B(n_4040),
.Y(n_4658)
);

INVx2_ASAP7_75t_L g4659 ( 
.A(n_4449),
.Y(n_4659)
);

NOR3xp33_ASAP7_75t_L g4660 ( 
.A(n_4516),
.B(n_792),
.C(n_786),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4441),
.B(n_3798),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4427),
.Y(n_4662)
);

INVx4_ASAP7_75t_L g4663 ( 
.A(n_4293),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4183),
.B(n_3848),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4368),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4201),
.B(n_3876),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4368),
.Y(n_4667)
);

INVx4_ASAP7_75t_L g4668 ( 
.A(n_4293),
.Y(n_4668)
);

A2O1A1Ixp33_ASAP7_75t_L g4669 ( 
.A1(n_4466),
.A2(n_1171),
.B(n_1193),
.C(n_1152),
.Y(n_4669)
);

BUFx6f_ASAP7_75t_L g4670 ( 
.A(n_4402),
.Y(n_4670)
);

HB1xp67_ASAP7_75t_L g4671 ( 
.A(n_4397),
.Y(n_4671)
);

OAI22xp5_ASAP7_75t_L g4672 ( 
.A1(n_4189),
.A2(n_3960),
.B1(n_3958),
.B2(n_3885),
.Y(n_4672)
);

NAND2x1p5_ASAP7_75t_L g4673 ( 
.A(n_4207),
.B(n_3929),
.Y(n_4673)
);

BUFx2_ASAP7_75t_SL g4674 ( 
.A(n_4203),
.Y(n_4674)
);

AOI22xp33_ASAP7_75t_L g4675 ( 
.A1(n_4188),
.A2(n_802),
.B1(n_806),
.B2(n_800),
.Y(n_4675)
);

AND2x4_ASAP7_75t_L g4676 ( 
.A(n_4469),
.B(n_3842),
.Y(n_4676)
);

AOI22xp33_ASAP7_75t_L g4677 ( 
.A1(n_4188),
.A2(n_4470),
.B1(n_4500),
.B2(n_4501),
.Y(n_4677)
);

NAND2x1p5_ASAP7_75t_L g4678 ( 
.A(n_4207),
.B(n_3983),
.Y(n_4678)
);

OAI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4175),
.A2(n_3958),
.B1(n_3960),
.B2(n_3885),
.Y(n_4679)
);

BUFx2_ASAP7_75t_L g4680 ( 
.A(n_4371),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4312),
.Y(n_4681)
);

INVx1_ASAP7_75t_SL g4682 ( 
.A(n_4178),
.Y(n_4682)
);

A2O1A1Ixp33_ASAP7_75t_SL g4683 ( 
.A1(n_4344),
.A2(n_806),
.B(n_830),
.C(n_802),
.Y(n_4683)
);

HB1xp67_ASAP7_75t_L g4684 ( 
.A(n_4170),
.Y(n_4684)
);

AOI21xp5_ASAP7_75t_L g4685 ( 
.A1(n_4291),
.A2(n_4033),
.B(n_4015),
.Y(n_4685)
);

HB1xp67_ASAP7_75t_L g4686 ( 
.A(n_4535),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4554),
.Y(n_4687)
);

AOI22xp33_ASAP7_75t_L g4688 ( 
.A1(n_4547),
.A2(n_830),
.B1(n_837),
.B2(n_834),
.Y(n_4688)
);

A2O1A1Ixp33_ASAP7_75t_L g4689 ( 
.A1(n_4513),
.A2(n_1211),
.B(n_1212),
.C(n_1206),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4185),
.B(n_3876),
.Y(n_4690)
);

O2A1O1Ixp33_ASAP7_75t_L g4691 ( 
.A1(n_4495),
.A2(n_837),
.B(n_838),
.C(n_834),
.Y(n_4691)
);

HB1xp67_ASAP7_75t_L g4692 ( 
.A(n_4549),
.Y(n_4692)
);

AND2x2_ASAP7_75t_L g4693 ( 
.A(n_4168),
.B(n_3885),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4449),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4250),
.B(n_3877),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4218),
.B(n_3877),
.Y(n_4696)
);

INVx3_ASAP7_75t_L g4697 ( 
.A(n_4475),
.Y(n_4697)
);

A2O1A1Ixp33_ASAP7_75t_SL g4698 ( 
.A1(n_4175),
.A2(n_839),
.B(n_843),
.C(n_838),
.Y(n_4698)
);

OAI22xp5_ASAP7_75t_L g4699 ( 
.A1(n_4176),
.A2(n_3960),
.B1(n_3958),
.B2(n_3345),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4554),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4319),
.Y(n_4701)
);

INVx2_ASAP7_75t_L g4702 ( 
.A(n_4504),
.Y(n_4702)
);

O2A1O1Ixp33_ASAP7_75t_L g4703 ( 
.A1(n_4496),
.A2(n_847),
.B(n_869),
.C(n_843),
.Y(n_4703)
);

OAI22xp5_ASAP7_75t_L g4704 ( 
.A1(n_4176),
.A2(n_3345),
.B1(n_3337),
.B2(n_869),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_SL g4705 ( 
.A(n_4202),
.B(n_4206),
.Y(n_4705)
);

INVx2_ASAP7_75t_L g4706 ( 
.A(n_4504),
.Y(n_4706)
);

NOR2xp33_ASAP7_75t_L g4707 ( 
.A(n_4180),
.B(n_847),
.Y(n_4707)
);

BUFx6f_ASAP7_75t_L g4708 ( 
.A(n_4402),
.Y(n_4708)
);

HB1xp67_ASAP7_75t_L g4709 ( 
.A(n_4403),
.Y(n_4709)
);

INVx4_ASAP7_75t_L g4710 ( 
.A(n_4293),
.Y(n_4710)
);

BUFx2_ASAP7_75t_L g4711 ( 
.A(n_4378),
.Y(n_4711)
);

INVx2_ASAP7_75t_L g4712 ( 
.A(n_4403),
.Y(n_4712)
);

NOR2xp33_ASAP7_75t_L g4713 ( 
.A(n_4447),
.B(n_871),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4342),
.Y(n_4714)
);

INVxp67_ASAP7_75t_SL g4715 ( 
.A(n_4538),
.Y(n_4715)
);

BUFx2_ASAP7_75t_L g4716 ( 
.A(n_4290),
.Y(n_4716)
);

INVxp67_ASAP7_75t_L g4717 ( 
.A(n_4345),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_SL g4718 ( 
.A(n_4458),
.B(n_4033),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4417),
.Y(n_4719)
);

AOI21xp5_ASAP7_75t_L g4720 ( 
.A1(n_4307),
.A2(n_4015),
.B(n_3983),
.Y(n_4720)
);

OAI22xp5_ASAP7_75t_L g4721 ( 
.A1(n_4468),
.A2(n_3345),
.B1(n_3337),
.B2(n_876),
.Y(n_4721)
);

OAI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_4190),
.A2(n_3345),
.B1(n_3337),
.B2(n_876),
.Y(n_4722)
);

OR2x6_ASAP7_75t_SL g4723 ( 
.A(n_4350),
.B(n_3792),
.Y(n_4723)
);

INVx4_ASAP7_75t_SL g4724 ( 
.A(n_4207),
.Y(n_4724)
);

AO32x1_ASAP7_75t_L g4725 ( 
.A1(n_4417),
.A2(n_3878),
.A3(n_3790),
.B1(n_3791),
.B2(n_3787),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_4404),
.Y(n_4726)
);

BUFx2_ASAP7_75t_L g4727 ( 
.A(n_4411),
.Y(n_4727)
);

AOI22xp5_ASAP7_75t_L g4728 ( 
.A1(n_4313),
.A2(n_4010),
.B1(n_3792),
.B2(n_3149),
.Y(n_4728)
);

INVx2_ASAP7_75t_SL g4729 ( 
.A(n_4212),
.Y(n_4729)
);

BUFx2_ASAP7_75t_L g4730 ( 
.A(n_4416),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4215),
.B(n_3878),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4215),
.B(n_3784),
.Y(n_4732)
);

BUFx12f_ASAP7_75t_L g4733 ( 
.A(n_4293),
.Y(n_4733)
);

CKINVDCx5p33_ASAP7_75t_R g4734 ( 
.A(n_4558),
.Y(n_4734)
);

AOI22xp33_ASAP7_75t_L g4735 ( 
.A1(n_4168),
.A2(n_878),
.B1(n_886),
.B2(n_871),
.Y(n_4735)
);

BUFx8_ASAP7_75t_SL g4736 ( 
.A(n_4469),
.Y(n_4736)
);

CKINVDCx8_ASAP7_75t_R g4737 ( 
.A(n_4469),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_SL g4738 ( 
.A(n_4283),
.B(n_2574),
.Y(n_4738)
);

HB1xp67_ASAP7_75t_L g4739 ( 
.A(n_4471),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_SL g4740 ( 
.A(n_4387),
.B(n_2574),
.Y(n_4740)
);

NOR2xp33_ASAP7_75t_L g4741 ( 
.A(n_4187),
.B(n_878),
.Y(n_4741)
);

HB1xp67_ASAP7_75t_L g4742 ( 
.A(n_4471),
.Y(n_4742)
);

OAI22xp5_ASAP7_75t_L g4743 ( 
.A1(n_4200),
.A2(n_3337),
.B1(n_905),
.B2(n_906),
.Y(n_4743)
);

BUFx2_ASAP7_75t_L g4744 ( 
.A(n_4476),
.Y(n_4744)
);

AND2x4_ASAP7_75t_SL g4745 ( 
.A(n_4469),
.B(n_3998),
.Y(n_4745)
);

BUFx3_ASAP7_75t_L g4746 ( 
.A(n_4294),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4483),
.Y(n_4747)
);

CKINVDCx8_ASAP7_75t_R g4748 ( 
.A(n_4294),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_SL g4749 ( 
.A(n_4461),
.B(n_2574),
.Y(n_4749)
);

AOI222xp33_ASAP7_75t_SL g4750 ( 
.A1(n_4512),
.A2(n_914),
.B1(n_905),
.B2(n_921),
.C1(n_906),
.C2(n_886),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4404),
.Y(n_4751)
);

OR2x2_ASAP7_75t_L g4752 ( 
.A(n_4451),
.B(n_3809),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4483),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4489),
.Y(n_4754)
);

INVx2_ASAP7_75t_L g4755 ( 
.A(n_4408),
.Y(n_4755)
);

AOI21xp5_ASAP7_75t_L g4756 ( 
.A1(n_4465),
.A2(n_4041),
.B(n_3167),
.Y(n_4756)
);

INVx3_ASAP7_75t_L g4757 ( 
.A(n_4476),
.Y(n_4757)
);

OAI22xp5_ASAP7_75t_L g4758 ( 
.A1(n_4321),
.A2(n_921),
.B1(n_928),
.B2(n_914),
.Y(n_4758)
);

A2O1A1Ixp33_ASAP7_75t_L g4759 ( 
.A1(n_4532),
.A2(n_1226),
.B(n_1230),
.C(n_1215),
.Y(n_4759)
);

BUFx12f_ASAP7_75t_L g4760 ( 
.A(n_4294),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4408),
.Y(n_4761)
);

INVx3_ASAP7_75t_L g4762 ( 
.A(n_4476),
.Y(n_4762)
);

BUFx3_ASAP7_75t_L g4763 ( 
.A(n_4294),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_SL g4764 ( 
.A(n_4463),
.B(n_2574),
.Y(n_4764)
);

O2A1O1Ixp33_ASAP7_75t_L g4765 ( 
.A1(n_4343),
.A2(n_928),
.B(n_933),
.C(n_931),
.Y(n_4765)
);

CKINVDCx5p33_ASAP7_75t_R g4766 ( 
.A(n_4214),
.Y(n_4766)
);

BUFx6f_ASAP7_75t_L g4767 ( 
.A(n_4221),
.Y(n_4767)
);

BUFx2_ASAP7_75t_L g4768 ( 
.A(n_4476),
.Y(n_4768)
);

NOR2x1_ASAP7_75t_L g4769 ( 
.A(n_4184),
.B(n_1387),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4489),
.Y(n_4770)
);

AOI22xp33_ASAP7_75t_L g4771 ( 
.A1(n_4551),
.A2(n_931),
.B1(n_941),
.B2(n_933),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4502),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4502),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_4409),
.Y(n_4774)
);

INVx2_ASAP7_75t_L g4775 ( 
.A(n_4409),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4505),
.Y(n_4776)
);

AOI21xp5_ASAP7_75t_L g4777 ( 
.A1(n_4465),
.A2(n_4259),
.B(n_4443),
.Y(n_4777)
);

BUFx12f_ASAP7_75t_L g4778 ( 
.A(n_4221),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4505),
.Y(n_4779)
);

AOI22xp5_ASAP7_75t_L g4780 ( 
.A1(n_4253),
.A2(n_4010),
.B1(n_3149),
.B2(n_3175),
.Y(n_4780)
);

CKINVDCx20_ASAP7_75t_R g4781 ( 
.A(n_4256),
.Y(n_4781)
);

O2A1O1Ixp33_ASAP7_75t_L g4782 ( 
.A1(n_4177),
.A2(n_4193),
.B(n_4205),
.C(n_4477),
.Y(n_4782)
);

OAI22xp33_ASAP7_75t_L g4783 ( 
.A1(n_4195),
.A2(n_942),
.B1(n_961),
.B2(n_948),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4414),
.Y(n_4784)
);

A2O1A1Ixp33_ASAP7_75t_L g4785 ( 
.A1(n_4472),
.A2(n_1240),
.B(n_942),
.C(n_948),
.Y(n_4785)
);

INVx3_ASAP7_75t_L g4786 ( 
.A(n_4221),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4524),
.Y(n_4787)
);

INVxp67_ASAP7_75t_L g4788 ( 
.A(n_4533),
.Y(n_4788)
);

AOI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4553),
.A2(n_4041),
.B(n_3167),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_4414),
.Y(n_4790)
);

AO21x1_ASAP7_75t_L g4791 ( 
.A1(n_4385),
.A2(n_957),
.B(n_941),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_SL g4792 ( 
.A(n_4384),
.B(n_2574),
.Y(n_4792)
);

INVx2_ASAP7_75t_SL g4793 ( 
.A(n_4503),
.Y(n_4793)
);

AND2x4_ASAP7_75t_L g4794 ( 
.A(n_4221),
.B(n_3819),
.Y(n_4794)
);

NOR2xp33_ASAP7_75t_L g4795 ( 
.A(n_4171),
.B(n_957),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4257),
.B(n_3822),
.Y(n_4796)
);

INVx2_ASAP7_75t_L g4797 ( 
.A(n_4352),
.Y(n_4797)
);

CKINVDCx5p33_ASAP7_75t_R g4798 ( 
.A(n_4258),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4352),
.Y(n_4799)
);

INVxp67_ASAP7_75t_SL g4800 ( 
.A(n_4265),
.Y(n_4800)
);

AND2x4_ASAP7_75t_L g4801 ( 
.A(n_4241),
.B(n_3841),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4524),
.Y(n_4802)
);

A2O1A1Ixp33_ASAP7_75t_L g4803 ( 
.A1(n_4473),
.A2(n_4233),
.B(n_4219),
.C(n_4531),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4525),
.Y(n_4804)
);

OAI22xp5_ASAP7_75t_L g4805 ( 
.A1(n_4448),
.A2(n_4514),
.B1(n_4365),
.B2(n_4369),
.Y(n_4805)
);

HB1xp67_ASAP7_75t_L g4806 ( 
.A(n_4525),
.Y(n_4806)
);

HB1xp67_ASAP7_75t_L g4807 ( 
.A(n_4224),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4353),
.Y(n_4808)
);

AND2x4_ASAP7_75t_L g4809 ( 
.A(n_4241),
.B(n_3853),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_L g4810 ( 
.A(n_4195),
.B(n_3855),
.Y(n_4810)
);

INVx3_ASAP7_75t_L g4811 ( 
.A(n_4241),
.Y(n_4811)
);

A2O1A1Ixp33_ASAP7_75t_L g4812 ( 
.A1(n_4454),
.A2(n_962),
.B(n_971),
.C(n_961),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4169),
.Y(n_4813)
);

OAI22x1_ASAP7_75t_L g4814 ( 
.A1(n_4220),
.A2(n_971),
.B1(n_973),
.B2(n_962),
.Y(n_4814)
);

OAI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4448),
.A2(n_977),
.B1(n_986),
.B2(n_973),
.Y(n_4815)
);

A2O1A1Ixp33_ASAP7_75t_L g4816 ( 
.A1(n_4455),
.A2(n_4041),
.B(n_986),
.C(n_988),
.Y(n_4816)
);

A2O1A1Ixp33_ASAP7_75t_L g4817 ( 
.A1(n_4508),
.A2(n_988),
.B(n_989),
.C(n_977),
.Y(n_4817)
);

INVx2_ASAP7_75t_L g4818 ( 
.A(n_4353),
.Y(n_4818)
);

NOR2xp33_ASAP7_75t_L g4819 ( 
.A(n_4204),
.B(n_989),
.Y(n_4819)
);

INVx3_ASAP7_75t_L g4820 ( 
.A(n_4241),
.Y(n_4820)
);

AND2x2_ASAP7_75t_L g4821 ( 
.A(n_4363),
.B(n_994),
.Y(n_4821)
);

AND2x4_ASAP7_75t_L g4822 ( 
.A(n_4230),
.B(n_3857),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4366),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4366),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4377),
.Y(n_4825)
);

INVx2_ASAP7_75t_SL g4826 ( 
.A(n_4498),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4380),
.B(n_3859),
.Y(n_4827)
);

INVx2_ASAP7_75t_L g4828 ( 
.A(n_4377),
.Y(n_4828)
);

INVx3_ASAP7_75t_L g4829 ( 
.A(n_4459),
.Y(n_4829)
);

OAI22xp33_ASAP7_75t_L g4830 ( 
.A1(n_4540),
.A2(n_999),
.B1(n_1001),
.B2(n_994),
.Y(n_4830)
);

OAI21xp33_ASAP7_75t_L g4831 ( 
.A1(n_4166),
.A2(n_831),
.B(n_827),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4542),
.Y(n_4832)
);

A2O1A1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4509),
.A2(n_4280),
.B(n_4281),
.C(n_4494),
.Y(n_4833)
);

A2O1A1Ixp33_ASAP7_75t_L g4834 ( 
.A1(n_4267),
.A2(n_1001),
.B(n_1002),
.C(n_999),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4546),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4367),
.A2(n_1014),
.B1(n_1016),
.B2(n_1002),
.Y(n_4836)
);

AOI22xp33_ASAP7_75t_L g4837 ( 
.A1(n_4165),
.A2(n_1014),
.B1(n_1017),
.B2(n_1016),
.Y(n_4837)
);

INVx2_ASAP7_75t_L g4838 ( 
.A(n_4548),
.Y(n_4838)
);

BUFx3_ASAP7_75t_L g4839 ( 
.A(n_4550),
.Y(n_4839)
);

INVx2_ASAP7_75t_L g4840 ( 
.A(n_4552),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4246),
.B(n_4247),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4273),
.Y(n_4842)
);

NOR2xp33_ASAP7_75t_SL g4843 ( 
.A(n_4428),
.B(n_3861),
.Y(n_4843)
);

NAND2x1p5_ASAP7_75t_L g4844 ( 
.A(n_4462),
.B(n_3864),
.Y(n_4844)
);

INVx4_ASAP7_75t_L g4845 ( 
.A(n_4216),
.Y(n_4845)
);

OAI22xp5_ASAP7_75t_L g4846 ( 
.A1(n_4370),
.A2(n_1019),
.B1(n_1022),
.B2(n_1017),
.Y(n_4846)
);

INVx2_ASAP7_75t_L g4847 ( 
.A(n_4248),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4286),
.Y(n_4848)
);

INVx2_ASAP7_75t_L g4849 ( 
.A(n_4288),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4225),
.Y(n_4850)
);

BUFx6f_ASAP7_75t_L g4851 ( 
.A(n_4326),
.Y(n_4851)
);

CKINVDCx14_ASAP7_75t_R g4852 ( 
.A(n_4217),
.Y(n_4852)
);

O2A1O1Ixp33_ASAP7_75t_L g4853 ( 
.A1(n_4478),
.A2(n_1019),
.B(n_1026),
.C(n_1022),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4322),
.B(n_3865),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4226),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4228),
.B(n_3867),
.Y(n_4856)
);

NOR2xp33_ASAP7_75t_L g4857 ( 
.A(n_4266),
.B(n_1026),
.Y(n_4857)
);

INVx2_ASAP7_75t_L g4858 ( 
.A(n_4249),
.Y(n_4858)
);

INVx2_ASAP7_75t_SL g4859 ( 
.A(n_4346),
.Y(n_4859)
);

INVx4_ASAP7_75t_L g4860 ( 
.A(n_4208),
.Y(n_4860)
);

AOI21xp5_ASAP7_75t_L g4861 ( 
.A1(n_4555),
.A2(n_3167),
.B(n_3132),
.Y(n_4861)
);

BUFx4f_ASAP7_75t_L g4862 ( 
.A(n_4410),
.Y(n_4862)
);

BUFx6f_ASAP7_75t_L g4863 ( 
.A(n_4335),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4522),
.Y(n_4864)
);

BUFx6f_ASAP7_75t_L g4865 ( 
.A(n_4373),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_SL g4866 ( 
.A(n_4382),
.B(n_2576),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4364),
.B(n_3870),
.Y(n_4867)
);

HB1xp67_ASAP7_75t_L g4868 ( 
.A(n_4269),
.Y(n_4868)
);

INVx2_ASAP7_75t_L g4869 ( 
.A(n_4251),
.Y(n_4869)
);

INVx3_ASAP7_75t_L g4870 ( 
.A(n_4459),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4523),
.Y(n_4871)
);

A2O1A1Ixp33_ASAP7_75t_L g4872 ( 
.A1(n_4453),
.A2(n_1037),
.B(n_1050),
.C(n_1028),
.Y(n_4872)
);

BUFx3_ASAP7_75t_L g4873 ( 
.A(n_4428),
.Y(n_4873)
);

O2A1O1Ixp5_ASAP7_75t_L g4874 ( 
.A1(n_4300),
.A2(n_2789),
.B(n_2791),
.C(n_2788),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4526),
.Y(n_4875)
);

BUFx12f_ASAP7_75t_L g4876 ( 
.A(n_4347),
.Y(n_4876)
);

NAND2xp33_ASAP7_75t_L g4877 ( 
.A(n_4213),
.B(n_3350),
.Y(n_4877)
);

HB1xp67_ASAP7_75t_L g4878 ( 
.A(n_4242),
.Y(n_4878)
);

INVxp67_ASAP7_75t_SL g4879 ( 
.A(n_4301),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_4234),
.B(n_4492),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4527),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4351),
.B(n_3871),
.Y(n_4882)
);

O2A1O1Ixp33_ASAP7_75t_L g4883 ( 
.A1(n_4488),
.A2(n_1028),
.B(n_1050),
.C(n_1037),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4252),
.Y(n_4884)
);

INVxp67_ASAP7_75t_L g4885 ( 
.A(n_4510),
.Y(n_4885)
);

AOI22xp5_ASAP7_75t_L g4886 ( 
.A1(n_4235),
.A2(n_3073),
.B1(n_3175),
.B2(n_3149),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_SL g4887 ( 
.A(n_4439),
.B(n_2576),
.Y(n_4887)
);

INVx4_ASAP7_75t_L g4888 ( 
.A(n_4406),
.Y(n_4888)
);

NAND2x1p5_ASAP7_75t_L g4889 ( 
.A(n_4464),
.B(n_3874),
.Y(n_4889)
);

O2A1O1Ixp33_ASAP7_75t_L g4890 ( 
.A1(n_4270),
.A2(n_1063),
.B(n_1069),
.C(n_1064),
.Y(n_4890)
);

INVx1_ASAP7_75t_L g4891 ( 
.A(n_4243),
.Y(n_4891)
);

BUFx12f_ASAP7_75t_L g4892 ( 
.A(n_4348),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4254),
.A2(n_3227),
.B(n_3132),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4244),
.Y(n_4894)
);

AOI21x1_ASAP7_75t_L g4895 ( 
.A1(n_4407),
.A2(n_1390),
.B(n_1388),
.Y(n_4895)
);

INVx6_ASAP7_75t_SL g4896 ( 
.A(n_4339),
.Y(n_4896)
);

CKINVDCx6p67_ASAP7_75t_R g4897 ( 
.A(n_4528),
.Y(n_4897)
);

BUFx2_ASAP7_75t_L g4898 ( 
.A(n_4422),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4268),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_SL g4900 ( 
.A(n_4272),
.B(n_2576),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_SL g4901 ( 
.A(n_4511),
.B(n_2576),
.Y(n_4901)
);

INVx2_ASAP7_75t_L g4902 ( 
.A(n_4302),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4287),
.Y(n_4903)
);

HB1xp67_ASAP7_75t_L g4904 ( 
.A(n_4285),
.Y(n_4904)
);

BUFx6f_ASAP7_75t_L g4905 ( 
.A(n_4374),
.Y(n_4905)
);

INVx5_ASAP7_75t_L g4906 ( 
.A(n_4425),
.Y(n_4906)
);

AOI21xp5_ASAP7_75t_L g4907 ( 
.A1(n_4545),
.A2(n_3227),
.B(n_3132),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4562),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4355),
.B(n_3875),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4444),
.B(n_3893),
.Y(n_4910)
);

BUFx3_ASAP7_75t_L g4911 ( 
.A(n_4340),
.Y(n_4911)
);

BUFx6f_ASAP7_75t_L g4912 ( 
.A(n_4323),
.Y(n_4912)
);

AOI222xp33_ASAP7_75t_L g4913 ( 
.A1(n_4520),
.A2(n_1069),
.B1(n_1063),
.B2(n_1075),
.C1(n_1072),
.C2(n_1064),
.Y(n_4913)
);

BUFx2_ASAP7_75t_L g4914 ( 
.A(n_4431),
.Y(n_4914)
);

NAND2xp5_ASAP7_75t_L g4915 ( 
.A(n_4255),
.B(n_3937),
.Y(n_4915)
);

INVx4_ASAP7_75t_L g4916 ( 
.A(n_4426),
.Y(n_4916)
);

INVx3_ASAP7_75t_L g4917 ( 
.A(n_4433),
.Y(n_4917)
);

INVxp67_ASAP7_75t_L g4918 ( 
.A(n_4231),
.Y(n_4918)
);

INVx2_ASAP7_75t_L g4919 ( 
.A(n_4561),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4260),
.B(n_3944),
.Y(n_4920)
);

NOR2xp33_ASAP7_75t_L g4921 ( 
.A(n_4529),
.B(n_1072),
.Y(n_4921)
);

O2A1O1Ixp33_ASAP7_75t_L g4922 ( 
.A1(n_4474),
.A2(n_1075),
.B(n_1078),
.C(n_1076),
.Y(n_4922)
);

AOI22xp33_ASAP7_75t_L g4923 ( 
.A1(n_4521),
.A2(n_1076),
.B1(n_1085),
.B2(n_1078),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_SL g4924 ( 
.A(n_4222),
.B(n_2576),
.Y(n_4924)
);

BUFx3_ASAP7_75t_L g4925 ( 
.A(n_4239),
.Y(n_4925)
);

OAI22x1_ASAP7_75t_L g4926 ( 
.A1(n_4279),
.A2(n_1090),
.B1(n_1095),
.B2(n_1085),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4295),
.Y(n_4927)
);

BUFx2_ASAP7_75t_SL g4928 ( 
.A(n_4560),
.Y(n_4928)
);

O2A1O1Ixp33_ASAP7_75t_L g4929 ( 
.A1(n_4356),
.A2(n_1090),
.B(n_1107),
.C(n_1095),
.Y(n_4929)
);

INVx3_ASAP7_75t_L g4930 ( 
.A(n_4303),
.Y(n_4930)
);

O2A1O1Ixp5_ASAP7_75t_L g4931 ( 
.A1(n_4232),
.A2(n_2791),
.B(n_2792),
.C(n_2789),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4530),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4534),
.Y(n_4933)
);

BUFx6f_ASAP7_75t_L g4934 ( 
.A(n_4324),
.Y(n_4934)
);

OR2x2_ASAP7_75t_L g4935 ( 
.A(n_4223),
.B(n_3951),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4536),
.Y(n_4936)
);

BUFx4f_ASAP7_75t_L g4937 ( 
.A(n_4556),
.Y(n_4937)
);

INVx2_ASAP7_75t_L g4938 ( 
.A(n_4237),
.Y(n_4938)
);

O2A1O1Ixp33_ASAP7_75t_L g4939 ( 
.A1(n_4357),
.A2(n_1107),
.B(n_1116),
.C(n_1108),
.Y(n_4939)
);

BUFx6f_ASAP7_75t_L g4940 ( 
.A(n_4325),
.Y(n_4940)
);

BUFx6f_ASAP7_75t_L g4941 ( 
.A(n_4327),
.Y(n_4941)
);

BUFx6f_ASAP7_75t_L g4942 ( 
.A(n_4328),
.Y(n_4942)
);

INVx1_ASAP7_75t_SL g4943 ( 
.A(n_4497),
.Y(n_4943)
);

BUFx2_ASAP7_75t_L g4944 ( 
.A(n_4388),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_SL g4945 ( 
.A(n_4445),
.B(n_4261),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4238),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4229),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4452),
.Y(n_4948)
);

AOI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_4329),
.A2(n_3227),
.B(n_2778),
.Y(n_4949)
);

INVx4_ASAP7_75t_L g4950 ( 
.A(n_4304),
.Y(n_4950)
);

INVx2_ASAP7_75t_SL g4951 ( 
.A(n_4306),
.Y(n_4951)
);

CKINVDCx20_ASAP7_75t_R g4952 ( 
.A(n_4499),
.Y(n_4952)
);

AOI21xp5_ASAP7_75t_L g4953 ( 
.A1(n_4330),
.A2(n_4333),
.B(n_4331),
.Y(n_4953)
);

INVxp67_ASAP7_75t_L g4954 ( 
.A(n_4262),
.Y(n_4954)
);

INVx4_ASAP7_75t_L g4955 ( 
.A(n_4308),
.Y(n_4955)
);

BUFx6f_ASAP7_75t_L g4956 ( 
.A(n_4334),
.Y(n_4956)
);

O2A1O1Ixp33_ASAP7_75t_L g4957 ( 
.A1(n_4263),
.A2(n_1108),
.B(n_1117),
.C(n_1116),
.Y(n_4957)
);

A2O1A1Ixp33_ASAP7_75t_L g4958 ( 
.A1(n_4393),
.A2(n_1124),
.B(n_1125),
.C(n_1117),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4349),
.Y(n_4959)
);

INVx2_ASAP7_75t_L g4960 ( 
.A(n_4482),
.Y(n_4960)
);

A2O1A1Ixp33_ASAP7_75t_L g4961 ( 
.A1(n_4398),
.A2(n_1125),
.B(n_1131),
.C(n_1124),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4360),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_SL g4963 ( 
.A(n_4518),
.B(n_4519),
.Y(n_4963)
);

BUFx8_ASAP7_75t_SL g4964 ( 
.A(n_4310),
.Y(n_4964)
);

AOI221xp5_ASAP7_75t_L g4965 ( 
.A1(n_4274),
.A2(n_1136),
.B1(n_1139),
.B2(n_1132),
.C(n_1131),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_SL g4966 ( 
.A(n_4457),
.B(n_2581),
.Y(n_4966)
);

BUFx3_ASAP7_75t_L g4967 ( 
.A(n_4311),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_SL g4968 ( 
.A(n_4460),
.B(n_2581),
.Y(n_4968)
);

INVx3_ASAP7_75t_L g4969 ( 
.A(n_4484),
.Y(n_4969)
);

AOI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4336),
.A2(n_2778),
.B(n_2775),
.Y(n_4970)
);

BUFx6f_ASAP7_75t_L g4971 ( 
.A(n_4337),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_L g4972 ( 
.A(n_4375),
.B(n_4376),
.Y(n_4972)
);

AOI21xp5_ASAP7_75t_L g4973 ( 
.A1(n_4372),
.A2(n_2872),
.B(n_2861),
.Y(n_4973)
);

AND2x4_ASAP7_75t_L g4974 ( 
.A(n_4315),
.B(n_3956),
.Y(n_4974)
);

AOI22xp5_ASAP7_75t_L g4975 ( 
.A1(n_4506),
.A2(n_3073),
.B1(n_3175),
.B2(n_3149),
.Y(n_4975)
);

INVx4_ASAP7_75t_L g4976 ( 
.A(n_4479),
.Y(n_4976)
);

BUFx6f_ASAP7_75t_L g4977 ( 
.A(n_4559),
.Y(n_4977)
);

NOR2xp33_ASAP7_75t_SL g4978 ( 
.A(n_4379),
.B(n_3969),
.Y(n_4978)
);

INVx2_ASAP7_75t_L g4979 ( 
.A(n_4486),
.Y(n_4979)
);

AND2x2_ASAP7_75t_L g4980 ( 
.A(n_4316),
.B(n_4317),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4487),
.Y(n_4981)
);

INVx3_ASAP7_75t_L g4982 ( 
.A(n_4587),
.Y(n_4982)
);

AOI21xp5_ASAP7_75t_L g4983 ( 
.A1(n_4877),
.A2(n_4491),
.B(n_4490),
.Y(n_4983)
);

AO31x2_ASAP7_75t_L g4984 ( 
.A1(n_4815),
.A2(n_3990),
.A3(n_3999),
.B(n_3982),
.Y(n_4984)
);

AOI21xp5_ASAP7_75t_L g4985 ( 
.A1(n_4705),
.A2(n_4596),
.B(n_4740),
.Y(n_4985)
);

AO31x2_ASAP7_75t_L g4986 ( 
.A1(n_4611),
.A2(n_4007),
.A3(n_4011),
.B(n_4003),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4601),
.B(n_4481),
.Y(n_4987)
);

OAI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_4596),
.A2(n_2442),
.B(n_2391),
.Y(n_4988)
);

O2A1O1Ixp5_ASAP7_75t_SL g4989 ( 
.A1(n_4717),
.A2(n_4297),
.B(n_4298),
.C(n_4296),
.Y(n_4989)
);

OAI21x1_ASAP7_75t_L g4990 ( 
.A1(n_4604),
.A2(n_4467),
.B(n_4276),
.Y(n_4990)
);

AND2x2_ASAP7_75t_L g4991 ( 
.A(n_4586),
.B(n_4493),
.Y(n_4991)
);

OAI21x1_ASAP7_75t_L g4992 ( 
.A1(n_4626),
.A2(n_4277),
.B(n_4275),
.Y(n_4992)
);

OAI21xp5_ASAP7_75t_L g4993 ( 
.A1(n_4573),
.A2(n_1136),
.B(n_1132),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4570),
.B(n_4318),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4671),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4601),
.B(n_1139),
.Y(n_4996)
);

OAI21x1_ASAP7_75t_L g4997 ( 
.A1(n_4652),
.A2(n_4278),
.B(n_4515),
.Y(n_4997)
);

CKINVDCx5p33_ASAP7_75t_R g4998 ( 
.A(n_4645),
.Y(n_4998)
);

AO32x2_ASAP7_75t_L g4999 ( 
.A1(n_4644),
.A2(n_4507),
.A3(n_4399),
.B1(n_4338),
.B2(n_4299),
.Y(n_4999)
);

OAI21xp5_ASAP7_75t_L g5000 ( 
.A1(n_4660),
.A2(n_1154),
.B(n_1145),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4570),
.B(n_4381),
.Y(n_5001)
);

INVx2_ASAP7_75t_L g5002 ( 
.A(n_4610),
.Y(n_5002)
);

AO31x2_ASAP7_75t_L g5003 ( 
.A1(n_4679),
.A2(n_1390),
.A3(n_1391),
.B(n_1388),
.Y(n_5003)
);

OAI21x1_ASAP7_75t_L g5004 ( 
.A1(n_4874),
.A2(n_4413),
.B(n_4412),
.Y(n_5004)
);

AOI221xp5_ASAP7_75t_L g5005 ( 
.A1(n_4783),
.A2(n_1155),
.B1(n_1161),
.B2(n_1154),
.C(n_1145),
.Y(n_5005)
);

AOI21xp5_ASAP7_75t_L g5006 ( 
.A1(n_4705),
.A2(n_4390),
.B(n_4383),
.Y(n_5006)
);

AOI21xp5_ASAP7_75t_L g5007 ( 
.A1(n_4740),
.A2(n_4866),
.B(n_4792),
.Y(n_5007)
);

INVx5_ASAP7_75t_L g5008 ( 
.A(n_4906),
.Y(n_5008)
);

NOR2xp67_ASAP7_75t_L g5009 ( 
.A(n_4906),
.B(n_4391),
.Y(n_5009)
);

OAI21x1_ASAP7_75t_L g5010 ( 
.A1(n_4874),
.A2(n_4394),
.B(n_4392),
.Y(n_5010)
);

INVx2_ASAP7_75t_SL g5011 ( 
.A(n_4577),
.Y(n_5011)
);

AOI21xp5_ASAP7_75t_L g5012 ( 
.A1(n_4792),
.A2(n_4396),
.B(n_4395),
.Y(n_5012)
);

OAI21x1_ASAP7_75t_L g5013 ( 
.A1(n_4931),
.A2(n_4400),
.B(n_4361),
.Y(n_5013)
);

AOI221x1_ASAP7_75t_L g5014 ( 
.A1(n_4566),
.A2(n_4819),
.B1(n_4707),
.B2(n_4713),
.C(n_4741),
.Y(n_5014)
);

AOI21xp5_ASAP7_75t_L g5015 ( 
.A1(n_4866),
.A2(n_4418),
.B(n_4415),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4671),
.Y(n_5016)
);

AO21x2_ASAP7_75t_L g5017 ( 
.A1(n_4618),
.A2(n_4421),
.B(n_4419),
.Y(n_5017)
);

NOR2xp33_ASAP7_75t_L g5018 ( 
.A(n_4628),
.B(n_149),
.Y(n_5018)
);

OAI22xp5_ASAP7_75t_L g5019 ( 
.A1(n_4677),
.A2(n_1161),
.B1(n_1172),
.B2(n_1155),
.Y(n_5019)
);

AOI21xp5_ASAP7_75t_L g5020 ( 
.A1(n_4738),
.A2(n_4424),
.B(n_4423),
.Y(n_5020)
);

AOI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_4738),
.A2(n_4430),
.B(n_4429),
.Y(n_5021)
);

INVx2_ASAP7_75t_L g5022 ( 
.A(n_4621),
.Y(n_5022)
);

A2O1A1Ixp33_ASAP7_75t_L g5023 ( 
.A1(n_4803),
.A2(n_1187),
.B(n_1192),
.C(n_1172),
.Y(n_5023)
);

O2A1O1Ixp33_ASAP7_75t_L g5024 ( 
.A1(n_4785),
.A2(n_1187),
.B(n_1196),
.C(n_1192),
.Y(n_5024)
);

CKINVDCx8_ASAP7_75t_R g5025 ( 
.A(n_4734),
.Y(n_5025)
);

AOI221x1_ASAP7_75t_L g5026 ( 
.A1(n_4819),
.A2(n_1196),
.B1(n_1202),
.B2(n_1201),
.C(n_1197),
.Y(n_5026)
);

CKINVDCx5p33_ASAP7_75t_R g5027 ( 
.A(n_4574),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4624),
.B(n_1197),
.Y(n_5028)
);

INVx1_ASAP7_75t_SL g5029 ( 
.A(n_4577),
.Y(n_5029)
);

AOI21xp5_ASAP7_75t_L g5030 ( 
.A1(n_4749),
.A2(n_4434),
.B(n_4432),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4749),
.A2(n_4436),
.B(n_4435),
.Y(n_5031)
);

AND2x2_ASAP7_75t_L g5032 ( 
.A(n_4571),
.B(n_1201),
.Y(n_5032)
);

OAI21x1_ASAP7_75t_L g5033 ( 
.A1(n_4931),
.A2(n_4440),
.B(n_4438),
.Y(n_5033)
);

AO31x2_ASAP7_75t_L g5034 ( 
.A1(n_4699),
.A2(n_1393),
.A3(n_1394),
.B(n_1391),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_4766),
.B(n_149),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4585),
.Y(n_5036)
);

O2A1O1Ixp33_ASAP7_75t_L g5037 ( 
.A1(n_4872),
.A2(n_1202),
.B(n_1223),
.C(n_1213),
.Y(n_5037)
);

OAI21x1_ASAP7_75t_L g5038 ( 
.A1(n_4777),
.A2(n_4895),
.B(n_4609),
.Y(n_5038)
);

AOI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4764),
.A2(n_4442),
.B(n_2587),
.Y(n_5039)
);

AOI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4764),
.A2(n_2587),
.B(n_2581),
.Y(n_5040)
);

AO31x2_ASAP7_75t_L g5041 ( 
.A1(n_4833),
.A2(n_1394),
.A3(n_1395),
.B(n_1393),
.Y(n_5041)
);

OAI21x1_ASAP7_75t_L g5042 ( 
.A1(n_4609),
.A2(n_2842),
.B(n_2643),
.Y(n_5042)
);

INVx4_ASAP7_75t_L g5043 ( 
.A(n_4845),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4624),
.Y(n_5044)
);

A2O1A1Ixp33_ASAP7_75t_L g5045 ( 
.A1(n_4660),
.A2(n_1213),
.B(n_1228),
.C(n_1223),
.Y(n_5045)
);

O2A1O1Ixp33_ASAP7_75t_L g5046 ( 
.A1(n_4872),
.A2(n_1228),
.B(n_1234),
.C(n_1232),
.Y(n_5046)
);

AND2x2_ASAP7_75t_SL g5047 ( 
.A(n_4564),
.B(n_1232),
.Y(n_5047)
);

INVx3_ASAP7_75t_L g5048 ( 
.A(n_4587),
.Y(n_5048)
);

AOI21xp5_ASAP7_75t_L g5049 ( 
.A1(n_4862),
.A2(n_2587),
.B(n_2581),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4717),
.B(n_1234),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_4839),
.B(n_4592),
.Y(n_5051)
);

AO31x2_ASAP7_75t_L g5052 ( 
.A1(n_4880),
.A2(n_1396),
.A3(n_1397),
.B(n_1395),
.Y(n_5052)
);

NOR2xp67_ASAP7_75t_L g5053 ( 
.A(n_4906),
.B(n_1397),
.Y(n_5053)
);

OAI21xp5_ASAP7_75t_L g5054 ( 
.A1(n_4602),
.A2(n_3149),
.B(n_3073),
.Y(n_5054)
);

INVx2_ASAP7_75t_L g5055 ( 
.A(n_4638),
.Y(n_5055)
);

AO31x2_ASAP7_75t_L g5056 ( 
.A1(n_4720),
.A2(n_1402),
.A3(n_1403),
.B(n_1398),
.Y(n_5056)
);

BUFx10_ASAP7_75t_L g5057 ( 
.A(n_4713),
.Y(n_5057)
);

NOR2xp33_ASAP7_75t_L g5058 ( 
.A(n_4654),
.B(n_150),
.Y(n_5058)
);

AO31x2_ASAP7_75t_L g5059 ( 
.A1(n_4858),
.A2(n_1402),
.A3(n_1403),
.B(n_1398),
.Y(n_5059)
);

OAI21x1_ASAP7_75t_L g5060 ( 
.A1(n_4685),
.A2(n_2842),
.B(n_2643),
.Y(n_5060)
);

AOI21xp5_ASAP7_75t_L g5061 ( 
.A1(n_4862),
.A2(n_2587),
.B(n_2581),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4651),
.Y(n_5062)
);

AOI21xp5_ASAP7_75t_L g5063 ( 
.A1(n_4625),
.A2(n_2587),
.B(n_2861),
.Y(n_5063)
);

AOI21xp5_ASAP7_75t_L g5064 ( 
.A1(n_4625),
.A2(n_2872),
.B(n_2861),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4583),
.B(n_1404),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4651),
.Y(n_5066)
);

BUFx3_ASAP7_75t_L g5067 ( 
.A(n_4589),
.Y(n_5067)
);

OAI21x1_ASAP7_75t_L g5068 ( 
.A1(n_4575),
.A2(n_2854),
.B(n_2514),
.Y(n_5068)
);

AOI21xp5_ASAP7_75t_L g5069 ( 
.A1(n_4937),
.A2(n_2881),
.B(n_2872),
.Y(n_5069)
);

O2A1O1Ixp33_ASAP7_75t_L g5070 ( 
.A1(n_4689),
.A2(n_2308),
.B(n_2169),
.C(n_2158),
.Y(n_5070)
);

AND2x2_ASAP7_75t_L g5071 ( 
.A(n_4571),
.B(n_1404),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4608),
.B(n_1405),
.Y(n_5072)
);

AOI21xp5_ASAP7_75t_L g5073 ( 
.A1(n_4937),
.A2(n_2881),
.B(n_2872),
.Y(n_5073)
);

AOI21xp5_ASAP7_75t_L g5074 ( 
.A1(n_4718),
.A2(n_2881),
.B(n_2872),
.Y(n_5074)
);

OAI21x1_ASAP7_75t_L g5075 ( 
.A1(n_4917),
.A2(n_2854),
.B(n_2514),
.Y(n_5075)
);

INVx2_ASAP7_75t_SL g5076 ( 
.A(n_4595),
.Y(n_5076)
);

AOI21xp5_ASAP7_75t_L g5077 ( 
.A1(n_4718),
.A2(n_2894),
.B(n_2881),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4576),
.Y(n_5078)
);

AND2x4_ASAP7_75t_L g5079 ( 
.A(n_4594),
.B(n_1405),
.Y(n_5079)
);

AOI21xp5_ASAP7_75t_SL g5080 ( 
.A1(n_4728),
.A2(n_1409),
.B(n_1406),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_4629),
.B(n_1406),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4576),
.Y(n_5082)
);

HB1xp67_ASAP7_75t_L g5083 ( 
.A(n_4709),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4605),
.Y(n_5084)
);

AO31x2_ASAP7_75t_L g5085 ( 
.A1(n_4869),
.A2(n_1412),
.A3(n_1416),
.B(n_1409),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4567),
.B(n_4612),
.Y(n_5086)
);

CKINVDCx8_ASAP7_75t_R g5087 ( 
.A(n_4674),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4613),
.B(n_4622),
.Y(n_5088)
);

OAI22xp5_ASAP7_75t_L g5089 ( 
.A1(n_4677),
.A2(n_831),
.B1(n_836),
.B2(n_827),
.Y(n_5089)
);

NOR3xp33_ASAP7_75t_L g5090 ( 
.A(n_4563),
.B(n_1181),
.C(n_836),
.Y(n_5090)
);

OAI21x1_ASAP7_75t_L g5091 ( 
.A1(n_4917),
.A2(n_2514),
.B(n_2510),
.Y(n_5091)
);

BUFx8_ASAP7_75t_L g5092 ( 
.A(n_4876),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4627),
.Y(n_5093)
);

BUFx4_ASAP7_75t_SL g5094 ( 
.A(n_4781),
.Y(n_5094)
);

AOI22xp33_ASAP7_75t_L g5095 ( 
.A1(n_4606),
.A2(n_3149),
.B1(n_3175),
.B2(n_3073),
.Y(n_5095)
);

AOI221xp5_ASAP7_75t_L g5096 ( 
.A1(n_4783),
.A2(n_879),
.B1(n_887),
.B2(n_885),
.C(n_875),
.Y(n_5096)
);

INVx1_ASAP7_75t_SL g5097 ( 
.A(n_4595),
.Y(n_5097)
);

A2O1A1Ixp33_ASAP7_75t_L g5098 ( 
.A1(n_4606),
.A2(n_1189),
.B(n_1218),
.C(n_840),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4630),
.Y(n_5099)
);

OAI21x1_ASAP7_75t_L g5100 ( 
.A1(n_4756),
.A2(n_2540),
.B(n_2510),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_4639),
.Y(n_5101)
);

INVx3_ASAP7_75t_L g5102 ( 
.A(n_4619),
.Y(n_5102)
);

AND2x2_ASAP7_75t_L g5103 ( 
.A(n_4709),
.B(n_1412),
.Y(n_5103)
);

INVx3_ASAP7_75t_L g5104 ( 
.A(n_4619),
.Y(n_5104)
);

A2O1A1Ixp33_ASAP7_75t_L g5105 ( 
.A1(n_4691),
.A2(n_1189),
.B(n_1218),
.C(n_840),
.Y(n_5105)
);

AOI21xp33_ASAP7_75t_L g5106 ( 
.A1(n_4569),
.A2(n_1465),
.B(n_1416),
.Y(n_5106)
);

OAI21x1_ASAP7_75t_L g5107 ( 
.A1(n_4789),
.A2(n_2543),
.B(n_2540),
.Y(n_5107)
);

AOI221x1_ASAP7_75t_L g5108 ( 
.A1(n_4707),
.A2(n_1634),
.B1(n_1636),
.B2(n_1632),
.C(n_1465),
.Y(n_5108)
);

NAND2xp5_ASAP7_75t_L g5109 ( 
.A(n_4715),
.B(n_1632),
.Y(n_5109)
);

HB1xp67_ASAP7_75t_L g5110 ( 
.A(n_4686),
.Y(n_5110)
);

BUFx6f_ASAP7_75t_L g5111 ( 
.A(n_4600),
.Y(n_5111)
);

O2A1O1Ixp5_ASAP7_75t_L g5112 ( 
.A1(n_4597),
.A2(n_1636),
.B(n_1637),
.C(n_1634),
.Y(n_5112)
);

A2O1A1Ixp33_ASAP7_75t_L g5113 ( 
.A1(n_4691),
.A2(n_1077),
.B(n_1180),
.C(n_949),
.Y(n_5113)
);

INVx2_ASAP7_75t_L g5114 ( 
.A(n_4656),
.Y(n_5114)
);

NOR2xp67_ASAP7_75t_L g5115 ( 
.A(n_4906),
.B(n_1637),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_4715),
.B(n_1638),
.Y(n_5116)
);

INVx2_ASAP7_75t_SL g5117 ( 
.A(n_4658),
.Y(n_5117)
);

OAI21x1_ASAP7_75t_L g5118 ( 
.A1(n_4861),
.A2(n_2543),
.B(n_2540),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_SL g5119 ( 
.A(n_4845),
.B(n_1638),
.Y(n_5119)
);

AOI221x1_ASAP7_75t_L g5120 ( 
.A1(n_4741),
.A2(n_1644),
.B1(n_1646),
.B2(n_1643),
.C(n_1642),
.Y(n_5120)
);

OAI21x1_ASAP7_75t_L g5121 ( 
.A1(n_4672),
.A2(n_2549),
.B(n_2543),
.Y(n_5121)
);

NOR2xp33_ASAP7_75t_L g5122 ( 
.A(n_4729),
.B(n_150),
.Y(n_5122)
);

AO31x2_ASAP7_75t_L g5123 ( 
.A1(n_4884),
.A2(n_1643),
.A3(n_1644),
.B(n_1642),
.Y(n_5123)
);

O2A1O1Ixp33_ASAP7_75t_SL g5124 ( 
.A1(n_4669),
.A2(n_2275),
.B(n_2284),
.C(n_2264),
.Y(n_5124)
);

BUFx3_ASAP7_75t_L g5125 ( 
.A(n_4736),
.Y(n_5125)
);

O2A1O1Ixp5_ASAP7_75t_L g5126 ( 
.A1(n_4597),
.A2(n_1649),
.B(n_1650),
.C(n_1646),
.Y(n_5126)
);

NOR2xp33_ASAP7_75t_SL g5127 ( 
.A(n_4737),
.B(n_3073),
.Y(n_5127)
);

NAND3xp33_ASAP7_75t_L g5128 ( 
.A(n_4636),
.B(n_1177),
.C(n_1114),
.Y(n_5128)
);

CKINVDCx5p33_ASAP7_75t_R g5129 ( 
.A(n_4892),
.Y(n_5129)
);

AOI21xp5_ASAP7_75t_L g5130 ( 
.A1(n_4716),
.A2(n_2894),
.B(n_2881),
.Y(n_5130)
);

OR2x2_ASAP7_75t_L g5131 ( 
.A(n_4578),
.B(n_4665),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4607),
.B(n_1649),
.Y(n_5132)
);

BUFx6f_ASAP7_75t_L g5133 ( 
.A(n_4600),
.Y(n_5133)
);

OAI21x1_ASAP7_75t_L g5134 ( 
.A1(n_4966),
.A2(n_2550),
.B(n_2549),
.Y(n_5134)
);

NOR2xp33_ASAP7_75t_L g5135 ( 
.A(n_4581),
.B(n_153),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_4659),
.Y(n_5136)
);

NOR2xp67_ASAP7_75t_L g5137 ( 
.A(n_4860),
.B(n_1650),
.Y(n_5137)
);

AOI21xp5_ASAP7_75t_L g5138 ( 
.A1(n_4860),
.A2(n_4944),
.B(n_4914),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_4667),
.B(n_1651),
.Y(n_5139)
);

OR2x2_ASAP7_75t_L g5140 ( 
.A(n_4641),
.B(n_1651),
.Y(n_5140)
);

INVx2_ASAP7_75t_SL g5141 ( 
.A(n_4565),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4620),
.B(n_1652),
.Y(n_5142)
);

AOI21xp5_ASAP7_75t_L g5143 ( 
.A1(n_4898),
.A2(n_2894),
.B(n_2625),
.Y(n_5143)
);

AOI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_4750),
.A2(n_3073),
.B1(n_3264),
.B2(n_3175),
.Y(n_5144)
);

A2O1A1Ixp33_ASAP7_75t_L g5145 ( 
.A1(n_4703),
.A2(n_1077),
.B(n_1180),
.C(n_949),
.Y(n_5145)
);

A2O1A1Ixp33_ASAP7_75t_L g5146 ( 
.A1(n_4703),
.A2(n_1183),
.B(n_1182),
.C(n_1181),
.Y(n_5146)
);

OAI22xp5_ASAP7_75t_L g5147 ( 
.A1(n_4735),
.A2(n_4675),
.B1(n_4688),
.B2(n_4923),
.Y(n_5147)
);

INVx2_ASAP7_75t_SL g5148 ( 
.A(n_4582),
.Y(n_5148)
);

AO31x2_ASAP7_75t_L g5149 ( 
.A1(n_4805),
.A2(n_1653),
.A3(n_1658),
.B(n_1652),
.Y(n_5149)
);

A2O1A1Ixp33_ASAP7_75t_L g5150 ( 
.A1(n_4572),
.A2(n_1214),
.B(n_1185),
.C(n_1183),
.Y(n_5150)
);

INVx5_ASAP7_75t_L g5151 ( 
.A(n_4643),
.Y(n_5151)
);

AOI22xp33_ASAP7_75t_L g5152 ( 
.A1(n_4735),
.A2(n_3264),
.B1(n_3285),
.B2(n_3175),
.Y(n_5152)
);

O2A1O1Ixp33_ASAP7_75t_L g5153 ( 
.A1(n_4758),
.A2(n_2284),
.B(n_2288),
.C(n_2275),
.Y(n_5153)
);

AND2x4_ASAP7_75t_L g5154 ( 
.A(n_4632),
.B(n_1653),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_L g5155 ( 
.A(n_4681),
.B(n_1658),
.Y(n_5155)
);

OAI21x1_ASAP7_75t_L g5156 ( 
.A1(n_4966),
.A2(n_2550),
.B(n_2549),
.Y(n_5156)
);

BUFx2_ASAP7_75t_SL g5157 ( 
.A(n_4614),
.Y(n_5157)
);

A2O1A1Ixp33_ASAP7_75t_L g5158 ( 
.A1(n_4572),
.A2(n_1188),
.B(n_1185),
.C(n_1182),
.Y(n_5158)
);

OAI21x1_ASAP7_75t_L g5159 ( 
.A1(n_4968),
.A2(n_2550),
.B(n_2487),
.Y(n_5159)
);

OAI21x1_ASAP7_75t_L g5160 ( 
.A1(n_4968),
.A2(n_2487),
.B(n_2792),
.Y(n_5160)
);

BUFx6f_ASAP7_75t_L g5161 ( 
.A(n_4600),
.Y(n_5161)
);

OAI21x1_ASAP7_75t_L g5162 ( 
.A1(n_4900),
.A2(n_2487),
.B(n_2798),
.Y(n_5162)
);

AOI31xp67_ASAP7_75t_L g5163 ( 
.A1(n_4945),
.A2(n_4899),
.A3(n_4902),
.B(n_4908),
.Y(n_5163)
);

BUFx4f_ASAP7_75t_SL g5164 ( 
.A(n_4896),
.Y(n_5164)
);

HB1xp67_ASAP7_75t_L g5165 ( 
.A(n_4686),
.Y(n_5165)
);

A2O1A1Ixp33_ASAP7_75t_L g5166 ( 
.A1(n_4563),
.A2(n_1214),
.B(n_1188),
.C(n_1660),
.Y(n_5166)
);

A2O1A1Ixp33_ASAP7_75t_L g5167 ( 
.A1(n_4853),
.A2(n_1663),
.B(n_1666),
.C(n_1661),
.Y(n_5167)
);

AOI22xp5_ASAP7_75t_L g5168 ( 
.A1(n_4580),
.A2(n_3264),
.B1(n_3350),
.B2(n_3285),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4649),
.Y(n_5169)
);

AOI21xp5_ASAP7_75t_L g5170 ( 
.A1(n_4680),
.A2(n_2894),
.B(n_2625),
.Y(n_5170)
);

INVx3_ASAP7_75t_L g5171 ( 
.A(n_4632),
.Y(n_5171)
);

AO32x2_ASAP7_75t_L g5172 ( 
.A1(n_4793),
.A2(n_2352),
.A3(n_1669),
.B1(n_1673),
.B2(n_1667),
.Y(n_5172)
);

OAI21x1_ASAP7_75t_L g5173 ( 
.A1(n_4900),
.A2(n_2818),
.B(n_2798),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_4568),
.Y(n_5174)
);

AOI21xp5_ASAP7_75t_L g5175 ( 
.A1(n_4711),
.A2(n_2894),
.B(n_2628),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4655),
.Y(n_5176)
);

AO31x2_ASAP7_75t_L g5177 ( 
.A1(n_4666),
.A2(n_4854),
.A3(n_4849),
.B(n_4915),
.Y(n_5177)
);

AND2x2_ASAP7_75t_L g5178 ( 
.A(n_4744),
.B(n_1666),
.Y(n_5178)
);

NAND2xp5_ASAP7_75t_L g5179 ( 
.A(n_4631),
.B(n_1667),
.Y(n_5179)
);

AND2x4_ASAP7_75t_L g5180 ( 
.A(n_4697),
.B(n_1669),
.Y(n_5180)
);

AND2x4_ASAP7_75t_L g5181 ( 
.A(n_4697),
.B(n_1674),
.Y(n_5181)
);

O2A1O1Ixp5_ASAP7_75t_L g5182 ( 
.A1(n_4963),
.A2(n_1674),
.B(n_1421),
.C(n_1424),
.Y(n_5182)
);

AOI22xp33_ASAP7_75t_L g5183 ( 
.A1(n_4675),
.A2(n_3285),
.B1(n_3350),
.B2(n_3264),
.Y(n_5183)
);

BUFx12f_ASAP7_75t_L g5184 ( 
.A(n_4798),
.Y(n_5184)
);

AO22x1_ASAP7_75t_L g5185 ( 
.A1(n_4581),
.A2(n_3285),
.B1(n_3350),
.B2(n_3264),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_4662),
.Y(n_5186)
);

INVx4_ASAP7_75t_L g5187 ( 
.A(n_4727),
.Y(n_5187)
);

AND2x4_ASAP7_75t_L g5188 ( 
.A(n_4757),
.B(n_1417),
.Y(n_5188)
);

OAI21x1_ASAP7_75t_L g5189 ( 
.A1(n_4973),
.A2(n_2819),
.B(n_2818),
.Y(n_5189)
);

AOI21xp5_ASAP7_75t_L g5190 ( 
.A1(n_4782),
.A2(n_2628),
.B(n_2624),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_4832),
.B(n_1421),
.Y(n_5191)
);

AOI21xp5_ASAP7_75t_L g5192 ( 
.A1(n_4782),
.A2(n_2630),
.B(n_2819),
.Y(n_5192)
);

OAI22xp5_ASAP7_75t_L g5193 ( 
.A1(n_4688),
.A2(n_4923),
.B1(n_4816),
.B2(n_4788),
.Y(n_5193)
);

OAI21x1_ASAP7_75t_L g5194 ( 
.A1(n_4907),
.A2(n_2824),
.B(n_2821),
.Y(n_5194)
);

BUFx2_ASAP7_75t_L g5195 ( 
.A(n_4730),
.Y(n_5195)
);

BUFx2_ASAP7_75t_R g5196 ( 
.A(n_4964),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4694),
.Y(n_5197)
);

OAI21x1_ASAP7_75t_L g5198 ( 
.A1(n_4924),
.A2(n_2824),
.B(n_2821),
.Y(n_5198)
);

OAI22xp5_ASAP7_75t_L g5199 ( 
.A1(n_4816),
.A2(n_1177),
.B1(n_1198),
.B2(n_1114),
.Y(n_5199)
);

INVx2_ASAP7_75t_L g5200 ( 
.A(n_4712),
.Y(n_5200)
);

AOI21xp5_ASAP7_75t_L g5201 ( 
.A1(n_4588),
.A2(n_4698),
.B(n_4901),
.Y(n_5201)
);

NOR2xp33_ASAP7_75t_L g5202 ( 
.A(n_4615),
.B(n_153),
.Y(n_5202)
);

INVx2_ASAP7_75t_L g5203 ( 
.A(n_4719),
.Y(n_5203)
);

AO21x1_ASAP7_75t_L g5204 ( 
.A1(n_4857),
.A2(n_919),
.B(n_1335),
.Y(n_5204)
);

A2O1A1Ixp33_ASAP7_75t_L g5205 ( 
.A1(n_4853),
.A2(n_889),
.B(n_894),
.C(n_888),
.Y(n_5205)
);

AOI21xp5_ASAP7_75t_L g5206 ( 
.A1(n_4588),
.A2(n_2630),
.B(n_2825),
.Y(n_5206)
);

AO31x2_ASAP7_75t_L g5207 ( 
.A1(n_4856),
.A2(n_3028),
.A3(n_3043),
.B(n_3019),
.Y(n_5207)
);

OAI21x1_ASAP7_75t_L g5208 ( 
.A1(n_4924),
.A2(n_2837),
.B(n_2825),
.Y(n_5208)
);

INVx3_ASAP7_75t_L g5209 ( 
.A(n_4757),
.Y(n_5209)
);

AO21x1_ASAP7_75t_L g5210 ( 
.A1(n_4857),
.A2(n_4795),
.B(n_4830),
.Y(n_5210)
);

AOI21xp5_ASAP7_75t_L g5211 ( 
.A1(n_4698),
.A2(n_2850),
.B(n_2837),
.Y(n_5211)
);

AOI221xp5_ASAP7_75t_L g5212 ( 
.A1(n_4650),
.A2(n_898),
.B1(n_899),
.B2(n_897),
.C(n_892),
.Y(n_5212)
);

AOI221x1_ASAP7_75t_L g5213 ( 
.A1(n_4814),
.A2(n_1198),
.B1(n_1177),
.B2(n_1114),
.C(n_1335),
.Y(n_5213)
);

AO21x1_ASAP7_75t_L g5214 ( 
.A1(n_4795),
.A2(n_919),
.B(n_1340),
.Y(n_5214)
);

AOI221xp5_ASAP7_75t_L g5215 ( 
.A1(n_4650),
.A2(n_907),
.B1(n_908),
.B2(n_901),
.C(n_900),
.Y(n_5215)
);

AO31x2_ASAP7_75t_L g5216 ( 
.A1(n_4919),
.A2(n_3028),
.A3(n_3043),
.B(n_3019),
.Y(n_5216)
);

BUFx2_ASAP7_75t_L g5217 ( 
.A(n_4852),
.Y(n_5217)
);

OAI21x1_ASAP7_75t_L g5218 ( 
.A1(n_4953),
.A2(n_2871),
.B(n_2850),
.Y(n_5218)
);

AOI21xp5_ASAP7_75t_L g5219 ( 
.A1(n_4901),
.A2(n_2884),
.B(n_2871),
.Y(n_5219)
);

INVx1_ASAP7_75t_SL g5220 ( 
.A(n_4897),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_4788),
.B(n_1114),
.Y(n_5221)
);

BUFx3_ASAP7_75t_L g5222 ( 
.A(n_4733),
.Y(n_5222)
);

OAI21x1_ASAP7_75t_L g5223 ( 
.A1(n_4887),
.A2(n_2892),
.B(n_2884),
.Y(n_5223)
);

AND2x4_ASAP7_75t_L g5224 ( 
.A(n_4762),
.B(n_4768),
.Y(n_5224)
);

CKINVDCx20_ASAP7_75t_R g5225 ( 
.A(n_4952),
.Y(n_5225)
);

INVx2_ASAP7_75t_L g5226 ( 
.A(n_4702),
.Y(n_5226)
);

AO31x2_ASAP7_75t_L g5227 ( 
.A1(n_4938),
.A2(n_3069),
.A3(n_3072),
.B(n_3052),
.Y(n_5227)
);

OAI22x1_ASAP7_75t_L g5228 ( 
.A1(n_4623),
.A2(n_915),
.B1(n_917),
.B2(n_911),
.Y(n_5228)
);

OA21x2_ASAP7_75t_L g5229 ( 
.A1(n_4879),
.A2(n_1433),
.B(n_1424),
.Y(n_5229)
);

AOI21x1_ASAP7_75t_SL g5230 ( 
.A1(n_4807),
.A2(n_7),
.B(n_8),
.Y(n_5230)
);

OAI21x1_ASAP7_75t_L g5231 ( 
.A1(n_4887),
.A2(n_2919),
.B(n_2892),
.Y(n_5231)
);

BUFx6f_ASAP7_75t_L g5232 ( 
.A(n_4600),
.Y(n_5232)
);

AOI21xp5_ASAP7_75t_L g5233 ( 
.A1(n_4963),
.A2(n_4945),
.B(n_4569),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_4885),
.B(n_1114),
.Y(n_5234)
);

OAI21x1_ASAP7_75t_L g5235 ( 
.A1(n_4704),
.A2(n_2919),
.B(n_3052),
.Y(n_5235)
);

AOI21xp5_ASAP7_75t_L g5236 ( 
.A1(n_4683),
.A2(n_3285),
.B(n_3264),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_4706),
.Y(n_5237)
);

AND2x4_ASAP7_75t_L g5238 ( 
.A(n_4762),
.B(n_4724),
.Y(n_5238)
);

OAI21x1_ASAP7_75t_L g5239 ( 
.A1(n_4648),
.A2(n_3072),
.B(n_3069),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4690),
.Y(n_5240)
);

NOR2xp33_ASAP7_75t_L g5241 ( 
.A(n_4682),
.B(n_154),
.Y(n_5241)
);

AOI21xp5_ASAP7_75t_L g5242 ( 
.A1(n_4683),
.A2(n_3350),
.B(n_3285),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_4739),
.Y(n_5243)
);

NAND2xp5_ASAP7_75t_L g5244 ( 
.A(n_4885),
.B(n_1114),
.Y(n_5244)
);

OR2x2_ASAP7_75t_L g5245 ( 
.A(n_4584),
.B(n_1433),
.Y(n_5245)
);

OAI22xp5_ASAP7_75t_L g5246 ( 
.A1(n_4834),
.A2(n_1198),
.B1(n_1177),
.B2(n_918),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_4920),
.Y(n_5247)
);

INVx3_ASAP7_75t_L g5248 ( 
.A(n_4950),
.Y(n_5248)
);

NAND3xp33_ASAP7_75t_L g5249 ( 
.A(n_4913),
.B(n_1198),
.C(n_1177),
.Y(n_5249)
);

AOI21xp5_ASAP7_75t_L g5250 ( 
.A1(n_4879),
.A2(n_3350),
.B(n_2518),
.Y(n_5250)
);

AO31x2_ASAP7_75t_L g5251 ( 
.A1(n_4946),
.A2(n_3081),
.A3(n_3090),
.B(n_3079),
.Y(n_5251)
);

OAI21x1_ASAP7_75t_SL g5252 ( 
.A1(n_4859),
.A2(n_4791),
.B(n_4841),
.Y(n_5252)
);

AO31x2_ASAP7_75t_L g5253 ( 
.A1(n_4882),
.A2(n_3081),
.A3(n_3090),
.B(n_3079),
.Y(n_5253)
);

AOI22xp5_ASAP7_75t_SL g5254 ( 
.A1(n_4643),
.A2(n_922),
.B1(n_926),
.B2(n_916),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_4701),
.B(n_4714),
.Y(n_5255)
);

O2A1O1Ixp33_ASAP7_75t_L g5256 ( 
.A1(n_4759),
.A2(n_2289),
.B(n_2291),
.C(n_2288),
.Y(n_5256)
);

AOI22xp33_ASAP7_75t_SL g5257 ( 
.A1(n_4693),
.A2(n_1198),
.B1(n_1177),
.B2(n_935),
.Y(n_5257)
);

INVx2_ASAP7_75t_L g5258 ( 
.A(n_4935),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_L g5259 ( 
.A(n_4739),
.B(n_1434),
.Y(n_5259)
);

INVx2_ASAP7_75t_SL g5260 ( 
.A(n_4635),
.Y(n_5260)
);

CKINVDCx20_ASAP7_75t_R g5261 ( 
.A(n_4911),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_L g5262 ( 
.A(n_4742),
.B(n_1434),
.Y(n_5262)
);

HB1xp67_ASAP7_75t_L g5263 ( 
.A(n_4684),
.Y(n_5263)
);

INVxp67_ASAP7_75t_L g5264 ( 
.A(n_4593),
.Y(n_5264)
);

NOR2xp33_ASAP7_75t_L g5265 ( 
.A(n_4603),
.B(n_154),
.Y(n_5265)
);

OAI22xp5_ASAP7_75t_L g5266 ( 
.A1(n_4834),
.A2(n_1198),
.B1(n_1177),
.B2(n_936),
.Y(n_5266)
);

BUFx4f_ASAP7_75t_SL g5267 ( 
.A(n_4896),
.Y(n_5267)
);

AOI21x1_ASAP7_75t_L g5268 ( 
.A1(n_4821),
.A2(n_1455),
.B(n_1449),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_4835),
.B(n_1198),
.Y(n_5269)
);

AOI21xp5_ASAP7_75t_L g5270 ( 
.A1(n_4978),
.A2(n_2518),
.B(n_2517),
.Y(n_5270)
);

OAI21xp5_ASAP7_75t_SL g5271 ( 
.A1(n_4657),
.A2(n_158),
.B(n_156),
.Y(n_5271)
);

O2A1O1Ixp33_ASAP7_75t_L g5272 ( 
.A1(n_4958),
.A2(n_2291),
.B(n_2294),
.C(n_2289),
.Y(n_5272)
);

O2A1O1Ixp33_ASAP7_75t_L g5273 ( 
.A1(n_4961),
.A2(n_2296),
.B(n_2303),
.C(n_2294),
.Y(n_5273)
);

AO31x2_ASAP7_75t_L g5274 ( 
.A1(n_4909),
.A2(n_4903),
.A3(n_4927),
.B(n_4867),
.Y(n_5274)
);

OAI22xp5_ASAP7_75t_L g5275 ( 
.A1(n_4771),
.A2(n_937),
.B1(n_945),
.B2(n_929),
.Y(n_5275)
);

AND2x2_ASAP7_75t_L g5276 ( 
.A(n_4661),
.B(n_8),
.Y(n_5276)
);

AO31x2_ASAP7_75t_L g5277 ( 
.A1(n_4960),
.A2(n_3106),
.A3(n_3109),
.B(n_3104),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_4742),
.Y(n_5278)
);

AOI21xp5_ASAP7_75t_L g5279 ( 
.A1(n_4800),
.A2(n_4692),
.B(n_4893),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_4806),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_4806),
.Y(n_5281)
);

AOI21xp5_ASAP7_75t_L g5282 ( 
.A1(n_4800),
.A2(n_2519),
.B(n_2517),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_4904),
.Y(n_5283)
);

AO31x2_ASAP7_75t_L g5284 ( 
.A1(n_4979),
.A2(n_3106),
.A3(n_3109),
.B(n_3104),
.Y(n_5284)
);

AO21x2_ASAP7_75t_L g5285 ( 
.A1(n_4910),
.A2(n_2303),
.B(n_2296),
.Y(n_5285)
);

OAI21x1_ASAP7_75t_L g5286 ( 
.A1(n_4886),
.A2(n_3115),
.B(n_3110),
.Y(n_5286)
);

AOI221x1_ASAP7_75t_L g5287 ( 
.A1(n_4926),
.A2(n_1340),
.B1(n_1347),
.B2(n_1346),
.C(n_1341),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4692),
.A2(n_2525),
.B(n_2519),
.Y(n_5288)
);

AO31x2_ASAP7_75t_L g5289 ( 
.A1(n_4981),
.A2(n_4696),
.A3(n_4848),
.B(n_4842),
.Y(n_5289)
);

OAI21xp5_ASAP7_75t_L g5290 ( 
.A1(n_4812),
.A2(n_950),
.B(n_946),
.Y(n_5290)
);

INVx2_ASAP7_75t_SL g5291 ( 
.A(n_4653),
.Y(n_5291)
);

OAI22xp5_ASAP7_75t_L g5292 ( 
.A1(n_4771),
.A2(n_965),
.B1(n_966),
.B2(n_953),
.Y(n_5292)
);

AOI21xp5_ASAP7_75t_L g5293 ( 
.A1(n_4975),
.A2(n_2527),
.B(n_2525),
.Y(n_5293)
);

OAI22xp5_ASAP7_75t_SL g5294 ( 
.A1(n_4748),
.A2(n_969),
.B1(n_975),
.B2(n_967),
.Y(n_5294)
);

OAI21x1_ASAP7_75t_L g5295 ( 
.A1(n_4844),
.A2(n_3115),
.B(n_3110),
.Y(n_5295)
);

OA21x2_ASAP7_75t_L g5296 ( 
.A1(n_4954),
.A2(n_4918),
.B(n_4664),
.Y(n_5296)
);

OAI21x1_ASAP7_75t_L g5297 ( 
.A1(n_4844),
.A2(n_3122),
.B(n_3118),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4904),
.Y(n_5298)
);

NAND2xp33_ASAP7_75t_SL g5299 ( 
.A(n_4634),
.B(n_4663),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_L g5300 ( 
.A1(n_4954),
.A2(n_2531),
.B(n_2527),
.Y(n_5300)
);

AOI31xp67_ASAP7_75t_L g5301 ( 
.A1(n_4847),
.A2(n_1449),
.A3(n_1470),
.B(n_1455),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_4838),
.B(n_9),
.Y(n_5302)
);

OA21x2_ASAP7_75t_L g5303 ( 
.A1(n_4918),
.A2(n_1485),
.B(n_1470),
.Y(n_5303)
);

CKINVDCx11_ASAP7_75t_R g5304 ( 
.A(n_4723),
.Y(n_5304)
);

OAI21x1_ASAP7_75t_L g5305 ( 
.A1(n_4889),
.A2(n_3122),
.B(n_3118),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_4840),
.B(n_9),
.Y(n_5306)
);

O2A1O1Ixp33_ASAP7_75t_L g5307 ( 
.A1(n_4830),
.A2(n_2305),
.B(n_2196),
.C(n_2197),
.Y(n_5307)
);

INVx2_ASAP7_75t_L g5308 ( 
.A(n_4752),
.Y(n_5308)
);

BUFx3_ASAP7_75t_L g5309 ( 
.A(n_4760),
.Y(n_5309)
);

AND2x2_ASAP7_75t_L g5310 ( 
.A(n_4579),
.B(n_4663),
.Y(n_5310)
);

OAI21x1_ASAP7_75t_L g5311 ( 
.A1(n_4889),
.A2(n_3136),
.B(n_3123),
.Y(n_5311)
);

CKINVDCx20_ASAP7_75t_R g5312 ( 
.A(n_4637),
.Y(n_5312)
);

NOR2x1_ASAP7_75t_SL g5313 ( 
.A(n_4668),
.B(n_2531),
.Y(n_5313)
);

OAI21x1_ASAP7_75t_L g5314 ( 
.A1(n_4780),
.A2(n_3136),
.B(n_3123),
.Y(n_5314)
);

AOI22xp5_ASAP7_75t_L g5315 ( 
.A1(n_4743),
.A2(n_979),
.B1(n_981),
.B2(n_978),
.Y(n_5315)
);

AO22x2_ASAP7_75t_L g5316 ( 
.A1(n_4687),
.A2(n_2533),
.B1(n_2535),
.B2(n_2532),
.Y(n_5316)
);

NAND2xp5_ASAP7_75t_L g5317 ( 
.A(n_4684),
.B(n_1485),
.Y(n_5317)
);

BUFx10_ASAP7_75t_L g5318 ( 
.A(n_4921),
.Y(n_5318)
);

AOI21xp5_ASAP7_75t_L g5319 ( 
.A1(n_4949),
.A2(n_2533),
.B(n_2532),
.Y(n_5319)
);

INVx2_ASAP7_75t_SL g5320 ( 
.A(n_4653),
.Y(n_5320)
);

OR2x2_ASAP7_75t_L g5321 ( 
.A(n_4829),
.B(n_1499),
.Y(n_5321)
);

O2A1O1Ixp5_ASAP7_75t_L g5322 ( 
.A1(n_4976),
.A2(n_1507),
.B(n_1508),
.C(n_1499),
.Y(n_5322)
);

BUFx2_ASAP7_75t_R g5323 ( 
.A(n_4746),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_4747),
.B(n_1507),
.Y(n_5324)
);

NOR2xp33_ASAP7_75t_L g5325 ( 
.A(n_4668),
.B(n_156),
.Y(n_5325)
);

BUFx2_ASAP7_75t_L g5326 ( 
.A(n_4967),
.Y(n_5326)
);

AND2x4_ASAP7_75t_L g5327 ( 
.A(n_4724),
.B(n_1508),
.Y(n_5327)
);

OAI21x1_ASAP7_75t_L g5328 ( 
.A1(n_4930),
.A2(n_3159),
.B(n_3157),
.Y(n_5328)
);

NOR2xp33_ASAP7_75t_L g5329 ( 
.A(n_4710),
.B(n_4634),
.Y(n_5329)
);

A2O1A1Ixp33_ASAP7_75t_L g5330 ( 
.A1(n_4590),
.A2(n_987),
.B(n_990),
.C(n_983),
.Y(n_5330)
);

OAI22xp33_ASAP7_75t_L g5331 ( 
.A1(n_4826),
.A2(n_3333),
.B1(n_3377),
.B2(n_3320),
.Y(n_5331)
);

AO31x2_ASAP7_75t_L g5332 ( 
.A1(n_4932),
.A2(n_3159),
.A3(n_3176),
.B(n_3157),
.Y(n_5332)
);

INVx2_ASAP7_75t_L g5333 ( 
.A(n_4813),
.Y(n_5333)
);

AND2x4_ASAP7_75t_L g5334 ( 
.A(n_4724),
.B(n_1531),
.Y(n_5334)
);

NAND2x1p5_ASAP7_75t_L g5335 ( 
.A(n_4598),
.B(n_3320),
.Y(n_5335)
);

AOI21xp5_ASAP7_75t_L g5336 ( 
.A1(n_4807),
.A2(n_2537),
.B(n_2535),
.Y(n_5336)
);

AO31x2_ASAP7_75t_L g5337 ( 
.A1(n_4850),
.A2(n_3178),
.A3(n_3185),
.B(n_3176),
.Y(n_5337)
);

OAI21x1_ASAP7_75t_L g5338 ( 
.A1(n_4930),
.A2(n_3185),
.B(n_3178),
.Y(n_5338)
);

AOI21xp5_ASAP7_75t_L g5339 ( 
.A1(n_4878),
.A2(n_2542),
.B(n_2537),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_L g5340 ( 
.A(n_4864),
.B(n_9),
.Y(n_5340)
);

AND3x2_ASAP7_75t_L g5341 ( 
.A(n_4921),
.B(n_4868),
.C(n_4878),
.Y(n_5341)
);

A2O1A1Ixp33_ASAP7_75t_L g5342 ( 
.A1(n_4590),
.A2(n_992),
.B(n_997),
.C(n_993),
.Y(n_5342)
);

INVx2_ASAP7_75t_L g5343 ( 
.A(n_4797),
.Y(n_5343)
);

BUFx12f_ASAP7_75t_L g5344 ( 
.A(n_4633),
.Y(n_5344)
);

INVx2_ASAP7_75t_L g5345 ( 
.A(n_4799),
.Y(n_5345)
);

A2O1A1Ixp33_ASAP7_75t_L g5346 ( 
.A1(n_4883),
.A2(n_998),
.B(n_1005),
.C(n_1004),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4695),
.Y(n_5347)
);

AOI21xp5_ASAP7_75t_L g5348 ( 
.A1(n_4868),
.A2(n_4972),
.B(n_4875),
.Y(n_5348)
);

NAND2xp5_ASAP7_75t_L g5349 ( 
.A(n_4753),
.B(n_1531),
.Y(n_5349)
);

BUFx2_ASAP7_75t_L g5350 ( 
.A(n_4925),
.Y(n_5350)
);

INVx3_ASAP7_75t_SL g5351 ( 
.A(n_4710),
.Y(n_5351)
);

AOI221xp5_ASAP7_75t_L g5352 ( 
.A1(n_4599),
.A2(n_1008),
.B1(n_1010),
.B2(n_1006),
.C(n_991),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_4871),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_4881),
.Y(n_5354)
);

OAI21x1_ASAP7_75t_L g5355 ( 
.A1(n_4673),
.A2(n_3206),
.B(n_3199),
.Y(n_5355)
);

O2A1O1Ixp5_ASAP7_75t_SL g5356 ( 
.A1(n_4962),
.A2(n_1346),
.B(n_1347),
.C(n_1341),
.Y(n_5356)
);

BUFx6f_ASAP7_75t_L g5357 ( 
.A(n_4616),
.Y(n_5357)
);

AOI22xp5_ASAP7_75t_L g5358 ( 
.A1(n_4721),
.A2(n_1012),
.B1(n_1013),
.B2(n_1011),
.Y(n_5358)
);

AND2x2_ASAP7_75t_L g5359 ( 
.A(n_4786),
.B(n_10),
.Y(n_5359)
);

AO31x2_ASAP7_75t_L g5360 ( 
.A1(n_4855),
.A2(n_3206),
.A3(n_3211),
.B(n_3199),
.Y(n_5360)
);

AOI21xp5_ASAP7_75t_L g5361 ( 
.A1(n_4933),
.A2(n_2546),
.B(n_2542),
.Y(n_5361)
);

OAI21x1_ASAP7_75t_L g5362 ( 
.A1(n_4673),
.A2(n_3215),
.B(n_3211),
.Y(n_5362)
);

OAI22xp5_ASAP7_75t_L g5363 ( 
.A1(n_4837),
.A2(n_4700),
.B1(n_4817),
.B2(n_4936),
.Y(n_5363)
);

HB1xp67_ASAP7_75t_L g5364 ( 
.A(n_4891),
.Y(n_5364)
);

OA21x2_ASAP7_75t_L g5365 ( 
.A1(n_4894),
.A2(n_1550),
.B(n_1543),
.Y(n_5365)
);

BUFx2_ASAP7_75t_L g5366 ( 
.A(n_4950),
.Y(n_5366)
);

AO31x2_ASAP7_75t_L g5367 ( 
.A1(n_4726),
.A2(n_3218),
.A3(n_3229),
.B(n_3215),
.Y(n_5367)
);

AND2x2_ASAP7_75t_L g5368 ( 
.A(n_4786),
.B(n_11),
.Y(n_5368)
);

AO31x2_ASAP7_75t_L g5369 ( 
.A1(n_4751),
.A2(n_3229),
.A3(n_3232),
.B(n_3218),
.Y(n_5369)
);

AOI22xp33_ASAP7_75t_L g5370 ( 
.A1(n_4974),
.A2(n_3283),
.B1(n_3288),
.B2(n_3278),
.Y(n_5370)
);

AOI21xp5_ASAP7_75t_L g5371 ( 
.A1(n_4843),
.A2(n_2547),
.B(n_2546),
.Y(n_5371)
);

OAI221xp5_ASAP7_75t_L g5372 ( 
.A1(n_4765),
.A2(n_1020),
.B1(n_1021),
.B2(n_1018),
.C(n_1015),
.Y(n_5372)
);

OAI21x1_ASAP7_75t_L g5373 ( 
.A1(n_4678),
.A2(n_4647),
.B(n_4947),
.Y(n_5373)
);

AOI21xp33_ASAP7_75t_L g5374 ( 
.A1(n_4883),
.A2(n_1027),
.B(n_1025),
.Y(n_5374)
);

INVx2_ASAP7_75t_L g5375 ( 
.A(n_4808),
.Y(n_5375)
);

O2A1O1Ixp33_ASAP7_75t_L g5376 ( 
.A1(n_4765),
.A2(n_2305),
.B(n_2196),
.C(n_2197),
.Y(n_5376)
);

NAND2xp5_ASAP7_75t_SL g5377 ( 
.A(n_4863),
.B(n_2286),
.Y(n_5377)
);

OAI21x1_ASAP7_75t_L g5378 ( 
.A1(n_4678),
.A2(n_3241),
.B(n_3232),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_4754),
.Y(n_5379)
);

OAI21x1_ASAP7_75t_L g5380 ( 
.A1(n_4647),
.A2(n_3244),
.B(n_3241),
.Y(n_5380)
);

INVx3_ASAP7_75t_L g5381 ( 
.A(n_4955),
.Y(n_5381)
);

AOI221x1_ASAP7_75t_L g5382 ( 
.A1(n_4959),
.A2(n_4831),
.B1(n_4836),
.B2(n_4846),
.C(n_4969),
.Y(n_5382)
);

CKINVDCx20_ASAP7_75t_R g5383 ( 
.A(n_4763),
.Y(n_5383)
);

AOI21xp5_ASAP7_75t_L g5384 ( 
.A1(n_4951),
.A2(n_2557),
.B(n_2547),
.Y(n_5384)
);

AND2x2_ASAP7_75t_L g5385 ( 
.A(n_4811),
.B(n_11),
.Y(n_5385)
);

NAND2xp33_ASAP7_75t_L g5386 ( 
.A(n_4643),
.B(n_1032),
.Y(n_5386)
);

OAI22xp5_ASAP7_75t_L g5387 ( 
.A1(n_4837),
.A2(n_1040),
.B1(n_1044),
.B2(n_1034),
.Y(n_5387)
);

OAI21x1_ASAP7_75t_L g5388 ( 
.A1(n_5038),
.A2(n_4969),
.B(n_4591),
.Y(n_5388)
);

OAI21x1_ASAP7_75t_L g5389 ( 
.A1(n_5130),
.A2(n_5143),
.B(n_5170),
.Y(n_5389)
);

BUFx6f_ASAP7_75t_L g5390 ( 
.A(n_5008),
.Y(n_5390)
);

AOI221xp5_ASAP7_75t_L g5391 ( 
.A1(n_5210),
.A2(n_5089),
.B1(n_5019),
.B2(n_4993),
.C(n_5271),
.Y(n_5391)
);

AOI22xp33_ASAP7_75t_L g5392 ( 
.A1(n_5147),
.A2(n_5249),
.B1(n_5089),
.B2(n_5019),
.Y(n_5392)
);

BUFx10_ASAP7_75t_L g5393 ( 
.A(n_5265),
.Y(n_5393)
);

AND2x6_ASAP7_75t_L g5394 ( 
.A(n_5238),
.B(n_4676),
.Y(n_5394)
);

NOR2xp33_ASAP7_75t_L g5395 ( 
.A(n_5195),
.B(n_4976),
.Y(n_5395)
);

INVx2_ASAP7_75t_L g5396 ( 
.A(n_5274),
.Y(n_5396)
);

HB1xp67_ASAP7_75t_L g5397 ( 
.A(n_5110),
.Y(n_5397)
);

AOI22x1_ASAP7_75t_L g5398 ( 
.A1(n_5043),
.A2(n_4916),
.B1(n_4888),
.B2(n_4955),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5289),
.Y(n_5399)
);

OAI221xp5_ASAP7_75t_L g5400 ( 
.A1(n_5271),
.A2(n_4922),
.B1(n_4965),
.B2(n_4890),
.C(n_4939),
.Y(n_5400)
);

INVx4_ASAP7_75t_L g5401 ( 
.A(n_5043),
.Y(n_5401)
);

HB1xp67_ASAP7_75t_L g5402 ( 
.A(n_5165),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_5289),
.Y(n_5403)
);

NOR2xp67_ASAP7_75t_L g5404 ( 
.A(n_5008),
.B(n_5187),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5289),
.Y(n_5405)
);

INVxp67_ASAP7_75t_L g5406 ( 
.A(n_5263),
.Y(n_5406)
);

BUFx6f_ASAP7_75t_L g5407 ( 
.A(n_5008),
.Y(n_5407)
);

CKINVDCx5p33_ASAP7_75t_R g5408 ( 
.A(n_4998),
.Y(n_5408)
);

BUFx10_ASAP7_75t_L g5409 ( 
.A(n_5058),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_4995),
.Y(n_5410)
);

INVx4_ASAP7_75t_L g5411 ( 
.A(n_5027),
.Y(n_5411)
);

OAI21x1_ASAP7_75t_L g5412 ( 
.A1(n_5175),
.A2(n_4985),
.B(n_5279),
.Y(n_5412)
);

AOI22xp33_ASAP7_75t_SL g5413 ( 
.A1(n_5047),
.A2(n_4643),
.B1(n_4943),
.B2(n_4676),
.Y(n_5413)
);

INVx3_ASAP7_75t_L g5414 ( 
.A(n_5187),
.Y(n_5414)
);

OAI22xp33_ASAP7_75t_L g5415 ( 
.A1(n_5014),
.A2(n_4598),
.B1(n_4646),
.B2(n_4873),
.Y(n_5415)
);

A2O1A1Ixp33_ASAP7_75t_L g5416 ( 
.A1(n_5254),
.A2(n_4890),
.B(n_4922),
.C(n_4957),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5274),
.Y(n_5417)
);

BUFx2_ASAP7_75t_L g5418 ( 
.A(n_5326),
.Y(n_5418)
);

AOI221xp5_ASAP7_75t_L g5419 ( 
.A1(n_4993),
.A2(n_1053),
.B1(n_1058),
.B2(n_1048),
.C(n_1045),
.Y(n_5419)
);

AND2x2_ASAP7_75t_L g5420 ( 
.A(n_5117),
.B(n_4811),
.Y(n_5420)
);

NAND3xp33_ASAP7_75t_L g5421 ( 
.A(n_5348),
.B(n_5382),
.C(n_5233),
.Y(n_5421)
);

CKINVDCx20_ASAP7_75t_R g5422 ( 
.A(n_5225),
.Y(n_5422)
);

OAI21xp33_ASAP7_75t_SL g5423 ( 
.A1(n_5029),
.A2(n_5097),
.B(n_5076),
.Y(n_5423)
);

INVx2_ASAP7_75t_SL g5424 ( 
.A(n_5067),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5016),
.Y(n_5425)
);

OAI21x1_ASAP7_75t_L g5426 ( 
.A1(n_5201),
.A2(n_4591),
.B(n_4948),
.Y(n_5426)
);

INVx1_ASAP7_75t_SL g5427 ( 
.A(n_5157),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_5243),
.B(n_4770),
.Y(n_5428)
);

BUFx2_ASAP7_75t_L g5429 ( 
.A(n_5350),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5044),
.Y(n_5430)
);

NOR2xp33_ASAP7_75t_L g5431 ( 
.A(n_5135),
.B(n_4888),
.Y(n_5431)
);

CKINVDCx6p67_ASAP7_75t_R g5432 ( 
.A(n_5304),
.Y(n_5432)
);

OAI21x1_ASAP7_75t_L g5433 ( 
.A1(n_5007),
.A2(n_4820),
.B(n_4829),
.Y(n_5433)
);

AOI21xp5_ASAP7_75t_L g5434 ( 
.A1(n_5127),
.A2(n_4725),
.B(n_4970),
.Y(n_5434)
);

OA21x2_ASAP7_75t_L g5435 ( 
.A1(n_5138),
.A2(n_4796),
.B(n_4732),
.Y(n_5435)
);

OAI21xp5_ASAP7_75t_L g5436 ( 
.A1(n_5023),
.A2(n_4957),
.B(n_4939),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5224),
.B(n_4820),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_5062),
.Y(n_5438)
);

INVx3_ASAP7_75t_L g5439 ( 
.A(n_5224),
.Y(n_5439)
);

OA21x2_ASAP7_75t_L g5440 ( 
.A1(n_5317),
.A2(n_4731),
.B(n_4810),
.Y(n_5440)
);

OAI21x1_ASAP7_75t_L g5441 ( 
.A1(n_4997),
.A2(n_4870),
.B(n_4827),
.Y(n_5441)
);

AND2x4_ASAP7_75t_L g5442 ( 
.A(n_5238),
.B(n_4870),
.Y(n_5442)
);

HB1xp67_ASAP7_75t_L g5443 ( 
.A(n_5083),
.Y(n_5443)
);

AO21x2_ASAP7_75t_L g5444 ( 
.A1(n_5317),
.A2(n_4825),
.B(n_4773),
.Y(n_5444)
);

OAI21x1_ASAP7_75t_L g5445 ( 
.A1(n_4990),
.A2(n_4769),
.B(n_4929),
.Y(n_5445)
);

AO21x2_ASAP7_75t_L g5446 ( 
.A1(n_5109),
.A2(n_4776),
.B(n_4772),
.Y(n_5446)
);

OAI21x1_ASAP7_75t_L g5447 ( 
.A1(n_5250),
.A2(n_4929),
.B(n_4980),
.Y(n_5447)
);

OAI21xp5_ASAP7_75t_L g5448 ( 
.A1(n_5128),
.A2(n_4722),
.B(n_4916),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5066),
.Y(n_5449)
);

AND2x2_ASAP7_75t_L g5450 ( 
.A(n_5029),
.B(n_4779),
.Y(n_5450)
);

CKINVDCx11_ASAP7_75t_R g5451 ( 
.A(n_5025),
.Y(n_5451)
);

AND2x2_ASAP7_75t_L g5452 ( 
.A(n_5097),
.B(n_4787),
.Y(n_5452)
);

INVx1_ASAP7_75t_SL g5453 ( 
.A(n_5296),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_5278),
.Y(n_5454)
);

AND2x2_ASAP7_75t_L g5455 ( 
.A(n_5011),
.B(n_4802),
.Y(n_5455)
);

AOI221xp5_ASAP7_75t_L g5456 ( 
.A1(n_5000),
.A2(n_1065),
.B1(n_1067),
.B2(n_1062),
.C(n_1061),
.Y(n_5456)
);

AND2x2_ASAP7_75t_L g5457 ( 
.A(n_5001),
.B(n_4804),
.Y(n_5457)
);

OA21x2_ASAP7_75t_L g5458 ( 
.A1(n_5234),
.A2(n_4823),
.B(n_4818),
.Y(n_5458)
);

INVx3_ASAP7_75t_L g5459 ( 
.A(n_5248),
.Y(n_5459)
);

OAI221xp5_ASAP7_75t_L g5460 ( 
.A1(n_5098),
.A2(n_1074),
.B1(n_1079),
.B2(n_1073),
.C(n_1071),
.Y(n_5460)
);

NAND2xp33_ASAP7_75t_L g5461 ( 
.A(n_5299),
.B(n_4643),
.Y(n_5461)
);

OR2x2_ASAP7_75t_L g5462 ( 
.A(n_5078),
.B(n_4824),
.Y(n_5462)
);

NOR2xp33_ASAP7_75t_L g5463 ( 
.A(n_5220),
.B(n_4934),
.Y(n_5463)
);

INVx2_ASAP7_75t_L g5464 ( 
.A(n_5274),
.Y(n_5464)
);

INVx2_ASAP7_75t_L g5465 ( 
.A(n_5333),
.Y(n_5465)
);

OAI21x1_ASAP7_75t_L g5466 ( 
.A1(n_4989),
.A2(n_4828),
.B(n_4761),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_5280),
.Y(n_5467)
);

OAI21x1_ASAP7_75t_L g5468 ( 
.A1(n_4992),
.A2(n_4774),
.B(n_4755),
.Y(n_5468)
);

OA21x2_ASAP7_75t_L g5469 ( 
.A1(n_5244),
.A2(n_4784),
.B(n_4775),
.Y(n_5469)
);

AOI22x1_ASAP7_75t_L g5470 ( 
.A1(n_5184),
.A2(n_4928),
.B1(n_1087),
.B2(n_1089),
.Y(n_5470)
);

AOI22xp5_ASAP7_75t_L g5471 ( 
.A1(n_5193),
.A2(n_4863),
.B1(n_4905),
.B2(n_4865),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5281),
.Y(n_5472)
);

OAI21x1_ASAP7_75t_L g5473 ( 
.A1(n_5074),
.A2(n_4790),
.B(n_4725),
.Y(n_5473)
);

AND2x4_ASAP7_75t_L g5474 ( 
.A(n_4982),
.B(n_4598),
.Y(n_5474)
);

NAND3xp33_ASAP7_75t_L g5475 ( 
.A(n_5364),
.B(n_4977),
.C(n_4905),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_5082),
.B(n_4977),
.Y(n_5476)
);

OAI21x1_ASAP7_75t_L g5477 ( 
.A1(n_5077),
.A2(n_4725),
.B(n_2200),
.Y(n_5477)
);

OAI21x1_ASAP7_75t_L g5478 ( 
.A1(n_5012),
.A2(n_2200),
.B(n_2192),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5353),
.Y(n_5479)
);

OR2x2_ASAP7_75t_L g5480 ( 
.A(n_5084),
.B(n_4767),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5354),
.Y(n_5481)
);

OAI21x1_ASAP7_75t_L g5482 ( 
.A1(n_5121),
.A2(n_2201),
.B(n_2192),
.Y(n_5482)
);

INVx5_ASAP7_75t_SL g5483 ( 
.A(n_5079),
.Y(n_5483)
);

NAND2xp5_ASAP7_75t_L g5484 ( 
.A(n_5283),
.B(n_4977),
.Y(n_5484)
);

INVx3_ASAP7_75t_L g5485 ( 
.A(n_5248),
.Y(n_5485)
);

OA21x2_ASAP7_75t_L g5486 ( 
.A1(n_5373),
.A2(n_4974),
.B(n_4822),
.Y(n_5486)
);

NAND2xp5_ASAP7_75t_L g5487 ( 
.A(n_5298),
.B(n_4977),
.Y(n_5487)
);

OAI21xp5_ASAP7_75t_L g5488 ( 
.A1(n_5128),
.A2(n_4822),
.B(n_1091),
.Y(n_5488)
);

NAND2xp5_ASAP7_75t_L g5489 ( 
.A(n_5086),
.B(n_4912),
.Y(n_5489)
);

AND2x2_ASAP7_75t_L g5490 ( 
.A(n_5051),
.B(n_4767),
.Y(n_5490)
);

INVx6_ASAP7_75t_L g5491 ( 
.A(n_5092),
.Y(n_5491)
);

OAI21x1_ASAP7_75t_L g5492 ( 
.A1(n_5010),
.A2(n_2203),
.B(n_2201),
.Y(n_5492)
);

OAI21x1_ASAP7_75t_L g5493 ( 
.A1(n_5030),
.A2(n_2207),
.B(n_2203),
.Y(n_5493)
);

NAND2xp5_ASAP7_75t_L g5494 ( 
.A(n_5264),
.B(n_4912),
.Y(n_5494)
);

OAI21x1_ASAP7_75t_L g5495 ( 
.A1(n_5031),
.A2(n_2216),
.B(n_2207),
.Y(n_5495)
);

OAI21x1_ASAP7_75t_L g5496 ( 
.A1(n_5013),
.A2(n_2216),
.B(n_4598),
.Y(n_5496)
);

BUFx6f_ASAP7_75t_L g5497 ( 
.A(n_5327),
.Y(n_5497)
);

INVx2_ASAP7_75t_L g5498 ( 
.A(n_5177),
.Y(n_5498)
);

OAI22xp5_ASAP7_75t_L g5499 ( 
.A1(n_5193),
.A2(n_4646),
.B1(n_4905),
.B2(n_4865),
.Y(n_5499)
);

OAI21x1_ASAP7_75t_L g5500 ( 
.A1(n_5015),
.A2(n_4646),
.B(n_3250),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5093),
.B(n_4912),
.Y(n_5501)
);

OAI21x1_ASAP7_75t_L g5502 ( 
.A1(n_5063),
.A2(n_4646),
.B(n_3250),
.Y(n_5502)
);

OAI21x1_ASAP7_75t_L g5503 ( 
.A1(n_5064),
.A2(n_3252),
.B(n_3244),
.Y(n_5503)
);

INVx1_ASAP7_75t_L g5504 ( 
.A(n_5177),
.Y(n_5504)
);

OAI21x1_ASAP7_75t_SL g5505 ( 
.A1(n_5313),
.A2(n_4633),
.B(n_4912),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_5177),
.Y(n_5506)
);

NAND2xp5_ASAP7_75t_L g5507 ( 
.A(n_5379),
.B(n_4934),
.Y(n_5507)
);

OR2x6_ASAP7_75t_L g5508 ( 
.A(n_5053),
.B(n_4778),
.Y(n_5508)
);

OA21x2_ASAP7_75t_L g5509 ( 
.A1(n_5109),
.A2(n_4801),
.B(n_4794),
.Y(n_5509)
);

AO21x2_ASAP7_75t_L g5510 ( 
.A1(n_5116),
.A2(n_4801),
.B(n_4794),
.Y(n_5510)
);

OAI21x1_ASAP7_75t_L g5511 ( 
.A1(n_5020),
.A2(n_3256),
.B(n_3252),
.Y(n_5511)
);

AND2x2_ASAP7_75t_L g5512 ( 
.A(n_5217),
.B(n_4767),
.Y(n_5512)
);

OAI21x1_ASAP7_75t_L g5513 ( 
.A1(n_5021),
.A2(n_5004),
.B(n_5091),
.Y(n_5513)
);

CKINVDCx5p33_ASAP7_75t_R g5514 ( 
.A(n_5094),
.Y(n_5514)
);

NOR2xp33_ASAP7_75t_L g5515 ( 
.A(n_5220),
.B(n_4934),
.Y(n_5515)
);

BUFx10_ASAP7_75t_L g5516 ( 
.A(n_5202),
.Y(n_5516)
);

OAI21xp5_ASAP7_75t_L g5517 ( 
.A1(n_5026),
.A2(n_1094),
.B(n_1083),
.Y(n_5517)
);

AND2x4_ASAP7_75t_L g5518 ( 
.A(n_4982),
.B(n_4767),
.Y(n_5518)
);

AND2x6_ASAP7_75t_L g5519 ( 
.A(n_5151),
.B(n_4653),
.Y(n_5519)
);

OAI21x1_ASAP7_75t_L g5520 ( 
.A1(n_5134),
.A2(n_3263),
.B(n_3256),
.Y(n_5520)
);

CKINVDCx5p33_ASAP7_75t_R g5521 ( 
.A(n_5261),
.Y(n_5521)
);

INVx3_ASAP7_75t_L g5522 ( 
.A(n_5381),
.Y(n_5522)
);

NAND2xp5_ASAP7_75t_L g5523 ( 
.A(n_5174),
.B(n_4934),
.Y(n_5523)
);

AOI22xp33_ASAP7_75t_SL g5524 ( 
.A1(n_5057),
.A2(n_4905),
.B1(n_4865),
.B2(n_4863),
.Y(n_5524)
);

OA21x2_ASAP7_75t_L g5525 ( 
.A1(n_5116),
.A2(n_4809),
.B(n_1550),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_5163),
.Y(n_5526)
);

OAI21x1_ASAP7_75t_L g5527 ( 
.A1(n_5156),
.A2(n_3266),
.B(n_3263),
.Y(n_5527)
);

OAI21x1_ASAP7_75t_L g5528 ( 
.A1(n_5033),
.A2(n_3278),
.B(n_3266),
.Y(n_5528)
);

OAI21x1_ASAP7_75t_L g5529 ( 
.A1(n_5159),
.A2(n_3288),
.B(n_3283),
.Y(n_5529)
);

INVx2_ASAP7_75t_L g5530 ( 
.A(n_5247),
.Y(n_5530)
);

AOI22xp33_ASAP7_75t_L g5531 ( 
.A1(n_5147),
.A2(n_2287),
.B1(n_2286),
.B2(n_4809),
.Y(n_5531)
);

INVx2_ASAP7_75t_L g5532 ( 
.A(n_5296),
.Y(n_5532)
);

OAI21x1_ASAP7_75t_L g5533 ( 
.A1(n_5006),
.A2(n_5100),
.B(n_5221),
.Y(n_5533)
);

OA21x2_ASAP7_75t_L g5534 ( 
.A1(n_5259),
.A2(n_1575),
.B(n_1543),
.Y(n_5534)
);

OAI21x1_ASAP7_75t_L g5535 ( 
.A1(n_5040),
.A2(n_3303),
.B(n_3302),
.Y(n_5535)
);

OAI21x1_ASAP7_75t_L g5536 ( 
.A1(n_5252),
.A2(n_3303),
.B(n_3302),
.Y(n_5536)
);

BUFx2_ASAP7_75t_L g5537 ( 
.A(n_5366),
.Y(n_5537)
);

INVx4_ASAP7_75t_L g5538 ( 
.A(n_5164),
.Y(n_5538)
);

INVx2_ASAP7_75t_L g5539 ( 
.A(n_5258),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_5240),
.Y(n_5540)
);

AND2x2_ASAP7_75t_L g5541 ( 
.A(n_5048),
.B(n_4616),
.Y(n_5541)
);

OAI21x1_ASAP7_75t_L g5542 ( 
.A1(n_5160),
.A2(n_2562),
.B(n_2557),
.Y(n_5542)
);

AO21x2_ASAP7_75t_L g5543 ( 
.A1(n_5269),
.A2(n_1590),
.B(n_1575),
.Y(n_5543)
);

NOR2xp33_ASAP7_75t_L g5544 ( 
.A(n_5050),
.B(n_4940),
.Y(n_5544)
);

AND2x2_ASAP7_75t_L g5545 ( 
.A(n_5048),
.B(n_4616),
.Y(n_5545)
);

OR2x2_ASAP7_75t_L g5546 ( 
.A(n_5131),
.B(n_4653),
.Y(n_5546)
);

HB1xp67_ASAP7_75t_L g5547 ( 
.A(n_5099),
.Y(n_5547)
);

INVx2_ASAP7_75t_SL g5548 ( 
.A(n_5125),
.Y(n_5548)
);

OAI21x1_ASAP7_75t_L g5549 ( 
.A1(n_5162),
.A2(n_2569),
.B(n_2562),
.Y(n_5549)
);

NAND2x1p5_ASAP7_75t_L g5550 ( 
.A(n_5151),
.B(n_4616),
.Y(n_5550)
);

NAND2xp5_ASAP7_75t_L g5551 ( 
.A(n_5088),
.B(n_5036),
.Y(n_5551)
);

A2O1A1Ixp33_ASAP7_75t_L g5552 ( 
.A1(n_5254),
.A2(n_4745),
.B(n_4863),
.C(n_4865),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5255),
.Y(n_5553)
);

NOR2xp33_ASAP7_75t_L g5554 ( 
.A(n_5087),
.B(n_4940),
.Y(n_5554)
);

OAI21xp5_ASAP7_75t_L g5555 ( 
.A1(n_5246),
.A2(n_1098),
.B(n_1097),
.Y(n_5555)
);

INVx3_ASAP7_75t_L g5556 ( 
.A(n_5381),
.Y(n_5556)
);

OAI22xp5_ASAP7_75t_L g5557 ( 
.A1(n_5144),
.A2(n_4941),
.B1(n_4942),
.B2(n_4940),
.Y(n_5557)
);

O2A1O1Ixp33_ASAP7_75t_SL g5558 ( 
.A1(n_5325),
.A2(n_160),
.B(n_161),
.C(n_159),
.Y(n_5558)
);

OAI21x1_ASAP7_75t_L g5559 ( 
.A1(n_5039),
.A2(n_2575),
.B(n_2569),
.Y(n_5559)
);

OAI21x1_ASAP7_75t_SL g5560 ( 
.A1(n_5028),
.A2(n_4941),
.B(n_4940),
.Y(n_5560)
);

INVxp67_ASAP7_75t_L g5561 ( 
.A(n_4996),
.Y(n_5561)
);

BUFx3_ASAP7_75t_L g5562 ( 
.A(n_5092),
.Y(n_5562)
);

OAI21x1_ASAP7_75t_L g5563 ( 
.A1(n_5229),
.A2(n_5262),
.B(n_5259),
.Y(n_5563)
);

BUFx2_ASAP7_75t_L g5564 ( 
.A(n_5383),
.Y(n_5564)
);

A2O1A1Ixp33_ASAP7_75t_L g5565 ( 
.A1(n_5144),
.A2(n_1100),
.B(n_1109),
.C(n_1099),
.Y(n_5565)
);

OA21x2_ASAP7_75t_L g5566 ( 
.A1(n_5262),
.A2(n_1607),
.B(n_1590),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_5308),
.Y(n_5567)
);

OAI21x1_ASAP7_75t_L g5568 ( 
.A1(n_5229),
.A2(n_2579),
.B(n_2575),
.Y(n_5568)
);

AOI21x1_ASAP7_75t_L g5569 ( 
.A1(n_5065),
.A2(n_1611),
.B(n_1607),
.Y(n_5569)
);

INVx2_ASAP7_75t_L g5570 ( 
.A(n_5200),
.Y(n_5570)
);

INVx5_ASAP7_75t_L g5571 ( 
.A(n_5151),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_5255),
.Y(n_5572)
);

HB1xp67_ASAP7_75t_L g5573 ( 
.A(n_5101),
.Y(n_5573)
);

AOI21xp5_ASAP7_75t_L g5574 ( 
.A1(n_5127),
.A2(n_4942),
.B(n_4941),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5169),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_5197),
.Y(n_5576)
);

INVx3_ASAP7_75t_L g5577 ( 
.A(n_5102),
.Y(n_5577)
);

OAI21x1_ASAP7_75t_SL g5578 ( 
.A1(n_5028),
.A2(n_4942),
.B(n_4941),
.Y(n_5578)
);

AOI21xp5_ASAP7_75t_L g5579 ( 
.A1(n_5371),
.A2(n_5185),
.B(n_5270),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5176),
.Y(n_5580)
);

OAI22xp5_ASAP7_75t_L g5581 ( 
.A1(n_5249),
.A2(n_4956),
.B1(n_4971),
.B2(n_4942),
.Y(n_5581)
);

NAND2x1p5_ASAP7_75t_L g5582 ( 
.A(n_5053),
.B(n_4617),
.Y(n_5582)
);

O2A1O1Ixp33_ASAP7_75t_SL g5583 ( 
.A1(n_5018),
.A2(n_162),
.B(n_163),
.C(n_160),
.Y(n_5583)
);

OR2x6_ASAP7_75t_L g5584 ( 
.A(n_5115),
.B(n_4617),
.Y(n_5584)
);

INVxp67_ASAP7_75t_SL g5585 ( 
.A(n_4987),
.Y(n_5585)
);

OR2x2_ASAP7_75t_L g5586 ( 
.A(n_5186),
.B(n_4670),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5226),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_L g5588 ( 
.A(n_5032),
.B(n_4956),
.Y(n_5588)
);

BUFx10_ASAP7_75t_L g5589 ( 
.A(n_5129),
.Y(n_5589)
);

INVx2_ASAP7_75t_L g5590 ( 
.A(n_5203),
.Y(n_5590)
);

AOI22xp33_ASAP7_75t_SL g5591 ( 
.A1(n_5057),
.A2(n_5318),
.B1(n_4999),
.B2(n_5363),
.Y(n_5591)
);

OAI21x1_ASAP7_75t_L g5592 ( 
.A1(n_5223),
.A2(n_2579),
.B(n_4956),
.Y(n_5592)
);

INVx3_ASAP7_75t_L g5593 ( 
.A(n_5102),
.Y(n_5593)
);

NAND2x1p5_ASAP7_75t_L g5594 ( 
.A(n_5115),
.B(n_4617),
.Y(n_5594)
);

NAND2x1p5_ASAP7_75t_L g5595 ( 
.A(n_5009),
.B(n_4617),
.Y(n_5595)
);

BUFx6f_ASAP7_75t_L g5596 ( 
.A(n_5327),
.Y(n_5596)
);

INVx2_ASAP7_75t_L g5597 ( 
.A(n_5002),
.Y(n_5597)
);

BUFx2_ASAP7_75t_SL g5598 ( 
.A(n_5312),
.Y(n_5598)
);

OAI21xp5_ASAP7_75t_L g5599 ( 
.A1(n_5246),
.A2(n_5266),
.B(n_5000),
.Y(n_5599)
);

OAI22xp5_ASAP7_75t_L g5600 ( 
.A1(n_5168),
.A2(n_4971),
.B1(n_4956),
.B2(n_4708),
.Y(n_5600)
);

AOI21xp33_ASAP7_75t_L g5601 ( 
.A1(n_5122),
.A2(n_4971),
.B(n_4851),
.Y(n_5601)
);

NAND3xp33_ASAP7_75t_SL g5602 ( 
.A(n_5035),
.B(n_1112),
.C(n_1111),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5237),
.Y(n_5603)
);

INVx2_ASAP7_75t_L g5604 ( 
.A(n_5022),
.Y(n_5604)
);

BUFx6f_ASAP7_75t_L g5605 ( 
.A(n_5334),
.Y(n_5605)
);

INVxp33_ASAP7_75t_SL g5606 ( 
.A(n_5241),
.Y(n_5606)
);

INVx5_ASAP7_75t_L g5607 ( 
.A(n_5318),
.Y(n_5607)
);

AOI221xp5_ASAP7_75t_L g5608 ( 
.A1(n_5005),
.A2(n_1126),
.B1(n_1127),
.B2(n_1115),
.C(n_1113),
.Y(n_5608)
);

AOI22xp33_ASAP7_75t_L g5609 ( 
.A1(n_5090),
.A2(n_2287),
.B1(n_2286),
.B2(n_2186),
.Y(n_5609)
);

OAI21x1_ASAP7_75t_L g5610 ( 
.A1(n_5231),
.A2(n_4971),
.B(n_4851),
.Y(n_5610)
);

OA21x2_ASAP7_75t_L g5611 ( 
.A1(n_5191),
.A2(n_1618),
.B(n_1611),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5055),
.Y(n_5612)
);

NAND2x1p5_ASAP7_75t_L g5613 ( 
.A(n_5009),
.B(n_5137),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5114),
.Y(n_5614)
);

OAI21x1_ASAP7_75t_L g5615 ( 
.A1(n_5303),
.A2(n_4851),
.B(n_1639),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5136),
.Y(n_5616)
);

BUFx2_ASAP7_75t_L g5617 ( 
.A(n_5104),
.Y(n_5617)
);

INVx2_ASAP7_75t_SL g5618 ( 
.A(n_5267),
.Y(n_5618)
);

NAND2xp5_ASAP7_75t_L g5619 ( 
.A(n_5071),
.B(n_4851),
.Y(n_5619)
);

NAND2x1p5_ASAP7_75t_L g5620 ( 
.A(n_5137),
.B(n_4640),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_4988),
.A2(n_4708),
.B(n_4670),
.Y(n_5621)
);

OAI22xp5_ASAP7_75t_L g5622 ( 
.A1(n_5168),
.A2(n_4708),
.B1(n_4670),
.B2(n_4642),
.Y(n_5622)
);

OAI21x1_ASAP7_75t_L g5623 ( 
.A1(n_5303),
.A2(n_1639),
.B(n_1618),
.Y(n_5623)
);

OAI21x1_ASAP7_75t_L g5624 ( 
.A1(n_5042),
.A2(n_1654),
.B(n_1641),
.Y(n_5624)
);

BUFx3_ASAP7_75t_L g5625 ( 
.A(n_5222),
.Y(n_5625)
);

BUFx2_ASAP7_75t_L g5626 ( 
.A(n_5104),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5347),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5103),
.Y(n_5628)
);

CKINVDCx20_ASAP7_75t_R g5629 ( 
.A(n_5309),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_5191),
.Y(n_5630)
);

BUFx3_ASAP7_75t_L g5631 ( 
.A(n_5344),
.Y(n_5631)
);

AND2x4_ASAP7_75t_L g5632 ( 
.A(n_4994),
.B(n_4640),
.Y(n_5632)
);

NAND3xp33_ASAP7_75t_L g5633 ( 
.A(n_5340),
.B(n_4642),
.C(n_4640),
.Y(n_5633)
);

CKINVDCx20_ASAP7_75t_R g5634 ( 
.A(n_4991),
.Y(n_5634)
);

AOI211x1_ASAP7_75t_L g5635 ( 
.A1(n_5276),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_5635)
);

AOI22xp33_ASAP7_75t_L g5636 ( 
.A1(n_5199),
.A2(n_2287),
.B1(n_2186),
.B2(n_2193),
.Y(n_5636)
);

OAI21x1_ASAP7_75t_L g5637 ( 
.A1(n_5365),
.A2(n_1654),
.B(n_1641),
.Y(n_5637)
);

INVx6_ASAP7_75t_L g5638 ( 
.A(n_5111),
.Y(n_5638)
);

INVxp67_ASAP7_75t_SL g5639 ( 
.A(n_5178),
.Y(n_5639)
);

AND2x4_ASAP7_75t_L g5640 ( 
.A(n_5171),
.B(n_4640),
.Y(n_5640)
);

INVx2_ASAP7_75t_SL g5641 ( 
.A(n_5310),
.Y(n_5641)
);

HB1xp67_ASAP7_75t_L g5642 ( 
.A(n_5285),
.Y(n_5642)
);

AOI21x1_ASAP7_75t_L g5643 ( 
.A1(n_5072),
.A2(n_1664),
.B(n_1659),
.Y(n_5643)
);

AO31x2_ASAP7_75t_L g5644 ( 
.A1(n_5204),
.A2(n_1664),
.A3(n_1675),
.B(n_1659),
.Y(n_5644)
);

AND2x4_ASAP7_75t_L g5645 ( 
.A(n_5171),
.B(n_4642),
.Y(n_5645)
);

CKINVDCx5p33_ASAP7_75t_R g5646 ( 
.A(n_5196),
.Y(n_5646)
);

OAI21x1_ASAP7_75t_L g5647 ( 
.A1(n_5365),
.A2(n_1675),
.B(n_2582),
.Y(n_5647)
);

NAND2xp5_ASAP7_75t_L g5648 ( 
.A(n_5285),
.B(n_4642),
.Y(n_5648)
);

AND2x2_ASAP7_75t_L g5649 ( 
.A(n_5209),
.B(n_4670),
.Y(n_5649)
);

NAND2xp5_ASAP7_75t_L g5650 ( 
.A(n_5081),
.B(n_4708),
.Y(n_5650)
);

BUFx8_ASAP7_75t_SL g5651 ( 
.A(n_5111),
.Y(n_5651)
);

NAND2xp33_ASAP7_75t_R g5652 ( 
.A(n_5341),
.B(n_164),
.Y(n_5652)
);

HB1xp67_ASAP7_75t_L g5653 ( 
.A(n_5052),
.Y(n_5653)
);

AND2x2_ASAP7_75t_L g5654 ( 
.A(n_5209),
.B(n_12),
.Y(n_5654)
);

AO21x2_ASAP7_75t_L g5655 ( 
.A1(n_5324),
.A2(n_1351),
.B(n_1348),
.Y(n_5655)
);

AND2x2_ASAP7_75t_L g5656 ( 
.A(n_5141),
.B(n_12),
.Y(n_5656)
);

O2A1O1Ixp33_ASAP7_75t_L g5657 ( 
.A1(n_5346),
.A2(n_2306),
.B(n_2298),
.C(n_15),
.Y(n_5657)
);

A2O1A1Ixp33_ASAP7_75t_L g5658 ( 
.A1(n_5386),
.A2(n_1135),
.B(n_1138),
.C(n_1129),
.Y(n_5658)
);

HB1xp67_ASAP7_75t_L g5659 ( 
.A(n_5052),
.Y(n_5659)
);

AOI22xp33_ASAP7_75t_L g5660 ( 
.A1(n_5199),
.A2(n_2287),
.B1(n_2186),
.B2(n_2193),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_5343),
.Y(n_5661)
);

OAI21x1_ASAP7_75t_L g5662 ( 
.A1(n_5288),
.A2(n_2588),
.B(n_2582),
.Y(n_5662)
);

AOI22xp5_ASAP7_75t_L g5663 ( 
.A1(n_5266),
.A2(n_5363),
.B1(n_5294),
.B2(n_5228),
.Y(n_5663)
);

INVx2_ASAP7_75t_SL g5664 ( 
.A(n_5111),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5345),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5375),
.Y(n_5666)
);

HB1xp67_ASAP7_75t_L g5667 ( 
.A(n_5052),
.Y(n_5667)
);

OR2x6_ASAP7_75t_L g5668 ( 
.A(n_5148),
.B(n_3031),
.Y(n_5668)
);

OAI21x1_ASAP7_75t_L g5669 ( 
.A1(n_5218),
.A2(n_2589),
.B(n_2588),
.Y(n_5669)
);

OAI21x1_ASAP7_75t_L g5670 ( 
.A1(n_4983),
.A2(n_2592),
.B(n_2589),
.Y(n_5670)
);

BUFx3_ASAP7_75t_L g5671 ( 
.A(n_5260),
.Y(n_5671)
);

OAI22xp33_ASAP7_75t_L g5672 ( 
.A1(n_5054),
.A2(n_1143),
.B1(n_1144),
.B2(n_1142),
.Y(n_5672)
);

NAND2x1_ASAP7_75t_L g5673 ( 
.A(n_5329),
.B(n_3031),
.Y(n_5673)
);

AOI22xp33_ASAP7_75t_L g5674 ( 
.A1(n_5374),
.A2(n_2287),
.B1(n_2186),
.B2(n_2193),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5324),
.Y(n_5675)
);

OAI22xp5_ASAP7_75t_L g5676 ( 
.A1(n_5105),
.A2(n_1150),
.B1(n_1157),
.B2(n_1151),
.Y(n_5676)
);

NAND2xp5_ASAP7_75t_L g5677 ( 
.A(n_5316),
.B(n_13),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_5349),
.Y(n_5678)
);

OAI21xp5_ASAP7_75t_SL g5679 ( 
.A1(n_5358),
.A2(n_13),
.B(n_14),
.Y(n_5679)
);

CKINVDCx5p33_ASAP7_75t_R g5680 ( 
.A(n_5323),
.Y(n_5680)
);

BUFx8_ASAP7_75t_L g5681 ( 
.A(n_5359),
.Y(n_5681)
);

OAI222xp33_ASAP7_75t_L g5682 ( 
.A1(n_5140),
.A2(n_1162),
.B1(n_1158),
.B2(n_1167),
.C1(n_1163),
.C2(n_1148),
.Y(n_5682)
);

INVx1_ASAP7_75t_SL g5683 ( 
.A(n_5351),
.Y(n_5683)
);

INVx2_ASAP7_75t_L g5684 ( 
.A(n_4986),
.Y(n_5684)
);

AND2x4_ASAP7_75t_L g5685 ( 
.A(n_5291),
.B(n_1348),
.Y(n_5685)
);

NAND2x1p5_ASAP7_75t_L g5686 ( 
.A(n_5377),
.B(n_3333),
.Y(n_5686)
);

OAI21x1_ASAP7_75t_L g5687 ( 
.A1(n_5314),
.A2(n_2593),
.B(n_2592),
.Y(n_5687)
);

NOR2xp33_ASAP7_75t_L g5688 ( 
.A(n_5079),
.B(n_15),
.Y(n_5688)
);

NAND2x1p5_ASAP7_75t_L g5689 ( 
.A(n_5334),
.B(n_3377),
.Y(n_5689)
);

BUFx3_ASAP7_75t_L g5690 ( 
.A(n_5320),
.Y(n_5690)
);

AOI21x1_ASAP7_75t_L g5691 ( 
.A1(n_5132),
.A2(n_1352),
.B(n_1351),
.Y(n_5691)
);

NAND4xp25_ASAP7_75t_L g5692 ( 
.A(n_5352),
.B(n_2306),
.C(n_17),
.D(n_15),
.Y(n_5692)
);

OAI22xp33_ASAP7_75t_SL g5693 ( 
.A1(n_5302),
.A2(n_5306),
.B1(n_5142),
.B2(n_5179),
.Y(n_5693)
);

OAI21x1_ASAP7_75t_L g5694 ( 
.A1(n_5282),
.A2(n_2593),
.B(n_2832),
.Y(n_5694)
);

OAI21x1_ASAP7_75t_L g5695 ( 
.A1(n_5060),
.A2(n_2832),
.B(n_2826),
.Y(n_5695)
);

OAI21xp5_ASAP7_75t_L g5696 ( 
.A1(n_4988),
.A2(n_1168),
.B(n_1159),
.Y(n_5696)
);

BUFx2_ASAP7_75t_SL g5697 ( 
.A(n_5133),
.Y(n_5697)
);

AOI22xp33_ASAP7_75t_L g5698 ( 
.A1(n_5374),
.A2(n_2186),
.B1(n_2193),
.B2(n_2182),
.Y(n_5698)
);

NAND2x1p5_ASAP7_75t_L g5699 ( 
.A(n_5133),
.B(n_2627),
.Y(n_5699)
);

OA21x2_ASAP7_75t_L g5700 ( 
.A1(n_5155),
.A2(n_1357),
.B(n_1352),
.Y(n_5700)
);

OAI21x1_ASAP7_75t_L g5701 ( 
.A1(n_5349),
.A2(n_2826),
.B(n_2817),
.Y(n_5701)
);

AND2x4_ASAP7_75t_L g5702 ( 
.A(n_5133),
.B(n_1357),
.Y(n_5702)
);

OAI21x1_ASAP7_75t_L g5703 ( 
.A1(n_5173),
.A2(n_2826),
.B(n_2817),
.Y(n_5703)
);

NAND2x1_ASAP7_75t_L g5704 ( 
.A(n_5161),
.B(n_5232),
.Y(n_5704)
);

OA21x2_ASAP7_75t_L g5705 ( 
.A1(n_5155),
.A2(n_1358),
.B(n_1174),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5245),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_4986),
.Y(n_5707)
);

INVx2_ASAP7_75t_SL g5708 ( 
.A(n_5161),
.Y(n_5708)
);

OAI22xp5_ASAP7_75t_L g5709 ( 
.A1(n_5113),
.A2(n_1175),
.B1(n_1176),
.B2(n_1173),
.Y(n_5709)
);

AND2x2_ASAP7_75t_L g5710 ( 
.A(n_5161),
.B(n_16),
.Y(n_5710)
);

OAI21x1_ASAP7_75t_L g5711 ( 
.A1(n_5268),
.A2(n_2833),
.B(n_2817),
.Y(n_5711)
);

AOI21xp5_ASAP7_75t_L g5712 ( 
.A1(n_5069),
.A2(n_2632),
.B(n_2627),
.Y(n_5712)
);

INVx3_ASAP7_75t_L g5713 ( 
.A(n_5232),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5232),
.B(n_16),
.Y(n_5714)
);

AO21x2_ASAP7_75t_L g5715 ( 
.A1(n_5139),
.A2(n_1358),
.B(n_2311),
.Y(n_5715)
);

OA21x2_ASAP7_75t_L g5716 ( 
.A1(n_5179),
.A2(n_5139),
.B(n_5188),
.Y(n_5716)
);

OA21x2_ASAP7_75t_L g5717 ( 
.A1(n_5188),
.A2(n_1195),
.B(n_1194),
.Y(n_5717)
);

INVx2_ASAP7_75t_SL g5718 ( 
.A(n_5357),
.Y(n_5718)
);

OAI221xp5_ASAP7_75t_L g5719 ( 
.A1(n_5045),
.A2(n_1204),
.B1(n_1222),
.B2(n_1203),
.C(n_1199),
.Y(n_5719)
);

OAI21x1_ASAP7_75t_SL g5720 ( 
.A1(n_5300),
.A2(n_5384),
.B(n_5339),
.Y(n_5720)
);

NAND2x1p5_ASAP7_75t_L g5721 ( 
.A(n_5357),
.B(n_5154),
.Y(n_5721)
);

NOR2x1_ASAP7_75t_SL g5722 ( 
.A(n_5357),
.B(n_1280),
.Y(n_5722)
);

INVxp67_ASAP7_75t_SL g5723 ( 
.A(n_5154),
.Y(n_5723)
);

AND2x2_ASAP7_75t_L g5724 ( 
.A(n_4999),
.B(n_16),
.Y(n_5724)
);

OAI21x1_ASAP7_75t_L g5725 ( 
.A1(n_5198),
.A2(n_2833),
.B(n_2632),
.Y(n_5725)
);

OAI21x1_ASAP7_75t_L g5726 ( 
.A1(n_5208),
.A2(n_2833),
.B(n_2632),
.Y(n_5726)
);

AOI21x1_ASAP7_75t_L g5727 ( 
.A1(n_5368),
.A2(n_1333),
.B(n_1292),
.Y(n_5727)
);

INVx3_ASAP7_75t_L g5728 ( 
.A(n_5180),
.Y(n_5728)
);

AND2x4_ASAP7_75t_L g5729 ( 
.A(n_5180),
.B(n_17),
.Y(n_5729)
);

BUFx6f_ASAP7_75t_L g5730 ( 
.A(n_5181),
.Y(n_5730)
);

AOI22xp33_ASAP7_75t_L g5731 ( 
.A1(n_5372),
.A2(n_2193),
.B1(n_2229),
.B2(n_2182),
.Y(n_5731)
);

HB1xp67_ASAP7_75t_L g5732 ( 
.A(n_5056),
.Y(n_5732)
);

INVx4_ASAP7_75t_SL g5733 ( 
.A(n_5041),
.Y(n_5733)
);

AO31x2_ASAP7_75t_L g5734 ( 
.A1(n_5214),
.A2(n_1293),
.A3(n_1290),
.B(n_2310),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5316),
.Y(n_5735)
);

CKINVDCx6p67_ASAP7_75t_R g5736 ( 
.A(n_5432),
.Y(n_5736)
);

NOR2xp33_ASAP7_75t_L g5737 ( 
.A(n_5411),
.B(n_5119),
.Y(n_5737)
);

OR2x2_ASAP7_75t_L g5738 ( 
.A(n_5443),
.B(n_5181),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_L g5739 ( 
.A(n_5585),
.B(n_5385),
.Y(n_5739)
);

INVx5_ASAP7_75t_L g5740 ( 
.A(n_5491),
.Y(n_5740)
);

INVx2_ASAP7_75t_L g5741 ( 
.A(n_5532),
.Y(n_5741)
);

AOI22xp33_ASAP7_75t_L g5742 ( 
.A1(n_5391),
.A2(n_5370),
.B1(n_5290),
.B2(n_5294),
.Y(n_5742)
);

OAI221xp5_ASAP7_75t_L g5743 ( 
.A1(n_5591),
.A2(n_5330),
.B1(n_5342),
.B2(n_5205),
.C(n_5096),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5547),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5547),
.Y(n_5745)
);

OAI22xp5_ASAP7_75t_L g5746 ( 
.A1(n_5591),
.A2(n_5257),
.B1(n_5095),
.B2(n_5080),
.Y(n_5746)
);

INVx2_ASAP7_75t_SL g5747 ( 
.A(n_5491),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5573),
.Y(n_5748)
);

OAI22xp33_ASAP7_75t_L g5749 ( 
.A1(n_5391),
.A2(n_4999),
.B1(n_5054),
.B2(n_5331),
.Y(n_5749)
);

HB1xp67_ASAP7_75t_L g5750 ( 
.A(n_5397),
.Y(n_5750)
);

OAI22xp5_ASAP7_75t_L g5751 ( 
.A1(n_5392),
.A2(n_5358),
.B1(n_5146),
.B2(n_5145),
.Y(n_5751)
);

NAND2xp5_ASAP7_75t_SL g5752 ( 
.A(n_5607),
.B(n_5321),
.Y(n_5752)
);

INVx1_ASAP7_75t_L g5753 ( 
.A(n_5573),
.Y(n_5753)
);

OAI22xp5_ASAP7_75t_L g5754 ( 
.A1(n_5392),
.A2(n_5183),
.B1(n_5152),
.B2(n_5336),
.Y(n_5754)
);

NAND2xp5_ASAP7_75t_L g5755 ( 
.A(n_5585),
.B(n_5553),
.Y(n_5755)
);

AND2x4_ASAP7_75t_L g5756 ( 
.A(n_5639),
.B(n_5735),
.Y(n_5756)
);

NAND2xp5_ASAP7_75t_L g5757 ( 
.A(n_5572),
.B(n_5149),
.Y(n_5757)
);

AOI22xp33_ASAP7_75t_L g5758 ( 
.A1(n_5724),
.A2(n_5290),
.B1(n_5106),
.B2(n_5387),
.Y(n_5758)
);

CKINVDCx20_ASAP7_75t_R g5759 ( 
.A(n_5422),
.Y(n_5759)
);

AOI21xp5_ASAP7_75t_L g5760 ( 
.A1(n_5461),
.A2(n_5124),
.B(n_5061),
.Y(n_5760)
);

OR2x6_ASAP7_75t_L g5761 ( 
.A(n_5574),
.B(n_5335),
.Y(n_5761)
);

BUFx6f_ASAP7_75t_L g5762 ( 
.A(n_5491),
.Y(n_5762)
);

OAI22xp5_ASAP7_75t_L g5763 ( 
.A1(n_5421),
.A2(n_5166),
.B1(n_5150),
.B2(n_5158),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5443),
.Y(n_5764)
);

NAND2xp5_ASAP7_75t_L g5765 ( 
.A(n_5639),
.B(n_5149),
.Y(n_5765)
);

OAI22xp5_ASAP7_75t_L g5766 ( 
.A1(n_5431),
.A2(n_5315),
.B1(n_5361),
.B2(n_5293),
.Y(n_5766)
);

AOI22xp33_ASAP7_75t_L g5767 ( 
.A1(n_5599),
.A2(n_5106),
.B1(n_5387),
.B2(n_5292),
.Y(n_5767)
);

CKINVDCx20_ASAP7_75t_R g5768 ( 
.A(n_5629),
.Y(n_5768)
);

NAND3xp33_ASAP7_75t_SL g5769 ( 
.A(n_5663),
.B(n_5046),
.C(n_5037),
.Y(n_5769)
);

OAI22xp5_ASAP7_75t_L g5770 ( 
.A1(n_5431),
.A2(n_5679),
.B1(n_5696),
.B2(n_5599),
.Y(n_5770)
);

INVx2_ASAP7_75t_L g5771 ( 
.A(n_5465),
.Y(n_5771)
);

OR2x2_ASAP7_75t_L g5772 ( 
.A(n_5397),
.B(n_5402),
.Y(n_5772)
);

AOI22xp33_ASAP7_75t_L g5773 ( 
.A1(n_5692),
.A2(n_5292),
.B1(n_5275),
.B2(n_5212),
.Y(n_5773)
);

AOI22xp5_ASAP7_75t_L g5774 ( 
.A1(n_5696),
.A2(n_5400),
.B1(n_5555),
.B2(n_5488),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5454),
.Y(n_5775)
);

OR2x2_ASAP7_75t_L g5776 ( 
.A(n_5402),
.B(n_5003),
.Y(n_5776)
);

AOI22xp33_ASAP7_75t_L g5777 ( 
.A1(n_5555),
.A2(n_5275),
.B1(n_5215),
.B2(n_5315),
.Y(n_5777)
);

OR2x2_ASAP7_75t_L g5778 ( 
.A(n_5406),
.B(n_5003),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5509),
.Y(n_5779)
);

INVx2_ASAP7_75t_L g5780 ( 
.A(n_5509),
.Y(n_5780)
);

INVx2_ASAP7_75t_L g5781 ( 
.A(n_5510),
.Y(n_5781)
);

INVx3_ASAP7_75t_L g5782 ( 
.A(n_5651),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_5467),
.Y(n_5783)
);

AOI22xp33_ASAP7_75t_SL g5784 ( 
.A1(n_5499),
.A2(n_5230),
.B1(n_5017),
.B2(n_5172),
.Y(n_5784)
);

OR2x6_ASAP7_75t_SL g5785 ( 
.A(n_5680),
.B(n_1224),
.Y(n_5785)
);

INVx2_ASAP7_75t_SL g5786 ( 
.A(n_5564),
.Y(n_5786)
);

AND2x4_ASAP7_75t_L g5787 ( 
.A(n_5607),
.B(n_5418),
.Y(n_5787)
);

OAI22xp5_ASAP7_75t_L g5788 ( 
.A1(n_5413),
.A2(n_5049),
.B1(n_5190),
.B2(n_5073),
.Y(n_5788)
);

NAND2x1_ASAP7_75t_L g5789 ( 
.A(n_5439),
.B(n_5429),
.Y(n_5789)
);

OR2x6_ASAP7_75t_L g5790 ( 
.A(n_5574),
.B(n_5508),
.Y(n_5790)
);

BUFx3_ASAP7_75t_L g5791 ( 
.A(n_5514),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_5472),
.Y(n_5792)
);

INVx3_ASAP7_75t_L g5793 ( 
.A(n_5439),
.Y(n_5793)
);

AND2x2_ASAP7_75t_L g5794 ( 
.A(n_5437),
.B(n_5017),
.Y(n_5794)
);

O2A1O1Ixp33_ASAP7_75t_SL g5795 ( 
.A1(n_5427),
.A2(n_5024),
.B(n_5256),
.C(n_5167),
.Y(n_5795)
);

NAND2xp5_ASAP7_75t_SL g5796 ( 
.A(n_5607),
.B(n_5206),
.Y(n_5796)
);

NAND2xp5_ASAP7_75t_L g5797 ( 
.A(n_5406),
.B(n_5561),
.Y(n_5797)
);

INVx2_ASAP7_75t_SL g5798 ( 
.A(n_5625),
.Y(n_5798)
);

OAI22xp5_ASAP7_75t_L g5799 ( 
.A1(n_5413),
.A2(n_5192),
.B1(n_5236),
.B2(n_5242),
.Y(n_5799)
);

OAI22xp33_ASAP7_75t_L g5800 ( 
.A1(n_5652),
.A2(n_5213),
.B1(n_5108),
.B2(n_5120),
.Y(n_5800)
);

AOI22xp33_ASAP7_75t_SL g5801 ( 
.A1(n_5499),
.A2(n_5172),
.B1(n_5003),
.B2(n_5041),
.Y(n_5801)
);

INVx5_ASAP7_75t_L g5802 ( 
.A(n_5538),
.Y(n_5802)
);

AOI221xp5_ASAP7_75t_L g5803 ( 
.A1(n_5583),
.A2(n_1231),
.B1(n_1236),
.B2(n_1227),
.C(n_1225),
.Y(n_5803)
);

HB1xp67_ASAP7_75t_L g5804 ( 
.A(n_5430),
.Y(n_5804)
);

OR2x6_ASAP7_75t_L g5805 ( 
.A(n_5508),
.B(n_5235),
.Y(n_5805)
);

NAND2xp33_ASAP7_75t_R g5806 ( 
.A(n_5646),
.B(n_18),
.Y(n_5806)
);

CKINVDCx8_ASAP7_75t_R g5807 ( 
.A(n_5598),
.Y(n_5807)
);

OAI22xp33_ASAP7_75t_L g5808 ( 
.A1(n_5652),
.A2(n_5287),
.B1(n_5041),
.B2(n_5319),
.Y(n_5808)
);

AOI21xp5_ASAP7_75t_L g5809 ( 
.A1(n_5415),
.A2(n_5126),
.B(n_5112),
.Y(n_5809)
);

BUFx2_ASAP7_75t_L g5810 ( 
.A(n_5423),
.Y(n_5810)
);

NAND2xp5_ASAP7_75t_L g5811 ( 
.A(n_5561),
.B(n_5149),
.Y(n_5811)
);

OAI21x1_ASAP7_75t_L g5812 ( 
.A1(n_5412),
.A2(n_5356),
.B(n_5286),
.Y(n_5812)
);

AOI22xp33_ASAP7_75t_L g5813 ( 
.A1(n_5705),
.A2(n_2233),
.B1(n_2229),
.B2(n_5211),
.Y(n_5813)
);

NAND2xp33_ASAP7_75t_R g5814 ( 
.A(n_5521),
.B(n_18),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5479),
.Y(n_5815)
);

NOR2x1_ASAP7_75t_SL g5816 ( 
.A(n_5607),
.B(n_5034),
.Y(n_5816)
);

CKINVDCx6p67_ASAP7_75t_R g5817 ( 
.A(n_5562),
.Y(n_5817)
);

BUFx6f_ASAP7_75t_L g5818 ( 
.A(n_5538),
.Y(n_5818)
);

AOI22xp33_ASAP7_75t_SL g5819 ( 
.A1(n_5705),
.A2(n_5172),
.B1(n_4986),
.B2(n_1239),
.Y(n_5819)
);

AOI22xp33_ASAP7_75t_SL g5820 ( 
.A1(n_5677),
.A2(n_1241),
.B1(n_1238),
.B2(n_5239),
.Y(n_5820)
);

INVx1_ASAP7_75t_SL g5821 ( 
.A(n_5427),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5481),
.Y(n_5822)
);

OR2x6_ASAP7_75t_L g5823 ( 
.A(n_5508),
.B(n_5107),
.Y(n_5823)
);

INVx4_ASAP7_75t_L g5824 ( 
.A(n_5411),
.Y(n_5824)
);

OAI22xp5_ASAP7_75t_L g5825 ( 
.A1(n_5677),
.A2(n_5219),
.B1(n_5307),
.B2(n_5376),
.Y(n_5825)
);

AND2x4_ASAP7_75t_L g5826 ( 
.A(n_5394),
.B(n_5034),
.Y(n_5826)
);

AOI22xp33_ASAP7_75t_L g5827 ( 
.A1(n_5415),
.A2(n_2233),
.B1(n_2229),
.B2(n_2304),
.Y(n_5827)
);

NOR2x1_ASAP7_75t_SL g5828 ( 
.A(n_5571),
.B(n_5668),
.Y(n_5828)
);

AOI22xp33_ASAP7_75t_L g5829 ( 
.A1(n_5717),
.A2(n_2233),
.B1(n_2229),
.B2(n_2304),
.Y(n_5829)
);

OR2x2_ASAP7_75t_L g5830 ( 
.A(n_5489),
.B(n_5034),
.Y(n_5830)
);

BUFx2_ASAP7_75t_L g5831 ( 
.A(n_5414),
.Y(n_5831)
);

AOI221xp5_ASAP7_75t_L g5832 ( 
.A1(n_5583),
.A2(n_5070),
.B1(n_5153),
.B2(n_5273),
.C(n_5272),
.Y(n_5832)
);

AND2x2_ASAP7_75t_L g5833 ( 
.A(n_5537),
.B(n_5056),
.Y(n_5833)
);

OAI22xp33_ASAP7_75t_SL g5834 ( 
.A1(n_5453),
.A2(n_4984),
.B1(n_21),
.B2(n_19),
.Y(n_5834)
);

OA21x2_ASAP7_75t_L g5835 ( 
.A1(n_5399),
.A2(n_5322),
.B(n_5328),
.Y(n_5835)
);

BUFx3_ASAP7_75t_L g5836 ( 
.A(n_5408),
.Y(n_5836)
);

INVxp67_ASAP7_75t_L g5837 ( 
.A(n_5395),
.Y(n_5837)
);

OAI21xp5_ASAP7_75t_L g5838 ( 
.A1(n_5558),
.A2(n_5182),
.B(n_5338),
.Y(n_5838)
);

OAI22xp5_ASAP7_75t_L g5839 ( 
.A1(n_5723),
.A2(n_5565),
.B1(n_5634),
.B2(n_5471),
.Y(n_5839)
);

BUFx4f_ASAP7_75t_SL g5840 ( 
.A(n_5589),
.Y(n_5840)
);

CKINVDCx20_ASAP7_75t_R g5841 ( 
.A(n_5451),
.Y(n_5841)
);

INVx4_ASAP7_75t_L g5842 ( 
.A(n_5589),
.Y(n_5842)
);

CKINVDCx8_ASAP7_75t_R g5843 ( 
.A(n_5729),
.Y(n_5843)
);

AND2x4_ASAP7_75t_L g5844 ( 
.A(n_5394),
.B(n_5056),
.Y(n_5844)
);

INVx2_ASAP7_75t_L g5845 ( 
.A(n_5510),
.Y(n_5845)
);

CKINVDCx6p67_ASAP7_75t_R g5846 ( 
.A(n_5451),
.Y(n_5846)
);

AOI21xp33_ASAP7_75t_L g5847 ( 
.A1(n_5435),
.A2(n_5526),
.B(n_5716),
.Y(n_5847)
);

OR2x6_ASAP7_75t_L g5848 ( 
.A(n_5613),
.B(n_5355),
.Y(n_5848)
);

NAND2xp5_ASAP7_75t_L g5849 ( 
.A(n_5489),
.B(n_5059),
.Y(n_5849)
);

BUFx2_ASAP7_75t_L g5850 ( 
.A(n_5414),
.Y(n_5850)
);

OAI22xp33_ASAP7_75t_L g5851 ( 
.A1(n_5557),
.A2(n_5085),
.B1(n_5123),
.B2(n_5059),
.Y(n_5851)
);

OAI22xp5_ASAP7_75t_L g5852 ( 
.A1(n_5723),
.A2(n_2633),
.B1(n_2683),
.B2(n_2627),
.Y(n_5852)
);

AOI22xp33_ASAP7_75t_L g5853 ( 
.A1(n_5717),
.A2(n_2233),
.B1(n_2229),
.B2(n_2304),
.Y(n_5853)
);

BUFx3_ASAP7_75t_L g5854 ( 
.A(n_5618),
.Y(n_5854)
);

AOI22xp33_ASAP7_75t_L g5855 ( 
.A1(n_5400),
.A2(n_2233),
.B1(n_2307),
.B2(n_2304),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5540),
.Y(n_5856)
);

NOR2xp33_ASAP7_75t_L g5857 ( 
.A(n_5606),
.B(n_164),
.Y(n_5857)
);

AND2x4_ASAP7_75t_L g5858 ( 
.A(n_5394),
.B(n_5059),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5410),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5425),
.Y(n_5860)
);

AND2x2_ASAP7_75t_L g5861 ( 
.A(n_5641),
.B(n_5337),
.Y(n_5861)
);

AND2x2_ASAP7_75t_L g5862 ( 
.A(n_5420),
.B(n_5512),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5438),
.Y(n_5863)
);

NAND2x1_ASAP7_75t_L g5864 ( 
.A(n_5394),
.B(n_5085),
.Y(n_5864)
);

INVx2_ASAP7_75t_L g5865 ( 
.A(n_5498),
.Y(n_5865)
);

OAI22xp33_ASAP7_75t_L g5866 ( 
.A1(n_5557),
.A2(n_5123),
.B1(n_5085),
.B2(n_4984),
.Y(n_5866)
);

INVx2_ASAP7_75t_L g5867 ( 
.A(n_5435),
.Y(n_5867)
);

OR2x6_ASAP7_75t_L g5868 ( 
.A(n_5613),
.B(n_5362),
.Y(n_5868)
);

OR2x2_ASAP7_75t_L g5869 ( 
.A(n_5546),
.B(n_5123),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5486),
.Y(n_5870)
);

BUFx3_ASAP7_75t_L g5871 ( 
.A(n_5424),
.Y(n_5871)
);

NAND2xp5_ASAP7_75t_L g5872 ( 
.A(n_5457),
.B(n_5337),
.Y(n_5872)
);

OR2x2_ASAP7_75t_L g5873 ( 
.A(n_5628),
.B(n_5337),
.Y(n_5873)
);

AOI21xp5_ASAP7_75t_L g5874 ( 
.A1(n_5579),
.A2(n_5118),
.B(n_5189),
.Y(n_5874)
);

AND2x2_ASAP7_75t_L g5875 ( 
.A(n_5617),
.B(n_5360),
.Y(n_5875)
);

INVx2_ASAP7_75t_L g5876 ( 
.A(n_5486),
.Y(n_5876)
);

NOR2xp33_ASAP7_75t_SL g5877 ( 
.A(n_5571),
.B(n_5360),
.Y(n_5877)
);

AOI22xp33_ASAP7_75t_L g5878 ( 
.A1(n_5602),
.A2(n_2307),
.B1(n_5297),
.B2(n_5295),
.Y(n_5878)
);

INVx2_ASAP7_75t_L g5879 ( 
.A(n_5396),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5449),
.Y(n_5880)
);

OR2x6_ASAP7_75t_L g5881 ( 
.A(n_5550),
.B(n_5378),
.Y(n_5881)
);

INVx2_ASAP7_75t_L g5882 ( 
.A(n_5417),
.Y(n_5882)
);

INVx3_ASAP7_75t_L g5883 ( 
.A(n_5577),
.Y(n_5883)
);

OAI22xp5_ASAP7_75t_L g5884 ( 
.A1(n_5565),
.A2(n_2633),
.B1(n_2691),
.B2(n_2683),
.Y(n_5884)
);

AO31x2_ASAP7_75t_L g5885 ( 
.A1(n_5403),
.A2(n_5301),
.A3(n_4984),
.B(n_5360),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5627),
.Y(n_5886)
);

INVx2_ASAP7_75t_L g5887 ( 
.A(n_5464),
.Y(n_5887)
);

AOI21xp33_ASAP7_75t_L g5888 ( 
.A1(n_5716),
.A2(n_19),
.B(n_20),
.Y(n_5888)
);

AOI222xp33_ASAP7_75t_L g5889 ( 
.A1(n_5419),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.C1(n_21),
.C2(n_23),
.Y(n_5889)
);

CKINVDCx16_ASAP7_75t_R g5890 ( 
.A(n_5516),
.Y(n_5890)
);

AOI221xp5_ASAP7_75t_L g5891 ( 
.A1(n_5558),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.C(n_23),
.Y(n_5891)
);

AOI221xp5_ASAP7_75t_L g5892 ( 
.A1(n_5635),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.C(n_26),
.Y(n_5892)
);

INVxp67_ASAP7_75t_L g5893 ( 
.A(n_5395),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5428),
.Y(n_5894)
);

AOI22xp33_ASAP7_75t_L g5895 ( 
.A1(n_5602),
.A2(n_2307),
.B1(n_5311),
.B2(n_5305),
.Y(n_5895)
);

INVx1_ASAP7_75t_SL g5896 ( 
.A(n_5626),
.Y(n_5896)
);

NAND2xp5_ASAP7_75t_L g5897 ( 
.A(n_5523),
.B(n_5253),
.Y(n_5897)
);

NAND3xp33_ASAP7_75t_SL g5898 ( 
.A(n_5579),
.B(n_24),
.C(n_26),
.Y(n_5898)
);

OAI21xp5_ASAP7_75t_L g5899 ( 
.A1(n_5416),
.A2(n_5380),
.B(n_5068),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5428),
.Y(n_5900)
);

INVx3_ASAP7_75t_L g5901 ( 
.A(n_5577),
.Y(n_5901)
);

BUFx6f_ASAP7_75t_L g5902 ( 
.A(n_5390),
.Y(n_5902)
);

AND2x2_ASAP7_75t_L g5903 ( 
.A(n_5649),
.B(n_5253),
.Y(n_5903)
);

OAI211xp5_ASAP7_75t_L g5904 ( 
.A1(n_5419),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_5904)
);

OAI21x1_ASAP7_75t_L g5905 ( 
.A1(n_5433),
.A2(n_5075),
.B(n_5194),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_5575),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5580),
.Y(n_5907)
);

BUFx6f_ASAP7_75t_L g5908 ( 
.A(n_5390),
.Y(n_5908)
);

HB1xp67_ASAP7_75t_L g5909 ( 
.A(n_5484),
.Y(n_5909)
);

NAND2xp5_ASAP7_75t_L g5910 ( 
.A(n_5523),
.B(n_5551),
.Y(n_5910)
);

AOI221xp5_ASAP7_75t_L g5911 ( 
.A1(n_5693),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.C(n_30),
.Y(n_5911)
);

A2O1A1Ixp33_ASAP7_75t_SL g5912 ( 
.A1(n_5459),
.A2(n_2306),
.B(n_2683),
.C(n_2633),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5576),
.Y(n_5913)
);

AOI21x1_ASAP7_75t_L g5914 ( 
.A1(n_5405),
.A2(n_5253),
.B(n_5216),
.Y(n_5914)
);

HB1xp67_ASAP7_75t_L g5915 ( 
.A(n_5484),
.Y(n_5915)
);

A2O1A1Ixp33_ASAP7_75t_L g5916 ( 
.A1(n_5657),
.A2(n_31),
.B(n_27),
.C(n_30),
.Y(n_5916)
);

OR2x6_ASAP7_75t_L g5917 ( 
.A(n_5550),
.B(n_5207),
.Y(n_5917)
);

HB1xp67_ASAP7_75t_L g5918 ( 
.A(n_5487),
.Y(n_5918)
);

AOI22xp33_ASAP7_75t_L g5919 ( 
.A1(n_5517),
.A2(n_2307),
.B1(n_2314),
.B2(n_2310),
.Y(n_5919)
);

INVx2_ASAP7_75t_L g5920 ( 
.A(n_5504),
.Y(n_5920)
);

AND2x4_ASAP7_75t_L g5921 ( 
.A(n_5394),
.B(n_5207),
.Y(n_5921)
);

CKINVDCx5p33_ASAP7_75t_R g5922 ( 
.A(n_5548),
.Y(n_5922)
);

OAI22xp5_ASAP7_75t_L g5923 ( 
.A1(n_5483),
.A2(n_2691),
.B1(n_2701),
.B2(n_2692),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5551),
.Y(n_5924)
);

BUFx3_ASAP7_75t_L g5925 ( 
.A(n_5681),
.Y(n_5925)
);

OAI22xp5_ASAP7_75t_L g5926 ( 
.A1(n_5483),
.A2(n_2691),
.B1(n_2701),
.B2(n_2692),
.Y(n_5926)
);

AND2x2_ASAP7_75t_L g5927 ( 
.A(n_5541),
.B(n_5207),
.Y(n_5927)
);

OAI22xp5_ASAP7_75t_L g5928 ( 
.A1(n_5483),
.A2(n_2692),
.B1(n_2722),
.B2(n_2701),
.Y(n_5928)
);

OAI22xp33_ASAP7_75t_L g5929 ( 
.A1(n_5600),
.A2(n_3031),
.B1(n_2722),
.B2(n_2762),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5506),
.Y(n_5930)
);

NAND2xp5_ASAP7_75t_L g5931 ( 
.A(n_5446),
.B(n_5216),
.Y(n_5931)
);

AND2x2_ASAP7_75t_L g5932 ( 
.A(n_5545),
.B(n_5216),
.Y(n_5932)
);

CKINVDCx5p33_ASAP7_75t_R g5933 ( 
.A(n_5631),
.Y(n_5933)
);

AND2x4_ASAP7_75t_L g5934 ( 
.A(n_5404),
.B(n_5227),
.Y(n_5934)
);

INVx4_ASAP7_75t_L g5935 ( 
.A(n_5401),
.Y(n_5935)
);

AND2x2_ASAP7_75t_L g5936 ( 
.A(n_5490),
.B(n_5227),
.Y(n_5936)
);

BUFx3_ASAP7_75t_L g5937 ( 
.A(n_5681),
.Y(n_5937)
);

NAND2xp5_ASAP7_75t_L g5938 ( 
.A(n_5446),
.B(n_5501),
.Y(n_5938)
);

AND2x4_ASAP7_75t_L g5939 ( 
.A(n_5442),
.B(n_5227),
.Y(n_5939)
);

AOI21xp5_ASAP7_75t_L g5940 ( 
.A1(n_5720),
.A2(n_2751),
.B(n_2722),
.Y(n_5940)
);

AOI22xp33_ASAP7_75t_L g5941 ( 
.A1(n_5517),
.A2(n_2307),
.B1(n_2319),
.B2(n_2314),
.Y(n_5941)
);

NAND2xp33_ASAP7_75t_R g5942 ( 
.A(n_5654),
.B(n_30),
.Y(n_5942)
);

AOI22xp33_ASAP7_75t_L g5943 ( 
.A1(n_5531),
.A2(n_2319),
.B1(n_2316),
.B2(n_2317),
.Y(n_5943)
);

INVx6_ASAP7_75t_L g5944 ( 
.A(n_5516),
.Y(n_5944)
);

NAND2xp5_ASAP7_75t_L g5945 ( 
.A(n_5501),
.B(n_5251),
.Y(n_5945)
);

NAND3xp33_ASAP7_75t_SL g5946 ( 
.A(n_5524),
.B(n_31),
.C(n_32),
.Y(n_5946)
);

NAND2xp33_ASAP7_75t_SL g5947 ( 
.A(n_5401),
.B(n_31),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5632),
.B(n_5251),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_5507),
.B(n_5251),
.Y(n_5949)
);

CKINVDCx6p67_ASAP7_75t_R g5950 ( 
.A(n_5393),
.Y(n_5950)
);

AOI22xp33_ASAP7_75t_L g5951 ( 
.A1(n_5531),
.A2(n_5715),
.B1(n_5706),
.B2(n_5436),
.Y(n_5951)
);

AND2x4_ASAP7_75t_L g5952 ( 
.A(n_5442),
.B(n_5332),
.Y(n_5952)
);

AOI22xp33_ASAP7_75t_L g5953 ( 
.A1(n_5715),
.A2(n_2316),
.B1(n_2317),
.B2(n_2311),
.Y(n_5953)
);

AOI22xp33_ASAP7_75t_L g5954 ( 
.A1(n_5436),
.A2(n_5633),
.B1(n_5488),
.B2(n_5630),
.Y(n_5954)
);

NAND2xp5_ASAP7_75t_L g5955 ( 
.A(n_5507),
.B(n_5332),
.Y(n_5955)
);

AOI22xp33_ASAP7_75t_L g5956 ( 
.A1(n_5581),
.A2(n_2762),
.B1(n_2805),
.B2(n_2751),
.Y(n_5956)
);

NAND2xp5_ASAP7_75t_L g5957 ( 
.A(n_5476),
.B(n_5332),
.Y(n_5957)
);

NAND3xp33_ASAP7_75t_SL g5958 ( 
.A(n_5524),
.B(n_32),
.C(n_33),
.Y(n_5958)
);

HB1xp67_ASAP7_75t_L g5959 ( 
.A(n_5487),
.Y(n_5959)
);

A2O1A1Ixp33_ASAP7_75t_L g5960 ( 
.A1(n_5657),
.A2(n_5416),
.B(n_5601),
.C(n_5552),
.Y(n_5960)
);

OAI22xp33_ASAP7_75t_L g5961 ( 
.A1(n_5600),
.A2(n_3031),
.B1(n_2762),
.B2(n_2805),
.Y(n_5961)
);

INVx2_ASAP7_75t_L g5962 ( 
.A(n_5453),
.Y(n_5962)
);

NAND2xp5_ASAP7_75t_L g5963 ( 
.A(n_5476),
.B(n_5450),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5462),
.Y(n_5964)
);

NAND2xp5_ASAP7_75t_L g5965 ( 
.A(n_5452),
.B(n_5277),
.Y(n_5965)
);

CKINVDCx16_ASAP7_75t_R g5966 ( 
.A(n_5393),
.Y(n_5966)
);

INVx2_ASAP7_75t_L g5967 ( 
.A(n_5597),
.Y(n_5967)
);

BUFx2_ASAP7_75t_SL g5968 ( 
.A(n_5671),
.Y(n_5968)
);

OR2x2_ASAP7_75t_L g5969 ( 
.A(n_5480),
.B(n_5367),
.Y(n_5969)
);

BUFx4f_ASAP7_75t_SL g5970 ( 
.A(n_5409),
.Y(n_5970)
);

INVx2_ASAP7_75t_L g5971 ( 
.A(n_5604),
.Y(n_5971)
);

HB1xp67_ASAP7_75t_L g5972 ( 
.A(n_5441),
.Y(n_5972)
);

NAND2x1p5_ASAP7_75t_L g5973 ( 
.A(n_5571),
.B(n_2751),
.Y(n_5973)
);

OAI22xp5_ASAP7_75t_L g5974 ( 
.A1(n_5728),
.A2(n_2807),
.B1(n_2805),
.B2(n_35),
.Y(n_5974)
);

BUFx2_ASAP7_75t_L g5975 ( 
.A(n_5593),
.Y(n_5975)
);

INVx2_ASAP7_75t_L g5976 ( 
.A(n_5661),
.Y(n_5976)
);

OAI222xp33_ASAP7_75t_L g5977 ( 
.A1(n_5581),
.A2(n_5284),
.B1(n_5277),
.B2(n_5369),
.C1(n_5367),
.C2(n_35),
.Y(n_5977)
);

OAI22xp5_ASAP7_75t_L g5978 ( 
.A1(n_5728),
.A2(n_2807),
.B1(n_35),
.B2(n_33),
.Y(n_5978)
);

NAND2xp5_ASAP7_75t_L g5979 ( 
.A(n_5494),
.B(n_5277),
.Y(n_5979)
);

INVx3_ASAP7_75t_L g5980 ( 
.A(n_5593),
.Y(n_5980)
);

AOI21xp5_ASAP7_75t_L g5981 ( 
.A1(n_5648),
.A2(n_2807),
.B(n_5284),
.Y(n_5981)
);

CKINVDCx16_ASAP7_75t_R g5982 ( 
.A(n_5409),
.Y(n_5982)
);

OR2x4_ASAP7_75t_L g5983 ( 
.A(n_5463),
.B(n_1280),
.Y(n_5983)
);

NOR2xp33_ASAP7_75t_R g5984 ( 
.A(n_5554),
.B(n_5683),
.Y(n_5984)
);

INVx3_ASAP7_75t_L g5985 ( 
.A(n_5459),
.Y(n_5985)
);

NAND3xp33_ASAP7_75t_L g5986 ( 
.A(n_5448),
.B(n_1294),
.C(n_1280),
.Y(n_5986)
);

HB1xp67_ASAP7_75t_L g5987 ( 
.A(n_5586),
.Y(n_5987)
);

AND2x4_ASAP7_75t_L g5988 ( 
.A(n_5475),
.B(n_5284),
.Y(n_5988)
);

AOI221xp5_ASAP7_75t_L g5989 ( 
.A1(n_5682),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.C(n_38),
.Y(n_5989)
);

NAND2xp33_ASAP7_75t_SL g5990 ( 
.A(n_5673),
.B(n_34),
.Y(n_5990)
);

NAND2xp5_ASAP7_75t_L g5991 ( 
.A(n_5494),
.B(n_5367),
.Y(n_5991)
);

AOI21xp33_ASAP7_75t_L g5992 ( 
.A1(n_5560),
.A2(n_34),
.B(n_37),
.Y(n_5992)
);

INVx3_ASAP7_75t_L g5993 ( 
.A(n_5485),
.Y(n_5993)
);

AOI22xp33_ASAP7_75t_L g5994 ( 
.A1(n_5675),
.A2(n_1294),
.B1(n_1383),
.B2(n_1280),
.Y(n_5994)
);

OAI22xp5_ASAP7_75t_L g5995 ( 
.A1(n_5729),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_5995)
);

AOI22xp5_ASAP7_75t_L g5996 ( 
.A1(n_5672),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_5996)
);

AOI221xp5_ASAP7_75t_SL g5997 ( 
.A1(n_5460),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.C(n_44),
.Y(n_5997)
);

AOI22xp33_ASAP7_75t_L g5998 ( 
.A1(n_5678),
.A2(n_1294),
.B1(n_1432),
.B2(n_1383),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5570),
.Y(n_5999)
);

CKINVDCx11_ASAP7_75t_R g6000 ( 
.A(n_5683),
.Y(n_6000)
);

AOI22xp33_ASAP7_75t_L g6001 ( 
.A1(n_5544),
.A2(n_1294),
.B1(n_1432),
.B2(n_1383),
.Y(n_6001)
);

HB1xp67_ASAP7_75t_L g6002 ( 
.A(n_5588),
.Y(n_6002)
);

CKINVDCx5p33_ASAP7_75t_R g6003 ( 
.A(n_5690),
.Y(n_6003)
);

AND2x2_ASAP7_75t_L g6004 ( 
.A(n_5632),
.B(n_5369),
.Y(n_6004)
);

OAI22xp5_ASAP7_75t_L g6005 ( 
.A1(n_5463),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_6005)
);

CKINVDCx5p33_ASAP7_75t_R g6006 ( 
.A(n_5515),
.Y(n_6006)
);

AO21x2_ASAP7_75t_L g6007 ( 
.A1(n_5653),
.A2(n_5369),
.B(n_1293),
.Y(n_6007)
);

AND2x2_ASAP7_75t_L g6008 ( 
.A(n_5485),
.B(n_5522),
.Y(n_6008)
);

AOI22xp33_ASAP7_75t_L g6009 ( 
.A1(n_5544),
.A2(n_5601),
.B1(n_5622),
.B2(n_5672),
.Y(n_6009)
);

INVxp67_ASAP7_75t_L g6010 ( 
.A(n_5515),
.Y(n_6010)
);

NAND2xp5_ASAP7_75t_SL g6011 ( 
.A(n_5571),
.B(n_1294),
.Y(n_6011)
);

AND2x4_ASAP7_75t_L g6012 ( 
.A(n_5474),
.B(n_46),
.Y(n_6012)
);

NOR2x1_ASAP7_75t_L g6013 ( 
.A(n_5522),
.B(n_1383),
.Y(n_6013)
);

INVx2_ASAP7_75t_L g6014 ( 
.A(n_5590),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_5444),
.Y(n_6015)
);

INVx2_ASAP7_75t_SL g6016 ( 
.A(n_5455),
.Y(n_6016)
);

AND2x6_ASAP7_75t_L g6017 ( 
.A(n_5730),
.B(n_1383),
.Y(n_6017)
);

INVx2_ASAP7_75t_L g6018 ( 
.A(n_5530),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5539),
.Y(n_6019)
);

NAND2xp5_ASAP7_75t_L g6020 ( 
.A(n_5588),
.B(n_46),
.Y(n_6020)
);

INVx6_ASAP7_75t_L g6021 ( 
.A(n_5740),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5779),
.Y(n_6022)
);

CKINVDCx11_ASAP7_75t_R g6023 ( 
.A(n_5841),
.Y(n_6023)
);

CKINVDCx11_ASAP7_75t_R g6024 ( 
.A(n_5768),
.Y(n_6024)
);

A2O1A1Ixp33_ASAP7_75t_L g6025 ( 
.A1(n_5774),
.A2(n_5960),
.B(n_5810),
.C(n_5997),
.Y(n_6025)
);

AOI221xp5_ASAP7_75t_L g6026 ( 
.A1(n_5749),
.A2(n_5682),
.B1(n_5460),
.B2(n_5709),
.C(n_5676),
.Y(n_6026)
);

BUFx3_ASAP7_75t_L g6027 ( 
.A(n_5759),
.Y(n_6027)
);

OAI22xp5_ASAP7_75t_L g6028 ( 
.A1(n_5774),
.A2(n_5398),
.B1(n_5554),
.B2(n_5619),
.Y(n_6028)
);

AOI22xp33_ASAP7_75t_L g6029 ( 
.A1(n_5769),
.A2(n_5622),
.B1(n_5732),
.B2(n_5659),
.Y(n_6029)
);

NAND2xp5_ASAP7_75t_L g6030 ( 
.A(n_5924),
.B(n_5642),
.Y(n_6030)
);

OAI22xp5_ASAP7_75t_L g6031 ( 
.A1(n_5770),
.A2(n_5619),
.B1(n_5721),
.B2(n_5552),
.Y(n_6031)
);

OAI211xp5_ASAP7_75t_SL g6032 ( 
.A1(n_5797),
.A2(n_5456),
.B(n_5556),
.C(n_5676),
.Y(n_6032)
);

AOI22xp33_ASAP7_75t_L g6033 ( 
.A1(n_5946),
.A2(n_5732),
.B1(n_5653),
.B2(n_5667),
.Y(n_6033)
);

HB1xp67_ASAP7_75t_L g6034 ( 
.A(n_5750),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_5894),
.B(n_5642),
.Y(n_6035)
);

HB1xp67_ASAP7_75t_L g6036 ( 
.A(n_5772),
.Y(n_6036)
);

AOI22xp33_ASAP7_75t_L g6037 ( 
.A1(n_5958),
.A2(n_5659),
.B1(n_5667),
.B2(n_5525),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_5804),
.Y(n_6038)
);

CKINVDCx20_ASAP7_75t_R g6039 ( 
.A(n_6000),
.Y(n_6039)
);

OA21x2_ASAP7_75t_L g6040 ( 
.A1(n_5847),
.A2(n_5707),
.B(n_5684),
.Y(n_6040)
);

AOI22xp5_ASAP7_75t_L g6041 ( 
.A1(n_5814),
.A2(n_5997),
.B1(n_5742),
.B2(n_5806),
.Y(n_6041)
);

AOI22xp33_ASAP7_75t_SL g6042 ( 
.A1(n_5834),
.A2(n_5578),
.B1(n_5519),
.B2(n_5688),
.Y(n_6042)
);

AND2x4_ASAP7_75t_L g6043 ( 
.A(n_5756),
.B(n_5828),
.Y(n_6043)
);

AOI22xp5_ASAP7_75t_L g6044 ( 
.A1(n_5942),
.A2(n_5688),
.B1(n_5456),
.B2(n_5709),
.Y(n_6044)
);

INVx2_ASAP7_75t_L g6045 ( 
.A(n_5780),
.Y(n_6045)
);

AOI21xp5_ASAP7_75t_L g6046 ( 
.A1(n_5986),
.A2(n_5648),
.B(n_5448),
.Y(n_6046)
);

BUFx2_ASAP7_75t_L g6047 ( 
.A(n_5984),
.Y(n_6047)
);

OAI221xp5_ASAP7_75t_L g6048 ( 
.A1(n_5911),
.A2(n_5658),
.B1(n_5470),
.B2(n_5719),
.C(n_5731),
.Y(n_6048)
);

AOI221xp5_ASAP7_75t_L g6049 ( 
.A1(n_5891),
.A2(n_5719),
.B1(n_5608),
.B2(n_5658),
.C(n_5731),
.Y(n_6049)
);

AOI21xp5_ASAP7_75t_L g6050 ( 
.A1(n_5986),
.A2(n_5621),
.B(n_5704),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_5815),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5822),
.Y(n_6052)
);

OAI22xp5_ASAP7_75t_L g6053 ( 
.A1(n_6009),
.A2(n_5721),
.B1(n_5668),
.B2(n_5730),
.Y(n_6053)
);

AND2x4_ASAP7_75t_L g6054 ( 
.A(n_5756),
.B(n_5474),
.Y(n_6054)
);

AOI22xp33_ASAP7_75t_L g6055 ( 
.A1(n_5898),
.A2(n_5892),
.B1(n_5746),
.B2(n_5743),
.Y(n_6055)
);

NAND2xp5_ASAP7_75t_L g6056 ( 
.A(n_5900),
.B(n_5444),
.Y(n_6056)
);

NAND2xp5_ASAP7_75t_L g6057 ( 
.A(n_5910),
.B(n_5685),
.Y(n_6057)
);

NAND2xp5_ASAP7_75t_L g6058 ( 
.A(n_5755),
.B(n_5685),
.Y(n_6058)
);

OAI222xp33_ASAP7_75t_L g6059 ( 
.A1(n_5839),
.A2(n_5666),
.B1(n_5665),
.B2(n_5614),
.C1(n_5587),
.C2(n_5616),
.Y(n_6059)
);

INVx2_ASAP7_75t_L g6060 ( 
.A(n_5969),
.Y(n_6060)
);

OAI21xp5_ASAP7_75t_L g6061 ( 
.A1(n_5916),
.A2(n_5857),
.B(n_5784),
.Y(n_6061)
);

INVx3_ASAP7_75t_L g6062 ( 
.A(n_5762),
.Y(n_6062)
);

INVx3_ASAP7_75t_L g6063 ( 
.A(n_5762),
.Y(n_6063)
);

AOI22xp5_ASAP7_75t_L g6064 ( 
.A1(n_5751),
.A2(n_5609),
.B1(n_5608),
.B2(n_5674),
.Y(n_6064)
);

AO21x2_ASAP7_75t_L g6065 ( 
.A1(n_6015),
.A2(n_5867),
.B(n_5938),
.Y(n_6065)
);

INVx2_ASAP7_75t_L g6066 ( 
.A(n_5932),
.Y(n_6066)
);

AND2x4_ASAP7_75t_L g6067 ( 
.A(n_5790),
.B(n_5730),
.Y(n_6067)
);

A2O1A1Ixp33_ASAP7_75t_L g6068 ( 
.A1(n_5888),
.A2(n_5434),
.B(n_5714),
.C(n_5710),
.Y(n_6068)
);

AOI222xp33_ASAP7_75t_L g6069 ( 
.A1(n_5989),
.A2(n_5656),
.B1(n_5733),
.B2(n_5698),
.C1(n_5674),
.C2(n_5603),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5870),
.Y(n_6070)
);

BUFx6f_ASAP7_75t_L g6071 ( 
.A(n_5762),
.Y(n_6071)
);

AND2x2_ASAP7_75t_SL g6072 ( 
.A(n_6012),
.B(n_5390),
.Y(n_6072)
);

OR2x6_ASAP7_75t_L g6073 ( 
.A(n_5790),
.B(n_5584),
.Y(n_6073)
);

OAI22xp5_ASAP7_75t_L g6074 ( 
.A1(n_5767),
.A2(n_5668),
.B1(n_5621),
.B2(n_5556),
.Y(n_6074)
);

AO31x2_ASAP7_75t_L g6075 ( 
.A1(n_5781),
.A2(n_5845),
.A3(n_5811),
.B(n_5962),
.Y(n_6075)
);

INVxp67_ASAP7_75t_L g6076 ( 
.A(n_5738),
.Y(n_6076)
);

AOI21xp5_ASAP7_75t_L g6077 ( 
.A1(n_5766),
.A2(n_5505),
.B(n_5650),
.Y(n_6077)
);

OA21x2_ASAP7_75t_L g6078 ( 
.A1(n_5876),
.A2(n_5513),
.B(n_5473),
.Y(n_6078)
);

CKINVDCx11_ASAP7_75t_R g6079 ( 
.A(n_5785),
.Y(n_6079)
);

OAI21x1_ASAP7_75t_L g6080 ( 
.A1(n_5789),
.A2(n_5388),
.B(n_5563),
.Y(n_6080)
);

INVx2_ASAP7_75t_L g6081 ( 
.A(n_5873),
.Y(n_6081)
);

INVx3_ASAP7_75t_L g6082 ( 
.A(n_5740),
.Y(n_6082)
);

AOI21xp5_ASAP7_75t_L g6083 ( 
.A1(n_5760),
.A2(n_5650),
.B(n_5426),
.Y(n_6083)
);

NAND2xp5_ASAP7_75t_L g6084 ( 
.A(n_5764),
.B(n_5533),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_L g6085 ( 
.A(n_5909),
.B(n_5915),
.Y(n_6085)
);

OAI22xp5_ASAP7_75t_L g6086 ( 
.A1(n_5890),
.A2(n_5954),
.B1(n_5982),
.B2(n_5966),
.Y(n_6086)
);

OA21x2_ASAP7_75t_L g6087 ( 
.A1(n_5741),
.A2(n_5466),
.B(n_5389),
.Y(n_6087)
);

BUFx2_ASAP7_75t_L g6088 ( 
.A(n_5782),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5906),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5907),
.Y(n_6090)
);

AOI22xp5_ASAP7_75t_L g6091 ( 
.A1(n_5904),
.A2(n_5609),
.B1(n_5698),
.B2(n_5660),
.Y(n_6091)
);

OR2x2_ASAP7_75t_L g6092 ( 
.A(n_5739),
.B(n_5440),
.Y(n_6092)
);

OAI221xp5_ASAP7_75t_L g6093 ( 
.A1(n_5951),
.A2(n_5434),
.B1(n_5612),
.B2(n_5440),
.C(n_5567),
.Y(n_6093)
);

AOI22xp33_ASAP7_75t_L g6094 ( 
.A1(n_5834),
.A2(n_5525),
.B1(n_5700),
.B2(n_5655),
.Y(n_6094)
);

AOI22xp5_ASAP7_75t_L g6095 ( 
.A1(n_5773),
.A2(n_5660),
.B1(n_5636),
.B2(n_5519),
.Y(n_6095)
);

OAI22xp5_ASAP7_75t_L g6096 ( 
.A1(n_5837),
.A2(n_5893),
.B1(n_5843),
.B2(n_5821),
.Y(n_6096)
);

CKINVDCx11_ASAP7_75t_R g6097 ( 
.A(n_5736),
.Y(n_6097)
);

AOI22xp33_ASAP7_75t_L g6098 ( 
.A1(n_5758),
.A2(n_5700),
.B1(n_5655),
.B2(n_5733),
.Y(n_6098)
);

NAND2xp5_ASAP7_75t_L g6099 ( 
.A(n_5918),
.B(n_5447),
.Y(n_6099)
);

AOI21xp5_ASAP7_75t_L g6100 ( 
.A1(n_5796),
.A2(n_5518),
.B(n_5640),
.Y(n_6100)
);

OAI21xp5_ASAP7_75t_L g6101 ( 
.A1(n_5821),
.A2(n_5445),
.B(n_5500),
.Y(n_6101)
);

BUFx6f_ASAP7_75t_L g6102 ( 
.A(n_5818),
.Y(n_6102)
);

CKINVDCx8_ASAP7_75t_R g6103 ( 
.A(n_5968),
.Y(n_6103)
);

NAND2xp5_ASAP7_75t_L g6104 ( 
.A(n_5959),
.B(n_5458),
.Y(n_6104)
);

AOI22xp33_ASAP7_75t_SL g6105 ( 
.A1(n_5754),
.A2(n_5519),
.B1(n_5469),
.B2(n_5458),
.Y(n_6105)
);

AOI22xp33_ASAP7_75t_L g6106 ( 
.A1(n_5763),
.A2(n_5733),
.B1(n_5543),
.B2(n_5469),
.Y(n_6106)
);

AOI22xp33_ASAP7_75t_L g6107 ( 
.A1(n_5819),
.A2(n_5543),
.B1(n_5566),
.B2(n_5534),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_5913),
.Y(n_6108)
);

AO21x2_ASAP7_75t_L g6109 ( 
.A1(n_5972),
.A2(n_5643),
.B(n_5569),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_5775),
.Y(n_6110)
);

A2O1A1Ixp33_ASAP7_75t_L g6111 ( 
.A1(n_5996),
.A2(n_5636),
.B(n_5536),
.C(n_5477),
.Y(n_6111)
);

NAND2xp5_ASAP7_75t_L g6112 ( 
.A(n_6002),
.B(n_5702),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_5936),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_5783),
.Y(n_6114)
);

AOI22xp33_ASAP7_75t_L g6115 ( 
.A1(n_5889),
.A2(n_5566),
.B1(n_5534),
.B2(n_5611),
.Y(n_6115)
);

OAI22xp33_ASAP7_75t_L g6116 ( 
.A1(n_5761),
.A2(n_5584),
.B1(n_5595),
.B2(n_5620),
.Y(n_6116)
);

AND2x2_ASAP7_75t_L g6117 ( 
.A(n_5787),
.B(n_5518),
.Y(n_6117)
);

NAND3xp33_ASAP7_75t_L g6118 ( 
.A(n_5765),
.B(n_5718),
.C(n_5708),
.Y(n_6118)
);

AOI222xp33_ASAP7_75t_L g6119 ( 
.A1(n_5777),
.A2(n_5468),
.B1(n_5519),
.B2(n_5702),
.C1(n_5664),
.C2(n_5497),
.Y(n_6119)
);

OAI221xp5_ASAP7_75t_L g6120 ( 
.A1(n_5996),
.A2(n_5620),
.B1(n_5595),
.B2(n_5713),
.C(n_5582),
.Y(n_6120)
);

INVx1_ASAP7_75t_L g6121 ( 
.A(n_5792),
.Y(n_6121)
);

INVx4_ASAP7_75t_L g6122 ( 
.A(n_5740),
.Y(n_6122)
);

NAND2xp5_ASAP7_75t_L g6123 ( 
.A(n_5744),
.B(n_5745),
.Y(n_6123)
);

AOI22xp33_ASAP7_75t_L g6124 ( 
.A1(n_5889),
.A2(n_5829),
.B1(n_5853),
.B2(n_5801),
.Y(n_6124)
);

AOI221xp5_ASAP7_75t_L g6125 ( 
.A1(n_6005),
.A2(n_5713),
.B1(n_49),
.B2(n_47),
.C(n_48),
.Y(n_6125)
);

NAND2xp5_ASAP7_75t_L g6126 ( 
.A(n_5748),
.B(n_5640),
.Y(n_6126)
);

OAI22xp5_ASAP7_75t_L g6127 ( 
.A1(n_6010),
.A2(n_5638),
.B1(n_5645),
.B2(n_5686),
.Y(n_6127)
);

AOI221xp5_ASAP7_75t_L g6128 ( 
.A1(n_5995),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_6128)
);

AND2x4_ASAP7_75t_L g6129 ( 
.A(n_5790),
.B(n_5645),
.Y(n_6129)
);

OAI22xp5_ASAP7_75t_L g6130 ( 
.A1(n_6012),
.A2(n_5638),
.B1(n_5686),
.B2(n_5697),
.Y(n_6130)
);

OA21x2_ASAP7_75t_L g6131 ( 
.A1(n_5920),
.A2(n_5496),
.B(n_5610),
.Y(n_6131)
);

AOI22xp33_ASAP7_75t_L g6132 ( 
.A1(n_5803),
.A2(n_5611),
.B1(n_5519),
.B2(n_5596),
.Y(n_6132)
);

AND2x2_ASAP7_75t_L g6133 ( 
.A(n_5787),
.B(n_5638),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_5903),
.Y(n_6134)
);

INVx2_ASAP7_75t_L g6135 ( 
.A(n_5927),
.Y(n_6135)
);

OAI22xp5_ASAP7_75t_L g6136 ( 
.A1(n_5944),
.A2(n_5584),
.B1(n_5689),
.B2(n_5699),
.Y(n_6136)
);

INVx2_ASAP7_75t_L g6137 ( 
.A(n_5869),
.Y(n_6137)
);

O2A1O1Ixp33_ASAP7_75t_L g6138 ( 
.A1(n_5795),
.A2(n_5689),
.B(n_5594),
.C(n_5582),
.Y(n_6138)
);

OAI221xp5_ASAP7_75t_L g6139 ( 
.A1(n_5872),
.A2(n_5965),
.B1(n_5897),
.B2(n_5830),
.C(n_5855),
.Y(n_6139)
);

HB1xp67_ASAP7_75t_L g6140 ( 
.A(n_5753),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5859),
.Y(n_6141)
);

AOI22xp5_ASAP7_75t_L g6142 ( 
.A1(n_5832),
.A2(n_5670),
.B1(n_5596),
.B2(n_5605),
.Y(n_6142)
);

NAND2xp5_ASAP7_75t_L g6143 ( 
.A(n_5856),
.B(n_5701),
.Y(n_6143)
);

AOI22xp5_ASAP7_75t_L g6144 ( 
.A1(n_5947),
.A2(n_5596),
.B1(n_5605),
.B2(n_5497),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_5860),
.Y(n_6145)
);

AOI21xp5_ASAP7_75t_L g6146 ( 
.A1(n_5788),
.A2(n_5722),
.B(n_5594),
.Y(n_6146)
);

OAI211xp5_ASAP7_75t_L g6147 ( 
.A1(n_5807),
.A2(n_5712),
.B(n_5559),
.C(n_5492),
.Y(n_6147)
);

AOI21xp5_ASAP7_75t_L g6148 ( 
.A1(n_5761),
.A2(n_5407),
.B(n_5497),
.Y(n_6148)
);

OAI22xp5_ASAP7_75t_SL g6149 ( 
.A1(n_5970),
.A2(n_5925),
.B1(n_5937),
.B2(n_5840),
.Y(n_6149)
);

AOI21xp5_ASAP7_75t_L g6150 ( 
.A1(n_5761),
.A2(n_5407),
.B(n_5605),
.Y(n_6150)
);

OAI211xp5_ASAP7_75t_L g6151 ( 
.A1(n_5896),
.A2(n_5712),
.B(n_5407),
.C(n_5727),
.Y(n_6151)
);

AOI21xp5_ASAP7_75t_L g6152 ( 
.A1(n_5757),
.A2(n_5699),
.B(n_5502),
.Y(n_6152)
);

OR2x2_ASAP7_75t_L g6153 ( 
.A(n_5987),
.B(n_5734),
.Y(n_6153)
);

NAND2x1p5_ASAP7_75t_L g6154 ( 
.A(n_5802),
.B(n_5662),
.Y(n_6154)
);

OR2x6_ASAP7_75t_L g6155 ( 
.A(n_5864),
.B(n_5493),
.Y(n_6155)
);

OAI221xp5_ASAP7_75t_L g6156 ( 
.A1(n_5849),
.A2(n_5691),
.B1(n_5734),
.B2(n_5644),
.C(n_1488),
.Y(n_6156)
);

AOI22xp33_ASAP7_75t_L g6157 ( 
.A1(n_5826),
.A2(n_5495),
.B1(n_5478),
.B2(n_5528),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5863),
.Y(n_6158)
);

INVx2_ASAP7_75t_L g6159 ( 
.A(n_5861),
.Y(n_6159)
);

AOI21xp5_ASAP7_75t_L g6160 ( 
.A1(n_5983),
.A2(n_5482),
.B(n_5592),
.Y(n_6160)
);

CKINVDCx11_ASAP7_75t_R g6161 ( 
.A(n_5846),
.Y(n_6161)
);

AOI22xp33_ASAP7_75t_L g6162 ( 
.A1(n_5826),
.A2(n_5568),
.B1(n_5511),
.B2(n_5615),
.Y(n_6162)
);

OAI33xp33_ASAP7_75t_L g6163 ( 
.A1(n_6020),
.A2(n_52),
.A3(n_54),
.B1(n_48),
.B2(n_49),
.B3(n_53),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_5880),
.Y(n_6164)
);

INVx2_ASAP7_75t_L g6165 ( 
.A(n_5875),
.Y(n_6165)
);

AOI221xp5_ASAP7_75t_L g6166 ( 
.A1(n_5808),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.C(n_55),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_5886),
.Y(n_6167)
);

AND2x2_ASAP7_75t_L g6168 ( 
.A(n_5862),
.B(n_5695),
.Y(n_6168)
);

OR2x6_ASAP7_75t_L g6169 ( 
.A(n_5805),
.B(n_5687),
.Y(n_6169)
);

AOI221xp5_ASAP7_75t_L g6170 ( 
.A1(n_5800),
.A2(n_5825),
.B1(n_5978),
.B2(n_5992),
.C(n_5899),
.Y(n_6170)
);

AOI22xp33_ASAP7_75t_L g6171 ( 
.A1(n_5844),
.A2(n_5503),
.B1(n_5711),
.B2(n_5535),
.Y(n_6171)
);

OAI221xp5_ASAP7_75t_L g6172 ( 
.A1(n_5945),
.A2(n_5734),
.B1(n_5644),
.B2(n_1488),
.C(n_1463),
.Y(n_6172)
);

AOI22xp33_ASAP7_75t_L g6173 ( 
.A1(n_5844),
.A2(n_5647),
.B1(n_5623),
.B2(n_5637),
.Y(n_6173)
);

AOI22xp33_ASAP7_75t_SL g6174 ( 
.A1(n_5816),
.A2(n_5694),
.B1(n_5734),
.B2(n_5644),
.Y(n_6174)
);

INVx3_ASAP7_75t_L g6175 ( 
.A(n_5842),
.Y(n_6175)
);

INVx2_ASAP7_75t_L g6176 ( 
.A(n_5771),
.Y(n_6176)
);

AOI221xp5_ASAP7_75t_L g6177 ( 
.A1(n_5899),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.C(n_56),
.Y(n_6177)
);

OR2x2_ASAP7_75t_L g6178 ( 
.A(n_5963),
.B(n_5896),
.Y(n_6178)
);

AOI21xp5_ASAP7_75t_L g6179 ( 
.A1(n_6011),
.A2(n_5726),
.B(n_5725),
.Y(n_6179)
);

AND2x4_ASAP7_75t_L g6180 ( 
.A(n_5823),
.B(n_5703),
.Y(n_6180)
);

AOI21xp5_ASAP7_75t_L g6181 ( 
.A1(n_5823),
.A2(n_5549),
.B(n_5542),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_5964),
.Y(n_6182)
);

OA21x2_ASAP7_75t_L g6183 ( 
.A1(n_5930),
.A2(n_5624),
.B(n_5669),
.Y(n_6183)
);

NOR2x1_ASAP7_75t_SL g6184 ( 
.A(n_5802),
.B(n_5644),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_5778),
.Y(n_6185)
);

CKINVDCx20_ASAP7_75t_R g6186 ( 
.A(n_5817),
.Y(n_6186)
);

AND2x2_ASAP7_75t_L g6187 ( 
.A(n_6008),
.B(n_5520),
.Y(n_6187)
);

OA21x2_ASAP7_75t_L g6188 ( 
.A1(n_5865),
.A2(n_5527),
.B(n_5529),
.Y(n_6188)
);

AOI21xp5_ASAP7_75t_L g6189 ( 
.A1(n_5823),
.A2(n_1463),
.B(n_1432),
.Y(n_6189)
);

AND2x2_ASAP7_75t_L g6190 ( 
.A(n_5794),
.B(n_55),
.Y(n_6190)
);

OAI22xp5_ASAP7_75t_L g6191 ( 
.A1(n_5944),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_6191)
);

AOI221xp5_ASAP7_75t_L g6192 ( 
.A1(n_5833),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_6192)
);

AOI21xp5_ASAP7_75t_L g6193 ( 
.A1(n_5809),
.A2(n_1463),
.B(n_1432),
.Y(n_6193)
);

OR2x2_ASAP7_75t_L g6194 ( 
.A(n_5776),
.B(n_57),
.Y(n_6194)
);

AOI22xp33_ASAP7_75t_L g6195 ( 
.A1(n_6004),
.A2(n_1463),
.B1(n_1488),
.B2(n_1432),
.Y(n_6195)
);

AND2x2_ASAP7_75t_L g6196 ( 
.A(n_6016),
.B(n_59),
.Y(n_6196)
);

AND2x2_ASAP7_75t_L g6197 ( 
.A(n_5831),
.B(n_60),
.Y(n_6197)
);

AOI22xp33_ASAP7_75t_L g6198 ( 
.A1(n_5813),
.A2(n_1488),
.B1(n_1463),
.B2(n_2141),
.Y(n_6198)
);

AOI22xp33_ASAP7_75t_L g6199 ( 
.A1(n_5948),
.A2(n_5866),
.B1(n_5858),
.B2(n_5988),
.Y(n_6199)
);

AOI22xp33_ASAP7_75t_L g6200 ( 
.A1(n_5858),
.A2(n_1488),
.B1(n_2142),
.B2(n_2141),
.Y(n_6200)
);

NAND2xp5_ASAP7_75t_L g6201 ( 
.A(n_5786),
.B(n_165),
.Y(n_6201)
);

OA21x2_ASAP7_75t_L g6202 ( 
.A1(n_5879),
.A2(n_1303),
.B(n_1302),
.Y(n_6202)
);

INVx3_ASAP7_75t_L g6203 ( 
.A(n_5842),
.Y(n_6203)
);

AOI22xp33_ASAP7_75t_SL g6204 ( 
.A1(n_5988),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_6204)
);

OA21x2_ASAP7_75t_L g6205 ( 
.A1(n_5882),
.A2(n_1305),
.B(n_1303),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5949),
.Y(n_6206)
);

AOI221xp5_ASAP7_75t_L g6207 ( 
.A1(n_5955),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.C(n_66),
.Y(n_6207)
);

AND2x2_ASAP7_75t_L g6208 ( 
.A(n_5850),
.B(n_62),
.Y(n_6208)
);

INVx2_ASAP7_75t_SL g6209 ( 
.A(n_5782),
.Y(n_6209)
);

AOI22xp33_ASAP7_75t_L g6210 ( 
.A1(n_5827),
.A2(n_2142),
.B1(n_2143),
.B2(n_1307),
.Y(n_6210)
);

INVxp67_ASAP7_75t_L g6211 ( 
.A(n_5737),
.Y(n_6211)
);

AOI21xp5_ASAP7_75t_L g6212 ( 
.A1(n_6013),
.A2(n_63),
.B(n_64),
.Y(n_6212)
);

INVx1_ASAP7_75t_SL g6213 ( 
.A(n_5922),
.Y(n_6213)
);

OAI22xp5_ASAP7_75t_L g6214 ( 
.A1(n_6006),
.A2(n_67),
.B1(n_63),
.B2(n_66),
.Y(n_6214)
);

BUFx12f_ASAP7_75t_L g6215 ( 
.A(n_5933),
.Y(n_6215)
);

AND2x2_ASAP7_75t_L g6216 ( 
.A(n_5793),
.B(n_67),
.Y(n_6216)
);

OA21x2_ASAP7_75t_L g6217 ( 
.A1(n_5887),
.A2(n_1307),
.B(n_1305),
.Y(n_6217)
);

CKINVDCx5p33_ASAP7_75t_R g6218 ( 
.A(n_5791),
.Y(n_6218)
);

OAI22xp5_ASAP7_75t_L g6219 ( 
.A1(n_5950),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_6219)
);

AND2x4_ASAP7_75t_L g6220 ( 
.A(n_5935),
.B(n_70),
.Y(n_6220)
);

OAI21x1_ASAP7_75t_L g6221 ( 
.A1(n_5979),
.A2(n_70),
.B(n_71),
.Y(n_6221)
);

OAI221xp5_ASAP7_75t_L g6222 ( 
.A1(n_5957),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.C(n_75),
.Y(n_6222)
);

NAND2xp5_ASAP7_75t_L g6223 ( 
.A(n_5975),
.B(n_165),
.Y(n_6223)
);

AND2x2_ASAP7_75t_L g6224 ( 
.A(n_5793),
.B(n_71),
.Y(n_6224)
);

HB1xp67_ASAP7_75t_L g6225 ( 
.A(n_5883),
.Y(n_6225)
);

AOI21xp5_ASAP7_75t_L g6226 ( 
.A1(n_6013),
.A2(n_72),
.B(n_73),
.Y(n_6226)
);

AOI22xp33_ASAP7_75t_L g6227 ( 
.A1(n_5851),
.A2(n_2142),
.B1(n_2143),
.B2(n_1311),
.Y(n_6227)
);

OAI21x1_ASAP7_75t_L g6228 ( 
.A1(n_5883),
.A2(n_5980),
.B(n_5901),
.Y(n_6228)
);

AND2x2_ASAP7_75t_L g6229 ( 
.A(n_5985),
.B(n_72),
.Y(n_6229)
);

NAND2xp5_ASAP7_75t_L g6230 ( 
.A(n_5985),
.B(n_166),
.Y(n_6230)
);

AND2x2_ASAP7_75t_L g6231 ( 
.A(n_5993),
.B(n_75),
.Y(n_6231)
);

AND2x4_ASAP7_75t_L g6232 ( 
.A(n_5935),
.B(n_76),
.Y(n_6232)
);

INVx3_ASAP7_75t_L g6233 ( 
.A(n_5901),
.Y(n_6233)
);

AOI22xp33_ASAP7_75t_L g6234 ( 
.A1(n_5799),
.A2(n_2142),
.B1(n_2143),
.B2(n_1311),
.Y(n_6234)
);

INVx5_ASAP7_75t_L g6235 ( 
.A(n_5818),
.Y(n_6235)
);

AO21x2_ASAP7_75t_L g6236 ( 
.A1(n_5931),
.A2(n_76),
.B(n_77),
.Y(n_6236)
);

AOI221xp5_ASAP7_75t_L g6237 ( 
.A1(n_5919),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.C(n_80),
.Y(n_6237)
);

NAND3xp33_ASAP7_75t_L g6238 ( 
.A(n_5820),
.B(n_78),
.C(n_79),
.Y(n_6238)
);

AND2x2_ASAP7_75t_L g6239 ( 
.A(n_5993),
.B(n_80),
.Y(n_6239)
);

OAI22xp5_ASAP7_75t_L g6240 ( 
.A1(n_5747),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_6240)
);

NAND2x1_ASAP7_75t_L g6241 ( 
.A(n_5980),
.B(n_5824),
.Y(n_6241)
);

OAI22xp33_ASAP7_75t_L g6242 ( 
.A1(n_5848),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_5991),
.Y(n_6243)
);

AND2x2_ASAP7_75t_L g6244 ( 
.A(n_5871),
.B(n_6003),
.Y(n_6244)
);

AOI22xp33_ASAP7_75t_L g6245 ( 
.A1(n_5941),
.A2(n_2142),
.B1(n_2143),
.B2(n_1313),
.Y(n_6245)
);

OAI221xp5_ASAP7_75t_L g6246 ( 
.A1(n_5990),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.C(n_86),
.Y(n_6246)
);

NAND2xp5_ASAP7_75t_L g6247 ( 
.A(n_5852),
.B(n_5798),
.Y(n_6247)
);

OA21x2_ASAP7_75t_L g6248 ( 
.A1(n_5905),
.A2(n_1313),
.B(n_1309),
.Y(n_6248)
);

AOI22xp33_ASAP7_75t_SL g6249 ( 
.A1(n_5877),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_6249)
);

HB1xp67_ASAP7_75t_L g6250 ( 
.A(n_5854),
.Y(n_6250)
);

OAI21x1_ASAP7_75t_L g6251 ( 
.A1(n_5914),
.A2(n_84),
.B(n_85),
.Y(n_6251)
);

OAI221xp5_ASAP7_75t_L g6252 ( 
.A1(n_5877),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.C(n_89),
.Y(n_6252)
);

AOI22xp33_ASAP7_75t_L g6253 ( 
.A1(n_6018),
.A2(n_6019),
.B1(n_5921),
.B2(n_5895),
.Y(n_6253)
);

AOI22xp33_ASAP7_75t_L g6254 ( 
.A1(n_5921),
.A2(n_2143),
.B1(n_1314),
.B2(n_1317),
.Y(n_6254)
);

AOI22xp33_ASAP7_75t_L g6255 ( 
.A1(n_5878),
.A2(n_2143),
.B1(n_1314),
.B2(n_1317),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5967),
.Y(n_6256)
);

AOI21x1_ASAP7_75t_L g6257 ( 
.A1(n_5934),
.A2(n_5874),
.B(n_5939),
.Y(n_6257)
);

BUFx4f_ASAP7_75t_SL g6258 ( 
.A(n_5836),
.Y(n_6258)
);

BUFx4f_ASAP7_75t_SL g6259 ( 
.A(n_5818),
.Y(n_6259)
);

AOI22xp33_ASAP7_75t_L g6260 ( 
.A1(n_5971),
.A2(n_1318),
.B1(n_1320),
.B2(n_1309),
.Y(n_6260)
);

AOI221xp5_ASAP7_75t_L g6261 ( 
.A1(n_5977),
.A2(n_91),
.B1(n_88),
.B2(n_90),
.C(n_92),
.Y(n_6261)
);

OR2x2_ASAP7_75t_L g6262 ( 
.A(n_5752),
.B(n_5939),
.Y(n_6262)
);

AND2x2_ASAP7_75t_L g6263 ( 
.A(n_5802),
.B(n_88),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_5976),
.Y(n_6264)
);

AOI22xp33_ASAP7_75t_SL g6265 ( 
.A1(n_5952),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_6265)
);

OAI211xp5_ASAP7_75t_SL g6266 ( 
.A1(n_5974),
.A2(n_94),
.B(n_90),
.C(n_93),
.Y(n_6266)
);

OAI22xp33_ASAP7_75t_L g6267 ( 
.A1(n_5848),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_6267)
);

AOI211xp5_ASAP7_75t_L g6268 ( 
.A1(n_5884),
.A2(n_98),
.B(n_94),
.C(n_97),
.Y(n_6268)
);

AOI21xp5_ASAP7_75t_L g6269 ( 
.A1(n_5848),
.A2(n_98),
.B(n_99),
.Y(n_6269)
);

AOI22xp33_ASAP7_75t_SL g6270 ( 
.A1(n_5952),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_6270)
);

OAI22xp33_ASAP7_75t_L g6271 ( 
.A1(n_5868),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_6271)
);

BUFx3_ASAP7_75t_L g6272 ( 
.A(n_5824),
.Y(n_6272)
);

NAND2xp5_ASAP7_75t_L g6273 ( 
.A(n_5902),
.B(n_166),
.Y(n_6273)
);

NOR2xp33_ASAP7_75t_R g6274 ( 
.A(n_6039),
.B(n_5902),
.Y(n_6274)
);

NAND2xp33_ASAP7_75t_R g6275 ( 
.A(n_6047),
.B(n_5868),
.Y(n_6275)
);

XNOR2xp5_ASAP7_75t_L g6276 ( 
.A(n_6041),
.B(n_5923),
.Y(n_6276)
);

AND2x2_ASAP7_75t_L g6277 ( 
.A(n_6117),
.B(n_5902),
.Y(n_6277)
);

AND2x4_ASAP7_75t_L g6278 ( 
.A(n_6088),
.B(n_5908),
.Y(n_6278)
);

NOR2xp33_ASAP7_75t_R g6279 ( 
.A(n_6161),
.B(n_5908),
.Y(n_6279)
);

AND2x4_ASAP7_75t_L g6280 ( 
.A(n_6175),
.B(n_6203),
.Y(n_6280)
);

AND2x2_ASAP7_75t_L g6281 ( 
.A(n_6133),
.B(n_5908),
.Y(n_6281)
);

OR2x6_ASAP7_75t_L g6282 ( 
.A(n_6021),
.B(n_5805),
.Y(n_6282)
);

NOR2xp33_ASAP7_75t_R g6283 ( 
.A(n_6186),
.B(n_101),
.Y(n_6283)
);

HB1xp67_ASAP7_75t_L g6284 ( 
.A(n_6034),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_6051),
.Y(n_6285)
);

INVxp67_ASAP7_75t_L g6286 ( 
.A(n_6250),
.Y(n_6286)
);

BUFx3_ASAP7_75t_L g6287 ( 
.A(n_6024),
.Y(n_6287)
);

XOR2xp5_ASAP7_75t_L g6288 ( 
.A(n_6041),
.B(n_5926),
.Y(n_6288)
);

INVx2_ASAP7_75t_SL g6289 ( 
.A(n_6027),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_6087),
.Y(n_6290)
);

AND2x4_ASAP7_75t_L g6291 ( 
.A(n_6175),
.B(n_5805),
.Y(n_6291)
);

BUFx3_ASAP7_75t_L g6292 ( 
.A(n_6023),
.Y(n_6292)
);

CKINVDCx8_ASAP7_75t_R g6293 ( 
.A(n_6218),
.Y(n_6293)
);

CKINVDCx8_ASAP7_75t_R g6294 ( 
.A(n_6235),
.Y(n_6294)
);

AND2x4_ASAP7_75t_L g6295 ( 
.A(n_6203),
.B(n_5934),
.Y(n_6295)
);

NOR2xp33_ASAP7_75t_R g6296 ( 
.A(n_6097),
.B(n_101),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_6052),
.Y(n_6297)
);

CKINVDCx8_ASAP7_75t_R g6298 ( 
.A(n_6235),
.Y(n_6298)
);

AND2x4_ASAP7_75t_L g6299 ( 
.A(n_6043),
.B(n_5868),
.Y(n_6299)
);

AND2x2_ASAP7_75t_L g6300 ( 
.A(n_6062),
.B(n_5973),
.Y(n_6300)
);

NAND2xp5_ASAP7_75t_L g6301 ( 
.A(n_6025),
.B(n_6190),
.Y(n_6301)
);

NAND2xp5_ASAP7_75t_L g6302 ( 
.A(n_6038),
.B(n_5981),
.Y(n_6302)
);

AND2x2_ASAP7_75t_L g6303 ( 
.A(n_6062),
.B(n_5812),
.Y(n_6303)
);

NAND2xp5_ASAP7_75t_SL g6304 ( 
.A(n_6043),
.B(n_5929),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6089),
.Y(n_6305)
);

OR2x6_ASAP7_75t_L g6306 ( 
.A(n_6021),
.B(n_5838),
.Y(n_6306)
);

AND2x2_ASAP7_75t_L g6307 ( 
.A(n_6063),
.B(n_5881),
.Y(n_6307)
);

NAND2xp5_ASAP7_75t_L g6308 ( 
.A(n_6194),
.B(n_5956),
.Y(n_6308)
);

NAND2xp33_ASAP7_75t_R g6309 ( 
.A(n_6061),
.B(n_102),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_6090),
.Y(n_6310)
);

INVxp67_ASAP7_75t_L g6311 ( 
.A(n_6086),
.Y(n_6311)
);

NOR2xp33_ASAP7_75t_R g6312 ( 
.A(n_6079),
.B(n_102),
.Y(n_6312)
);

CKINVDCx8_ASAP7_75t_R g6313 ( 
.A(n_6235),
.Y(n_6313)
);

XNOR2xp5_ASAP7_75t_L g6314 ( 
.A(n_6072),
.B(n_5928),
.Y(n_6314)
);

AND2x2_ASAP7_75t_L g6315 ( 
.A(n_6063),
.B(n_5881),
.Y(n_6315)
);

NOR2xp33_ASAP7_75t_R g6316 ( 
.A(n_6103),
.B(n_102),
.Y(n_6316)
);

AND2x4_ASAP7_75t_L g6317 ( 
.A(n_6082),
.B(n_5881),
.Y(n_6317)
);

NOR2xp33_ASAP7_75t_R g6318 ( 
.A(n_6259),
.B(n_103),
.Y(n_6318)
);

HB1xp67_ASAP7_75t_L g6319 ( 
.A(n_6036),
.Y(n_6319)
);

NOR2xp33_ASAP7_75t_R g6320 ( 
.A(n_6215),
.B(n_104),
.Y(n_6320)
);

AND2x4_ASAP7_75t_L g6321 ( 
.A(n_6082),
.B(n_5917),
.Y(n_6321)
);

NAND2xp33_ASAP7_75t_R g6322 ( 
.A(n_6220),
.B(n_104),
.Y(n_6322)
);

INVxp67_ASAP7_75t_L g6323 ( 
.A(n_6096),
.Y(n_6323)
);

NAND2xp5_ASAP7_75t_L g6324 ( 
.A(n_6236),
.B(n_6017),
.Y(n_6324)
);

NAND2xp33_ASAP7_75t_R g6325 ( 
.A(n_6220),
.B(n_105),
.Y(n_6325)
);

CKINVDCx5p33_ASAP7_75t_R g6326 ( 
.A(n_6258),
.Y(n_6326)
);

NOR2xp33_ASAP7_75t_R g6327 ( 
.A(n_6209),
.B(n_105),
.Y(n_6327)
);

NAND2xp5_ASAP7_75t_L g6328 ( 
.A(n_6236),
.B(n_6017),
.Y(n_6328)
);

NOR2xp33_ASAP7_75t_R g6329 ( 
.A(n_6213),
.B(n_105),
.Y(n_6329)
);

AND2x4_ASAP7_75t_L g6330 ( 
.A(n_6122),
.B(n_5917),
.Y(n_6330)
);

AND2x2_ASAP7_75t_L g6331 ( 
.A(n_6054),
.B(n_5917),
.Y(n_6331)
);

BUFx10_ASAP7_75t_L g6332 ( 
.A(n_6232),
.Y(n_6332)
);

AND2x2_ASAP7_75t_L g6333 ( 
.A(n_6054),
.B(n_6211),
.Y(n_6333)
);

NOR2xp33_ASAP7_75t_R g6334 ( 
.A(n_6102),
.B(n_6272),
.Y(n_6334)
);

INVxp67_ASAP7_75t_L g6335 ( 
.A(n_6247),
.Y(n_6335)
);

BUFx10_ASAP7_75t_L g6336 ( 
.A(n_6232),
.Y(n_6336)
);

AND2x2_ASAP7_75t_L g6337 ( 
.A(n_6076),
.B(n_5999),
.Y(n_6337)
);

NAND2xp33_ASAP7_75t_R g6338 ( 
.A(n_6263),
.B(n_106),
.Y(n_6338)
);

AND2x4_ASAP7_75t_L g6339 ( 
.A(n_6122),
.B(n_6017),
.Y(n_6339)
);

NAND2xp33_ASAP7_75t_SL g6340 ( 
.A(n_6241),
.B(n_5838),
.Y(n_6340)
);

BUFx3_ASAP7_75t_L g6341 ( 
.A(n_6244),
.Y(n_6341)
);

BUFx3_ASAP7_75t_L g6342 ( 
.A(n_6149),
.Y(n_6342)
);

NAND2xp33_ASAP7_75t_R g6343 ( 
.A(n_6073),
.B(n_106),
.Y(n_6343)
);

NOR2xp33_ASAP7_75t_R g6344 ( 
.A(n_6102),
.B(n_6071),
.Y(n_6344)
);

INVx2_ASAP7_75t_L g6345 ( 
.A(n_6087),
.Y(n_6345)
);

OR2x6_ASAP7_75t_L g6346 ( 
.A(n_6071),
.B(n_5940),
.Y(n_6346)
);

HB1xp67_ASAP7_75t_L g6347 ( 
.A(n_6140),
.Y(n_6347)
);

NAND2xp33_ASAP7_75t_R g6348 ( 
.A(n_6073),
.B(n_107),
.Y(n_6348)
);

NOR2xp33_ASAP7_75t_R g6349 ( 
.A(n_6102),
.B(n_107),
.Y(n_6349)
);

NAND2xp5_ASAP7_75t_L g6350 ( 
.A(n_6221),
.B(n_6017),
.Y(n_6350)
);

NAND2xp33_ASAP7_75t_SL g6351 ( 
.A(n_6197),
.B(n_5912),
.Y(n_6351)
);

BUFx3_ASAP7_75t_L g6352 ( 
.A(n_6149),
.Y(n_6352)
);

AND2x4_ASAP7_75t_L g6353 ( 
.A(n_6129),
.B(n_6014),
.Y(n_6353)
);

NOR2xp33_ASAP7_75t_R g6354 ( 
.A(n_6071),
.B(n_108),
.Y(n_6354)
);

NOR2xp33_ASAP7_75t_R g6355 ( 
.A(n_6208),
.B(n_109),
.Y(n_6355)
);

CKINVDCx5p33_ASAP7_75t_R g6356 ( 
.A(n_6044),
.Y(n_6356)
);

INVxp67_ASAP7_75t_L g6357 ( 
.A(n_6031),
.Y(n_6357)
);

CKINVDCx20_ASAP7_75t_R g6358 ( 
.A(n_6044),
.Y(n_6358)
);

NOR2xp33_ASAP7_75t_L g6359 ( 
.A(n_6032),
.B(n_167),
.Y(n_6359)
);

INVx3_ASAP7_75t_L g6360 ( 
.A(n_6129),
.Y(n_6360)
);

NOR2xp33_ASAP7_75t_R g6361 ( 
.A(n_6196),
.B(n_109),
.Y(n_6361)
);

XNOR2xp5_ASAP7_75t_L g6362 ( 
.A(n_6144),
.B(n_6042),
.Y(n_6362)
);

BUFx10_ASAP7_75t_L g6363 ( 
.A(n_6067),
.Y(n_6363)
);

AND2x4_ASAP7_75t_L g6364 ( 
.A(n_6067),
.B(n_6001),
.Y(n_6364)
);

AND2x4_ASAP7_75t_L g6365 ( 
.A(n_6118),
.B(n_6007),
.Y(n_6365)
);

NAND2xp33_ASAP7_75t_SL g6366 ( 
.A(n_6229),
.B(n_5943),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_6108),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_6040),
.Y(n_6368)
);

NAND2xp5_ASAP7_75t_L g6369 ( 
.A(n_6170),
.B(n_5961),
.Y(n_6369)
);

NAND2xp33_ASAP7_75t_R g6370 ( 
.A(n_6073),
.B(n_110),
.Y(n_6370)
);

AND2x4_ASAP7_75t_L g6371 ( 
.A(n_6182),
.B(n_6007),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_6110),
.B(n_5994),
.Y(n_6372)
);

BUFx10_ASAP7_75t_L g6373 ( 
.A(n_6219),
.Y(n_6373)
);

XNOR2xp5_ASAP7_75t_L g6374 ( 
.A(n_6144),
.B(n_6053),
.Y(n_6374)
);

NAND2xp33_ASAP7_75t_SL g6375 ( 
.A(n_6231),
.B(n_5953),
.Y(n_6375)
);

NOR2xp33_ASAP7_75t_L g6376 ( 
.A(n_6163),
.B(n_168),
.Y(n_6376)
);

NAND2xp5_ASAP7_75t_L g6377 ( 
.A(n_6114),
.B(n_5998),
.Y(n_6377)
);

NOR2xp33_ASAP7_75t_L g6378 ( 
.A(n_6201),
.B(n_168),
.Y(n_6378)
);

NOR2xp33_ASAP7_75t_R g6379 ( 
.A(n_6216),
.B(n_110),
.Y(n_6379)
);

NAND2xp5_ASAP7_75t_L g6380 ( 
.A(n_6121),
.B(n_5835),
.Y(n_6380)
);

CKINVDCx20_ASAP7_75t_R g6381 ( 
.A(n_6142),
.Y(n_6381)
);

CKINVDCx5p33_ASAP7_75t_R g6382 ( 
.A(n_6224),
.Y(n_6382)
);

NOR2xp33_ASAP7_75t_R g6383 ( 
.A(n_6223),
.B(n_110),
.Y(n_6383)
);

NAND2xp5_ASAP7_75t_L g6384 ( 
.A(n_6141),
.B(n_5835),
.Y(n_6384)
);

AND2x4_ASAP7_75t_L g6385 ( 
.A(n_6178),
.B(n_5885),
.Y(n_6385)
);

NAND2xp33_ASAP7_75t_R g6386 ( 
.A(n_6239),
.B(n_111),
.Y(n_6386)
);

NAND2xp5_ASAP7_75t_L g6387 ( 
.A(n_6145),
.B(n_5885),
.Y(n_6387)
);

NOR2xp33_ASAP7_75t_R g6388 ( 
.A(n_6230),
.B(n_111),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_6158),
.Y(n_6389)
);

NAND2xp5_ASAP7_75t_L g6390 ( 
.A(n_6164),
.B(n_6167),
.Y(n_6390)
);

NOR2xp33_ASAP7_75t_R g6391 ( 
.A(n_6273),
.B(n_6055),
.Y(n_6391)
);

AND2x2_ASAP7_75t_L g6392 ( 
.A(n_6168),
.B(n_5885),
.Y(n_6392)
);

HB1xp67_ASAP7_75t_L g6393 ( 
.A(n_6185),
.Y(n_6393)
);

INVxp67_ASAP7_75t_L g6394 ( 
.A(n_6028),
.Y(n_6394)
);

NAND2xp33_ASAP7_75t_R g6395 ( 
.A(n_6269),
.B(n_111),
.Y(n_6395)
);

NOR2xp33_ASAP7_75t_R g6396 ( 
.A(n_6033),
.B(n_112),
.Y(n_6396)
);

NAND2xp5_ASAP7_75t_L g6397 ( 
.A(n_6046),
.B(n_171),
.Y(n_6397)
);

AND2x2_ASAP7_75t_L g6398 ( 
.A(n_6077),
.B(n_112),
.Y(n_6398)
);

AND2x2_ASAP7_75t_L g6399 ( 
.A(n_6126),
.B(n_112),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_6123),
.Y(n_6400)
);

NOR2xp33_ASAP7_75t_R g6401 ( 
.A(n_6058),
.B(n_113),
.Y(n_6401)
);

INVxp67_ASAP7_75t_L g6402 ( 
.A(n_6093),
.Y(n_6402)
);

NAND2xp33_ASAP7_75t_R g6403 ( 
.A(n_6146),
.B(n_113),
.Y(n_6403)
);

NOR2xp33_ASAP7_75t_R g6404 ( 
.A(n_6233),
.B(n_113),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_6251),
.Y(n_6405)
);

AND2x4_ASAP7_75t_L g6406 ( 
.A(n_6142),
.B(n_114),
.Y(n_6406)
);

HB1xp67_ASAP7_75t_L g6407 ( 
.A(n_6085),
.Y(n_6407)
);

NAND2xp33_ASAP7_75t_R g6408 ( 
.A(n_6169),
.B(n_115),
.Y(n_6408)
);

NOR2xp33_ASAP7_75t_R g6409 ( 
.A(n_6233),
.B(n_115),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_6035),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_6030),
.Y(n_6411)
);

XNOR2xp5_ASAP7_75t_L g6412 ( 
.A(n_6026),
.B(n_116),
.Y(n_6412)
);

INVx1_ASAP7_75t_L g6413 ( 
.A(n_6057),
.Y(n_6413)
);

NAND2xp5_ASAP7_75t_SL g6414 ( 
.A(n_6116),
.B(n_1318),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_6056),
.Y(n_6415)
);

XNOR2xp5_ASAP7_75t_L g6416 ( 
.A(n_6064),
.B(n_116),
.Y(n_6416)
);

BUFx3_ASAP7_75t_L g6417 ( 
.A(n_6112),
.Y(n_6417)
);

NOR2xp33_ASAP7_75t_R g6418 ( 
.A(n_6257),
.B(n_118),
.Y(n_6418)
);

NAND2xp5_ASAP7_75t_L g6419 ( 
.A(n_6092),
.B(n_172),
.Y(n_6419)
);

AND2x4_ASAP7_75t_L g6420 ( 
.A(n_6169),
.B(n_6180),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_L g6421 ( 
.A(n_6083),
.B(n_172),
.Y(n_6421)
);

XNOR2xp5_ASAP7_75t_L g6422 ( 
.A(n_6064),
.B(n_118),
.Y(n_6422)
);

AND2x4_ASAP7_75t_L g6423 ( 
.A(n_6169),
.B(n_6180),
.Y(n_6423)
);

NAND2xp33_ASAP7_75t_SL g6424 ( 
.A(n_6225),
.B(n_119),
.Y(n_6424)
);

AND2x2_ASAP7_75t_L g6425 ( 
.A(n_6187),
.B(n_119),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6143),
.Y(n_6426)
);

CKINVDCx11_ASAP7_75t_R g6427 ( 
.A(n_6191),
.Y(n_6427)
);

NAND2xp5_ASAP7_75t_SL g6428 ( 
.A(n_6105),
.B(n_1320),
.Y(n_6428)
);

NAND2xp33_ASAP7_75t_R g6429 ( 
.A(n_6248),
.B(n_119),
.Y(n_6429)
);

NAND2xp33_ASAP7_75t_R g6430 ( 
.A(n_6248),
.B(n_120),
.Y(n_6430)
);

AND2x4_ASAP7_75t_L g6431 ( 
.A(n_6262),
.B(n_120),
.Y(n_6431)
);

INVxp67_ASAP7_75t_L g6432 ( 
.A(n_6222),
.Y(n_6432)
);

XOR2xp5_ASAP7_75t_L g6433 ( 
.A(n_6074),
.B(n_120),
.Y(n_6433)
);

INVxp67_ASAP7_75t_L g6434 ( 
.A(n_6119),
.Y(n_6434)
);

NAND2xp33_ASAP7_75t_R g6435 ( 
.A(n_6202),
.B(n_121),
.Y(n_6435)
);

AND2x2_ASAP7_75t_L g6436 ( 
.A(n_6100),
.B(n_121),
.Y(n_6436)
);

INVxp67_ASAP7_75t_L g6437 ( 
.A(n_6099),
.Y(n_6437)
);

NAND2xp33_ASAP7_75t_R g6438 ( 
.A(n_6202),
.B(n_122),
.Y(n_6438)
);

AND2x2_ASAP7_75t_L g6439 ( 
.A(n_6127),
.B(n_122),
.Y(n_6439)
);

NAND2xp5_ASAP7_75t_L g6440 ( 
.A(n_6204),
.B(n_173),
.Y(n_6440)
);

OR2x6_ASAP7_75t_L g6441 ( 
.A(n_6138),
.B(n_123),
.Y(n_6441)
);

BUFx10_ASAP7_75t_L g6442 ( 
.A(n_6214),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_6206),
.Y(n_6443)
);

AND2x4_ASAP7_75t_L g6444 ( 
.A(n_6101),
.B(n_123),
.Y(n_6444)
);

AND2x2_ASAP7_75t_L g6445 ( 
.A(n_6130),
.B(n_125),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6022),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_6228),
.B(n_125),
.Y(n_6447)
);

AND2x4_ASAP7_75t_L g6448 ( 
.A(n_6155),
.B(n_125),
.Y(n_6448)
);

XNOR2xp5_ASAP7_75t_L g6449 ( 
.A(n_6265),
.B(n_126),
.Y(n_6449)
);

INVxp67_ASAP7_75t_L g6450 ( 
.A(n_6069),
.Y(n_6450)
);

NOR2xp33_ASAP7_75t_L g6451 ( 
.A(n_6048),
.B(n_174),
.Y(n_6451)
);

BUFx10_ASAP7_75t_L g6452 ( 
.A(n_6240),
.Y(n_6452)
);

AND2x2_ASAP7_75t_L g6453 ( 
.A(n_6029),
.B(n_126),
.Y(n_6453)
);

NAND2xp33_ASAP7_75t_R g6454 ( 
.A(n_6205),
.B(n_126),
.Y(n_6454)
);

CKINVDCx5p33_ASAP7_75t_R g6455 ( 
.A(n_6270),
.Y(n_6455)
);

AND2x4_ASAP7_75t_L g6456 ( 
.A(n_6155),
.B(n_127),
.Y(n_6456)
);

NOR2xp33_ASAP7_75t_L g6457 ( 
.A(n_6120),
.B(n_174),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6045),
.Y(n_6458)
);

NOR2xp33_ASAP7_75t_R g6459 ( 
.A(n_6234),
.B(n_127),
.Y(n_6459)
);

BUFx3_ASAP7_75t_L g6460 ( 
.A(n_6246),
.Y(n_6460)
);

BUFx10_ASAP7_75t_L g6461 ( 
.A(n_6238),
.Y(n_6461)
);

AND2x4_ASAP7_75t_L g6462 ( 
.A(n_6155),
.B(n_127),
.Y(n_6462)
);

INVxp67_ASAP7_75t_L g6463 ( 
.A(n_6139),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6243),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_6070),
.Y(n_6465)
);

AND2x4_ASAP7_75t_L g6466 ( 
.A(n_6050),
.B(n_128),
.Y(n_6466)
);

NAND2xp5_ASAP7_75t_L g6467 ( 
.A(n_6068),
.B(n_175),
.Y(n_6467)
);

NOR2xp33_ASAP7_75t_R g6468 ( 
.A(n_6132),
.B(n_128),
.Y(n_6468)
);

NAND2xp5_ASAP7_75t_L g6469 ( 
.A(n_6177),
.B(n_177),
.Y(n_6469)
);

NAND2xp33_ASAP7_75t_R g6470 ( 
.A(n_6205),
.B(n_128),
.Y(n_6470)
);

AND2x2_ASAP7_75t_L g6471 ( 
.A(n_6199),
.B(n_129),
.Y(n_6471)
);

BUFx3_ASAP7_75t_L g6472 ( 
.A(n_6075),
.Y(n_6472)
);

AND2x4_ASAP7_75t_L g6473 ( 
.A(n_6152),
.B(n_130),
.Y(n_6473)
);

INVxp67_ASAP7_75t_L g6474 ( 
.A(n_6084),
.Y(n_6474)
);

INVxp67_ASAP7_75t_L g6475 ( 
.A(n_6252),
.Y(n_6475)
);

AND2x4_ASAP7_75t_L g6476 ( 
.A(n_6181),
.B(n_131),
.Y(n_6476)
);

NOR2xp33_ASAP7_75t_SL g6477 ( 
.A(n_6059),
.B(n_131),
.Y(n_6477)
);

NOR2xp33_ASAP7_75t_R g6478 ( 
.A(n_6037),
.B(n_132),
.Y(n_6478)
);

NAND2xp33_ASAP7_75t_R g6479 ( 
.A(n_6217),
.B(n_132),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6040),
.Y(n_6480)
);

AND2x4_ASAP7_75t_L g6481 ( 
.A(n_6165),
.B(n_133),
.Y(n_6481)
);

INVxp67_ASAP7_75t_L g6482 ( 
.A(n_6153),
.Y(n_6482)
);

AND2x4_ASAP7_75t_L g6483 ( 
.A(n_6080),
.B(n_133),
.Y(n_6483)
);

BUFx3_ASAP7_75t_L g6484 ( 
.A(n_6075),
.Y(n_6484)
);

NAND2xp5_ASAP7_75t_L g6485 ( 
.A(n_6207),
.B(n_179),
.Y(n_6485)
);

XNOR2xp5_ASAP7_75t_L g6486 ( 
.A(n_6136),
.B(n_133),
.Y(n_6486)
);

AND2x4_ASAP7_75t_L g6487 ( 
.A(n_6111),
.B(n_134),
.Y(n_6487)
);

BUFx3_ASAP7_75t_L g6488 ( 
.A(n_6075),
.Y(n_6488)
);

AND2x2_ASAP7_75t_L g6489 ( 
.A(n_6154),
.B(n_134),
.Y(n_6489)
);

INVxp67_ASAP7_75t_L g6490 ( 
.A(n_6212),
.Y(n_6490)
);

AND2x2_ASAP7_75t_L g6491 ( 
.A(n_6078),
.B(n_134),
.Y(n_6491)
);

XNOR2xp5_ASAP7_75t_L g6492 ( 
.A(n_6095),
.B(n_135),
.Y(n_6492)
);

AND2x4_ASAP7_75t_L g6493 ( 
.A(n_6148),
.B(n_135),
.Y(n_6493)
);

XNOR2xp5_ASAP7_75t_L g6494 ( 
.A(n_6095),
.B(n_6238),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_6065),
.Y(n_6495)
);

AND2x4_ASAP7_75t_L g6496 ( 
.A(n_6150),
.B(n_135),
.Y(n_6496)
);

AND2x4_ASAP7_75t_L g6497 ( 
.A(n_6134),
.B(n_136),
.Y(n_6497)
);

AND2x4_ASAP7_75t_L g6498 ( 
.A(n_6135),
.B(n_136),
.Y(n_6498)
);

NAND2xp5_ASAP7_75t_L g6499 ( 
.A(n_6242),
.B(n_179),
.Y(n_6499)
);

AND2x4_ASAP7_75t_L g6500 ( 
.A(n_6171),
.B(n_6159),
.Y(n_6500)
);

AND2x2_ASAP7_75t_L g6501 ( 
.A(n_6078),
.B(n_137),
.Y(n_6501)
);

NAND2xp5_ASAP7_75t_L g6502 ( 
.A(n_6267),
.B(n_180),
.Y(n_6502)
);

NAND2xp33_ASAP7_75t_R g6503 ( 
.A(n_6217),
.B(n_137),
.Y(n_6503)
);

NAND2xp33_ASAP7_75t_SL g6504 ( 
.A(n_6124),
.B(n_138),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_6065),
.Y(n_6505)
);

INVxp67_ASAP7_75t_L g6506 ( 
.A(n_6226),
.Y(n_6506)
);

CKINVDCx20_ASAP7_75t_R g6507 ( 
.A(n_6091),
.Y(n_6507)
);

AND2x4_ASAP7_75t_L g6508 ( 
.A(n_6184),
.B(n_138),
.Y(n_6508)
);

OR2x4_ASAP7_75t_L g6509 ( 
.A(n_6104),
.B(n_138),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_6081),
.Y(n_6510)
);

NAND2xp33_ASAP7_75t_R g6511 ( 
.A(n_6131),
.B(n_139),
.Y(n_6511)
);

INVx2_ASAP7_75t_L g6512 ( 
.A(n_6131),
.Y(n_6512)
);

INVxp67_ASAP7_75t_L g6513 ( 
.A(n_6166),
.Y(n_6513)
);

AND2x4_ASAP7_75t_L g6514 ( 
.A(n_6066),
.B(n_139),
.Y(n_6514)
);

NAND2xp5_ASAP7_75t_L g6515 ( 
.A(n_6271),
.B(n_181),
.Y(n_6515)
);

AND2x4_ASAP7_75t_L g6516 ( 
.A(n_6113),
.B(n_139),
.Y(n_6516)
);

AND2x2_ASAP7_75t_L g6517 ( 
.A(n_6253),
.B(n_140),
.Y(n_6517)
);

NAND2xp5_ASAP7_75t_L g6518 ( 
.A(n_6193),
.B(n_182),
.Y(n_6518)
);

OAI22xp5_ASAP7_75t_L g6519 ( 
.A1(n_6509),
.A2(n_6147),
.B1(n_6249),
.B2(n_6268),
.Y(n_6519)
);

INVx2_ASAP7_75t_L g6520 ( 
.A(n_6461),
.Y(n_6520)
);

INVx3_ASAP7_75t_L g6521 ( 
.A(n_6294),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_6390),
.Y(n_6522)
);

OR2x2_ASAP7_75t_L g6523 ( 
.A(n_6319),
.B(n_6137),
.Y(n_6523)
);

AND2x2_ASAP7_75t_L g6524 ( 
.A(n_6277),
.B(n_6060),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6393),
.Y(n_6525)
);

AND2x2_ASAP7_75t_L g6526 ( 
.A(n_6281),
.B(n_6333),
.Y(n_6526)
);

BUFx2_ASAP7_75t_L g6527 ( 
.A(n_6274),
.Y(n_6527)
);

INVx2_ASAP7_75t_L g6528 ( 
.A(n_6472),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6341),
.B(n_6098),
.Y(n_6529)
);

AOI21xp33_ASAP7_75t_L g6530 ( 
.A1(n_6309),
.A2(n_6151),
.B(n_6268),
.Y(n_6530)
);

AND2x2_ASAP7_75t_L g6531 ( 
.A(n_6278),
.B(n_6192),
.Y(n_6531)
);

INVx2_ASAP7_75t_L g6532 ( 
.A(n_6484),
.Y(n_6532)
);

AOI211xp5_ASAP7_75t_SL g6533 ( 
.A1(n_6311),
.A2(n_6125),
.B(n_6128),
.C(n_6261),
.Y(n_6533)
);

AND2x4_ASAP7_75t_L g6534 ( 
.A(n_6448),
.B(n_6189),
.Y(n_6534)
);

INVx2_ASAP7_75t_SL g6535 ( 
.A(n_6332),
.Y(n_6535)
);

HB1xp67_ASAP7_75t_L g6536 ( 
.A(n_6397),
.Y(n_6536)
);

AND2x2_ASAP7_75t_L g6537 ( 
.A(n_6278),
.B(n_6254),
.Y(n_6537)
);

BUFx8_ASAP7_75t_L g6538 ( 
.A(n_6292),
.Y(n_6538)
);

INVx2_ASAP7_75t_L g6539 ( 
.A(n_6488),
.Y(n_6539)
);

AND2x4_ASAP7_75t_L g6540 ( 
.A(n_6448),
.B(n_6160),
.Y(n_6540)
);

AND2x2_ASAP7_75t_L g6541 ( 
.A(n_6280),
.B(n_6157),
.Y(n_6541)
);

OR2x6_ASAP7_75t_L g6542 ( 
.A(n_6456),
.B(n_6179),
.Y(n_6542)
);

AND2x4_ASAP7_75t_L g6543 ( 
.A(n_6456),
.B(n_6256),
.Y(n_6543)
);

INVx2_ASAP7_75t_L g6544 ( 
.A(n_6368),
.Y(n_6544)
);

AND2x2_ASAP7_75t_L g6545 ( 
.A(n_6280),
.B(n_6425),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6491),
.B(n_6264),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_6480),
.Y(n_6547)
);

INVx2_ASAP7_75t_SL g6548 ( 
.A(n_6336),
.Y(n_6548)
);

INVx2_ASAP7_75t_L g6549 ( 
.A(n_6501),
.Y(n_6549)
);

AND2x2_ASAP7_75t_L g6550 ( 
.A(n_6344),
.B(n_6227),
.Y(n_6550)
);

INVx2_ASAP7_75t_L g6551 ( 
.A(n_6512),
.Y(n_6551)
);

INVx2_ASAP7_75t_L g6552 ( 
.A(n_6356),
.Y(n_6552)
);

INVx2_ASAP7_75t_L g6553 ( 
.A(n_6431),
.Y(n_6553)
);

HB1xp67_ASAP7_75t_L g6554 ( 
.A(n_6284),
.Y(n_6554)
);

INVx2_ASAP7_75t_L g6555 ( 
.A(n_6431),
.Y(n_6555)
);

AND2x4_ASAP7_75t_L g6556 ( 
.A(n_6462),
.B(n_6162),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6285),
.Y(n_6557)
);

HB1xp67_ASAP7_75t_L g6558 ( 
.A(n_6490),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_6481),
.Y(n_6559)
);

INVx2_ASAP7_75t_L g6560 ( 
.A(n_6481),
.Y(n_6560)
);

AND2x2_ASAP7_75t_L g6561 ( 
.A(n_6300),
.B(n_6106),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_6297),
.Y(n_6562)
);

OR2x2_ASAP7_75t_L g6563 ( 
.A(n_6413),
.B(n_6176),
.Y(n_6563)
);

INVx1_ASAP7_75t_L g6564 ( 
.A(n_6305),
.Y(n_6564)
);

AND2x2_ASAP7_75t_L g6565 ( 
.A(n_6360),
.B(n_6200),
.Y(n_6565)
);

NOR2xp33_ASAP7_75t_L g6566 ( 
.A(n_6287),
.B(n_6266),
.Y(n_6566)
);

INVx1_ASAP7_75t_L g6567 ( 
.A(n_6310),
.Y(n_6567)
);

INVx3_ASAP7_75t_L g6568 ( 
.A(n_6298),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6367),
.Y(n_6569)
);

BUFx2_ASAP7_75t_L g6570 ( 
.A(n_6279),
.Y(n_6570)
);

INVx4_ASAP7_75t_L g6571 ( 
.A(n_6326),
.Y(n_6571)
);

INVx4_ASAP7_75t_L g6572 ( 
.A(n_6342),
.Y(n_6572)
);

INVx2_ASAP7_75t_L g6573 ( 
.A(n_6494),
.Y(n_6573)
);

INVx1_ASAP7_75t_L g6574 ( 
.A(n_6389),
.Y(n_6574)
);

AND2x4_ASAP7_75t_L g6575 ( 
.A(n_6462),
.B(n_6109),
.Y(n_6575)
);

INVxp67_ASAP7_75t_L g6576 ( 
.A(n_6322),
.Y(n_6576)
);

AND2x2_ASAP7_75t_L g6577 ( 
.A(n_6299),
.B(n_6183),
.Y(n_6577)
);

AND2x4_ASAP7_75t_L g6578 ( 
.A(n_6508),
.B(n_6109),
.Y(n_6578)
);

AND2x2_ASAP7_75t_L g6579 ( 
.A(n_6299),
.B(n_6183),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_6347),
.Y(n_6580)
);

INVx2_ASAP7_75t_L g6581 ( 
.A(n_6497),
.Y(n_6581)
);

NAND2xp5_ASAP7_75t_L g6582 ( 
.A(n_6506),
.B(n_6091),
.Y(n_6582)
);

BUFx6f_ASAP7_75t_L g6583 ( 
.A(n_6518),
.Y(n_6583)
);

BUFx3_ASAP7_75t_L g6584 ( 
.A(n_6293),
.Y(n_6584)
);

INVx2_ASAP7_75t_SL g6585 ( 
.A(n_6508),
.Y(n_6585)
);

AND2x2_ASAP7_75t_L g6586 ( 
.A(n_6466),
.B(n_6174),
.Y(n_6586)
);

HB1xp67_ASAP7_75t_L g6587 ( 
.A(n_6286),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6405),
.Y(n_6588)
);

AND2x2_ASAP7_75t_L g6589 ( 
.A(n_6466),
.B(n_6195),
.Y(n_6589)
);

NOR2xp33_ASAP7_75t_L g6590 ( 
.A(n_6352),
.B(n_6359),
.Y(n_6590)
);

AND2x2_ASAP7_75t_L g6591 ( 
.A(n_6407),
.B(n_6094),
.Y(n_6591)
);

INVx1_ASAP7_75t_L g6592 ( 
.A(n_6443),
.Y(n_6592)
);

INVx3_ASAP7_75t_L g6593 ( 
.A(n_6313),
.Y(n_6593)
);

INVx2_ASAP7_75t_L g6594 ( 
.A(n_6497),
.Y(n_6594)
);

NAND2x1p5_ASAP7_75t_L g6595 ( 
.A(n_6339),
.B(n_6188),
.Y(n_6595)
);

INVx2_ASAP7_75t_SL g6596 ( 
.A(n_6363),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6464),
.Y(n_6597)
);

AND2x2_ASAP7_75t_L g6598 ( 
.A(n_6334),
.B(n_6255),
.Y(n_6598)
);

NAND2xp5_ASAP7_75t_L g6599 ( 
.A(n_6421),
.B(n_6049),
.Y(n_6599)
);

HB1xp67_ASAP7_75t_L g6600 ( 
.A(n_6380),
.Y(n_6600)
);

AND2x2_ASAP7_75t_L g6601 ( 
.A(n_6291),
.B(n_6331),
.Y(n_6601)
);

INVx2_ASAP7_75t_L g6602 ( 
.A(n_6498),
.Y(n_6602)
);

HB1xp67_ASAP7_75t_L g6603 ( 
.A(n_6384),
.Y(n_6603)
);

INVx1_ASAP7_75t_L g6604 ( 
.A(n_6400),
.Y(n_6604)
);

NAND2xp5_ASAP7_75t_L g6605 ( 
.A(n_6335),
.B(n_6237),
.Y(n_6605)
);

AND2x2_ASAP7_75t_L g6606 ( 
.A(n_6291),
.B(n_6115),
.Y(n_6606)
);

BUFx2_ASAP7_75t_L g6607 ( 
.A(n_6327),
.Y(n_6607)
);

INVx1_ASAP7_75t_SL g6608 ( 
.A(n_6312),
.Y(n_6608)
);

INVx4_ASAP7_75t_L g6609 ( 
.A(n_6489),
.Y(n_6609)
);

INVx2_ASAP7_75t_L g6610 ( 
.A(n_6498),
.Y(n_6610)
);

BUFx2_ASAP7_75t_L g6611 ( 
.A(n_6404),
.Y(n_6611)
);

AND2x2_ASAP7_75t_L g6612 ( 
.A(n_6323),
.B(n_6173),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_6510),
.Y(n_6613)
);

AND2x4_ASAP7_75t_L g6614 ( 
.A(n_6339),
.B(n_6260),
.Y(n_6614)
);

HB1xp67_ASAP7_75t_L g6615 ( 
.A(n_6387),
.Y(n_6615)
);

BUFx2_ASAP7_75t_L g6616 ( 
.A(n_6409),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_6419),
.Y(n_6617)
);

AND2x4_ASAP7_75t_L g6618 ( 
.A(n_6330),
.B(n_6107),
.Y(n_6618)
);

AND2x2_ASAP7_75t_L g6619 ( 
.A(n_6295),
.B(n_6188),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6337),
.Y(n_6620)
);

AND2x4_ASAP7_75t_L g6621 ( 
.A(n_6330),
.B(n_6198),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_6295),
.B(n_6210),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_6514),
.Y(n_6623)
);

AND2x2_ASAP7_75t_L g6624 ( 
.A(n_6307),
.B(n_140),
.Y(n_6624)
);

AND2x2_ASAP7_75t_L g6625 ( 
.A(n_6315),
.B(n_140),
.Y(n_6625)
);

AO21x2_ASAP7_75t_L g6626 ( 
.A1(n_6418),
.A2(n_6172),
.B(n_6156),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6514),
.Y(n_6627)
);

BUFx2_ASAP7_75t_L g6628 ( 
.A(n_6382),
.Y(n_6628)
);

AND2x2_ASAP7_75t_L g6629 ( 
.A(n_6317),
.B(n_141),
.Y(n_6629)
);

AND2x2_ASAP7_75t_SL g6630 ( 
.A(n_6444),
.B(n_6245),
.Y(n_6630)
);

INVx3_ASAP7_75t_L g6631 ( 
.A(n_6321),
.Y(n_6631)
);

AND2x2_ASAP7_75t_L g6632 ( 
.A(n_6317),
.B(n_141),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6516),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_6516),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6372),
.Y(n_6635)
);

INVx2_ASAP7_75t_L g6636 ( 
.A(n_6290),
.Y(n_6636)
);

NOR2x1_ASAP7_75t_L g6637 ( 
.A(n_6398),
.B(n_141),
.Y(n_6637)
);

AND2x2_ASAP7_75t_L g6638 ( 
.A(n_6304),
.B(n_142),
.Y(n_6638)
);

AND2x4_ASAP7_75t_L g6639 ( 
.A(n_6483),
.B(n_142),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6377),
.Y(n_6640)
);

AND2x2_ASAP7_75t_L g6641 ( 
.A(n_6483),
.B(n_6417),
.Y(n_6641)
);

HB1xp67_ASAP7_75t_L g6642 ( 
.A(n_6426),
.Y(n_6642)
);

AND2x2_ASAP7_75t_L g6643 ( 
.A(n_6399),
.B(n_143),
.Y(n_6643)
);

AND2x2_ASAP7_75t_L g6644 ( 
.A(n_6447),
.B(n_143),
.Y(n_6644)
);

OA21x2_ASAP7_75t_L g6645 ( 
.A1(n_6495),
.A2(n_143),
.B(n_144),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6505),
.Y(n_6646)
);

AND2x2_ASAP7_75t_L g6647 ( 
.A(n_6394),
.B(n_144),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_6345),
.Y(n_6648)
);

INVx3_ASAP7_75t_L g6649 ( 
.A(n_6321),
.Y(n_6649)
);

BUFx2_ASAP7_75t_L g6650 ( 
.A(n_6424),
.Y(n_6650)
);

AND2x4_ASAP7_75t_L g6651 ( 
.A(n_6473),
.B(n_145),
.Y(n_6651)
);

AND2x4_ASAP7_75t_L g6652 ( 
.A(n_6473),
.B(n_146),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_6517),
.Y(n_6653)
);

INVx2_ASAP7_75t_L g6654 ( 
.A(n_6442),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_6410),
.Y(n_6655)
);

AND2x2_ASAP7_75t_L g6656 ( 
.A(n_6411),
.B(n_146),
.Y(n_6656)
);

AOI22xp33_ASAP7_75t_L g6657 ( 
.A1(n_6460),
.A2(n_147),
.B1(n_148),
.B2(n_183),
.Y(n_6657)
);

INVx2_ASAP7_75t_L g6658 ( 
.A(n_6373),
.Y(n_6658)
);

HB1xp67_ASAP7_75t_L g6659 ( 
.A(n_6306),
.Y(n_6659)
);

INVx2_ASAP7_75t_SL g6660 ( 
.A(n_6289),
.Y(n_6660)
);

INVx2_ASAP7_75t_L g6661 ( 
.A(n_6358),
.Y(n_6661)
);

AND2x2_ASAP7_75t_L g6662 ( 
.A(n_6445),
.B(n_147),
.Y(n_6662)
);

OAI22xp33_ASAP7_75t_L g6663 ( 
.A1(n_6477),
.A2(n_147),
.B1(n_185),
.B2(n_184),
.Y(n_6663)
);

INVx2_ASAP7_75t_L g6664 ( 
.A(n_6324),
.Y(n_6664)
);

INVx2_ASAP7_75t_SL g6665 ( 
.A(n_6493),
.Y(n_6665)
);

INVx2_ASAP7_75t_L g6666 ( 
.A(n_6328),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_6446),
.Y(n_6667)
);

OAI22xp5_ASAP7_75t_L g6668 ( 
.A1(n_6357),
.A2(n_187),
.B1(n_184),
.B2(n_186),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6487),
.Y(n_6669)
);

OR2x2_ASAP7_75t_L g6670 ( 
.A(n_6308),
.B(n_188),
.Y(n_6670)
);

OAI321xp33_ASAP7_75t_L g6671 ( 
.A1(n_6450),
.A2(n_192),
.A3(n_194),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_6671)
);

OAI22xp5_ASAP7_75t_L g6672 ( 
.A1(n_6301),
.A2(n_195),
.B1(n_190),
.B2(n_193),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6487),
.Y(n_6673)
);

INVx4_ASAP7_75t_L g6674 ( 
.A(n_6436),
.Y(n_6674)
);

NOR4xp25_ASAP7_75t_SL g6675 ( 
.A(n_6275),
.B(n_197),
.C(n_195),
.D(n_196),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6458),
.Y(n_6676)
);

AOI22xp33_ASAP7_75t_L g6677 ( 
.A1(n_6507),
.A2(n_200),
.B1(n_196),
.B2(n_199),
.Y(n_6677)
);

INVx2_ASAP7_75t_L g6678 ( 
.A(n_6467),
.Y(n_6678)
);

INVx4_ASAP7_75t_L g6679 ( 
.A(n_6441),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_6465),
.Y(n_6680)
);

AND2x2_ASAP7_75t_L g6681 ( 
.A(n_6437),
.B(n_199),
.Y(n_6681)
);

AND2x2_ASAP7_75t_L g6682 ( 
.A(n_6306),
.B(n_6439),
.Y(n_6682)
);

AND2x4_ASAP7_75t_L g6683 ( 
.A(n_6476),
.B(n_202),
.Y(n_6683)
);

INVx2_ASAP7_75t_L g6684 ( 
.A(n_6385),
.Y(n_6684)
);

NAND2xp5_ASAP7_75t_L g6685 ( 
.A(n_6432),
.B(n_202),
.Y(n_6685)
);

AND2x2_ASAP7_75t_L g6686 ( 
.A(n_6476),
.B(n_203),
.Y(n_6686)
);

AOI22xp33_ASAP7_75t_L g6687 ( 
.A1(n_6402),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_6687)
);

BUFx6f_ASAP7_75t_L g6688 ( 
.A(n_6414),
.Y(n_6688)
);

NOR2x1p5_ASAP7_75t_L g6689 ( 
.A(n_6369),
.B(n_205),
.Y(n_6689)
);

BUFx6f_ASAP7_75t_L g6690 ( 
.A(n_6469),
.Y(n_6690)
);

INVx4_ASAP7_75t_L g6691 ( 
.A(n_6441),
.Y(n_6691)
);

HB1xp67_ASAP7_75t_L g6692 ( 
.A(n_6415),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_6350),
.Y(n_6693)
);

HB1xp67_ASAP7_75t_L g6694 ( 
.A(n_6474),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6453),
.Y(n_6695)
);

NAND3xp33_ASAP7_75t_L g6696 ( 
.A(n_6463),
.B(n_206),
.C(n_207),
.Y(n_6696)
);

INVx1_ASAP7_75t_L g6697 ( 
.A(n_6471),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_6302),
.Y(n_6698)
);

HB1xp67_ASAP7_75t_L g6699 ( 
.A(n_6482),
.Y(n_6699)
);

INVx2_ASAP7_75t_L g6700 ( 
.A(n_6385),
.Y(n_6700)
);

OR2x2_ASAP7_75t_L g6701 ( 
.A(n_6444),
.B(n_209),
.Y(n_6701)
);

AND2x2_ASAP7_75t_L g6702 ( 
.A(n_6314),
.B(n_210),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6486),
.Y(n_6703)
);

INVx1_ASAP7_75t_L g6704 ( 
.A(n_6492),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6433),
.Y(n_6705)
);

INVx2_ASAP7_75t_SL g6706 ( 
.A(n_6493),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6496),
.Y(n_6707)
);

INVx6_ASAP7_75t_L g6708 ( 
.A(n_6452),
.Y(n_6708)
);

NOR2x1_ASAP7_75t_L g6709 ( 
.A(n_6457),
.B(n_212),
.Y(n_6709)
);

BUFx3_ASAP7_75t_L g6710 ( 
.A(n_6427),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6303),
.B(n_212),
.Y(n_6711)
);

INVx2_ASAP7_75t_L g6712 ( 
.A(n_6371),
.Y(n_6712)
);

AND2x4_ASAP7_75t_L g6713 ( 
.A(n_6420),
.B(n_213),
.Y(n_6713)
);

BUFx2_ASAP7_75t_L g6714 ( 
.A(n_6318),
.Y(n_6714)
);

AND2x4_ASAP7_75t_L g6715 ( 
.A(n_6420),
.B(n_215),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6496),
.Y(n_6716)
);

INVx1_ASAP7_75t_L g6717 ( 
.A(n_6375),
.Y(n_6717)
);

AND2x4_ASAP7_75t_SL g6718 ( 
.A(n_6346),
.B(n_6423),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_6406),
.Y(n_6719)
);

AND2x2_ASAP7_75t_L g6720 ( 
.A(n_6346),
.B(n_215),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6406),
.Y(n_6721)
);

INVx2_ASAP7_75t_L g6722 ( 
.A(n_6371),
.Y(n_6722)
);

OAI22xp33_ASAP7_75t_L g6723 ( 
.A1(n_6408),
.A2(n_220),
.B1(n_217),
.B2(n_218),
.Y(n_6723)
);

OA21x2_ASAP7_75t_L g6724 ( 
.A1(n_6434),
.A2(n_1325),
.B(n_1323),
.Y(n_6724)
);

INVx1_ASAP7_75t_L g6725 ( 
.A(n_6366),
.Y(n_6725)
);

HB1xp67_ASAP7_75t_L g6726 ( 
.A(n_6499),
.Y(n_6726)
);

AND2x2_ASAP7_75t_L g6727 ( 
.A(n_6423),
.B(n_217),
.Y(n_6727)
);

AND2x2_ASAP7_75t_L g6728 ( 
.A(n_6378),
.B(n_218),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6502),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_6364),
.Y(n_6730)
);

AND2x2_ASAP7_75t_L g6731 ( 
.A(n_6282),
.B(n_220),
.Y(n_6731)
);

AOI22xp5_ASAP7_75t_L g6732 ( 
.A1(n_6395),
.A2(n_1325),
.B1(n_1326),
.B2(n_1323),
.Y(n_6732)
);

AND2x2_ASAP7_75t_L g6733 ( 
.A(n_6282),
.B(n_221),
.Y(n_6733)
);

AND2x2_ASAP7_75t_L g6734 ( 
.A(n_6500),
.B(n_221),
.Y(n_6734)
);

NAND2xp5_ASAP7_75t_L g6735 ( 
.A(n_6276),
.B(n_6288),
.Y(n_6735)
);

INVx3_ASAP7_75t_L g6736 ( 
.A(n_6353),
.Y(n_6736)
);

INVx2_ASAP7_75t_L g6737 ( 
.A(n_6364),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6515),
.Y(n_6738)
);

INVx2_ASAP7_75t_L g6739 ( 
.A(n_6416),
.Y(n_6739)
);

INVx3_ASAP7_75t_L g6740 ( 
.A(n_6353),
.Y(n_6740)
);

OR2x2_ASAP7_75t_L g6741 ( 
.A(n_6513),
.B(n_222),
.Y(n_6741)
);

HB1xp67_ASAP7_75t_L g6742 ( 
.A(n_6475),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6500),
.B(n_6392),
.Y(n_6743)
);

HB1xp67_ASAP7_75t_L g6744 ( 
.A(n_6325),
.Y(n_6744)
);

INVx1_ASAP7_75t_L g6745 ( 
.A(n_6351),
.Y(n_6745)
);

AND2x2_ASAP7_75t_L g6746 ( 
.A(n_6316),
.B(n_222),
.Y(n_6746)
);

NAND2xp5_ASAP7_75t_L g6747 ( 
.A(n_6428),
.B(n_223),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6422),
.Y(n_6748)
);

NAND3xp33_ASAP7_75t_L g6749 ( 
.A(n_6558),
.B(n_6451),
.C(n_6511),
.Y(n_6749)
);

NAND2xp5_ASAP7_75t_L g6750 ( 
.A(n_6536),
.B(n_6391),
.Y(n_6750)
);

NOR3xp33_ASAP7_75t_L g6751 ( 
.A(n_6572),
.B(n_6376),
.C(n_6485),
.Y(n_6751)
);

AND2x2_ASAP7_75t_L g6752 ( 
.A(n_6527),
.B(n_6296),
.Y(n_6752)
);

NAND2xp5_ASAP7_75t_L g6753 ( 
.A(n_6536),
.B(n_6383),
.Y(n_6753)
);

NAND2xp5_ASAP7_75t_L g6754 ( 
.A(n_6558),
.B(n_6355),
.Y(n_6754)
);

OA21x2_ASAP7_75t_L g6755 ( 
.A1(n_6582),
.A2(n_6362),
.B(n_6412),
.Y(n_6755)
);

OAI22xp5_ASAP7_75t_L g6756 ( 
.A1(n_6708),
.A2(n_6455),
.B1(n_6381),
.B2(n_6440),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_SL g6757 ( 
.A(n_6660),
.B(n_6340),
.Y(n_6757)
);

AND2x2_ASAP7_75t_L g6758 ( 
.A(n_6545),
.B(n_6628),
.Y(n_6758)
);

AND2x2_ASAP7_75t_L g6759 ( 
.A(n_6570),
.B(n_6388),
.Y(n_6759)
);

NAND2xp5_ASAP7_75t_SL g6760 ( 
.A(n_6660),
.B(n_6365),
.Y(n_6760)
);

AOI22xp5_ASAP7_75t_L g6761 ( 
.A1(n_6519),
.A2(n_6403),
.B1(n_6338),
.B2(n_6348),
.Y(n_6761)
);

AND2x2_ASAP7_75t_L g6762 ( 
.A(n_6526),
.B(n_6283),
.Y(n_6762)
);

AND2x2_ASAP7_75t_L g6763 ( 
.A(n_6572),
.B(n_6329),
.Y(n_6763)
);

NOR3xp33_ASAP7_75t_L g6764 ( 
.A(n_6671),
.B(n_6504),
.C(n_6365),
.Y(n_6764)
);

AND2x2_ASAP7_75t_L g6765 ( 
.A(n_6585),
.B(n_6401),
.Y(n_6765)
);

NAND2xp5_ASAP7_75t_L g6766 ( 
.A(n_6726),
.B(n_6379),
.Y(n_6766)
);

NOR2xp33_ASAP7_75t_SL g6767 ( 
.A(n_6679),
.B(n_6320),
.Y(n_6767)
);

AND2x2_ASAP7_75t_L g6768 ( 
.A(n_6585),
.B(n_6349),
.Y(n_6768)
);

NAND3xp33_ASAP7_75t_L g6769 ( 
.A(n_6690),
.B(n_6590),
.C(n_6533),
.Y(n_6769)
);

OAI21xp5_ASAP7_75t_SL g6770 ( 
.A1(n_6745),
.A2(n_6449),
.B(n_6374),
.Y(n_6770)
);

OAI21xp33_ASAP7_75t_L g6771 ( 
.A1(n_6590),
.A2(n_6396),
.B(n_6478),
.Y(n_6771)
);

NAND3xp33_ASAP7_75t_L g6772 ( 
.A(n_6690),
.B(n_6430),
.C(n_6429),
.Y(n_6772)
);

OAI22xp5_ASAP7_75t_L g6773 ( 
.A1(n_6708),
.A2(n_6370),
.B1(n_6343),
.B2(n_6386),
.Y(n_6773)
);

AOI22xp33_ASAP7_75t_L g6774 ( 
.A1(n_6744),
.A2(n_6468),
.B1(n_6459),
.B2(n_6361),
.Y(n_6774)
);

NAND2xp5_ASAP7_75t_L g6775 ( 
.A(n_6726),
.B(n_6354),
.Y(n_6775)
);

NAND2xp5_ASAP7_75t_SL g6776 ( 
.A(n_6713),
.B(n_6435),
.Y(n_6776)
);

NAND2xp5_ASAP7_75t_L g6777 ( 
.A(n_6742),
.B(n_224),
.Y(n_6777)
);

AND2x2_ASAP7_75t_L g6778 ( 
.A(n_6521),
.B(n_224),
.Y(n_6778)
);

NAND2xp5_ASAP7_75t_SL g6779 ( 
.A(n_6713),
.B(n_6438),
.Y(n_6779)
);

AND2x2_ASAP7_75t_L g6780 ( 
.A(n_6521),
.B(n_226),
.Y(n_6780)
);

NAND2xp5_ASAP7_75t_L g6781 ( 
.A(n_6742),
.B(n_229),
.Y(n_6781)
);

NAND2xp5_ASAP7_75t_L g6782 ( 
.A(n_6647),
.B(n_229),
.Y(n_6782)
);

NAND3xp33_ASAP7_75t_L g6783 ( 
.A(n_6690),
.B(n_6470),
.C(n_6454),
.Y(n_6783)
);

AND2x2_ASAP7_75t_L g6784 ( 
.A(n_6568),
.B(n_230),
.Y(n_6784)
);

NOR2xp33_ASAP7_75t_R g6785 ( 
.A(n_6538),
.B(n_6503),
.Y(n_6785)
);

OAI21xp5_ASAP7_75t_L g6786 ( 
.A1(n_6744),
.A2(n_6479),
.B(n_231),
.Y(n_6786)
);

NAND2xp5_ASAP7_75t_L g6787 ( 
.A(n_6678),
.B(n_6656),
.Y(n_6787)
);

AND2x2_ASAP7_75t_L g6788 ( 
.A(n_6568),
.B(n_231),
.Y(n_6788)
);

AOI22xp5_ASAP7_75t_L g6789 ( 
.A1(n_6599),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_6789)
);

AOI22x1_ASAP7_75t_SL g6790 ( 
.A1(n_6593),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_6790)
);

AOI21xp5_ASAP7_75t_L g6791 ( 
.A1(n_6530),
.A2(n_236),
.B(n_237),
.Y(n_6791)
);

NAND2xp5_ASAP7_75t_L g6792 ( 
.A(n_6678),
.B(n_238),
.Y(n_6792)
);

OAI21xp5_ASAP7_75t_L g6793 ( 
.A1(n_6576),
.A2(n_239),
.B(n_241),
.Y(n_6793)
);

OAI21xp5_ASAP7_75t_L g6794 ( 
.A1(n_6576),
.A2(n_239),
.B(n_241),
.Y(n_6794)
);

AND2x2_ASAP7_75t_L g6795 ( 
.A(n_6593),
.B(n_242),
.Y(n_6795)
);

NAND2xp5_ASAP7_75t_L g6796 ( 
.A(n_6690),
.B(n_242),
.Y(n_6796)
);

NAND2xp5_ASAP7_75t_L g6797 ( 
.A(n_6638),
.B(n_243),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_SL g6798 ( 
.A(n_6713),
.B(n_245),
.Y(n_6798)
);

AOI221xp5_ASAP7_75t_L g6799 ( 
.A1(n_6591),
.A2(n_248),
.B1(n_245),
.B2(n_246),
.C(n_249),
.Y(n_6799)
);

OAI21xp5_ASAP7_75t_L g6800 ( 
.A1(n_6723),
.A2(n_246),
.B(n_248),
.Y(n_6800)
);

AOI22xp33_ASAP7_75t_SL g6801 ( 
.A1(n_6743),
.A2(n_255),
.B1(n_250),
.B2(n_252),
.Y(n_6801)
);

OAI221xp5_ASAP7_75t_SL g6802 ( 
.A1(n_6650),
.A2(n_258),
.B1(n_250),
.B2(n_252),
.C(n_259),
.Y(n_6802)
);

NAND3xp33_ASAP7_75t_L g6803 ( 
.A(n_6583),
.B(n_258),
.C(n_259),
.Y(n_6803)
);

OAI21xp5_ASAP7_75t_SL g6804 ( 
.A1(n_6520),
.A2(n_260),
.B(n_263),
.Y(n_6804)
);

OA21x2_ASAP7_75t_L g6805 ( 
.A1(n_6735),
.A2(n_264),
.B(n_265),
.Y(n_6805)
);

OAI21xp5_ASAP7_75t_SL g6806 ( 
.A1(n_6520),
.A2(n_264),
.B(n_265),
.Y(n_6806)
);

OAI221xp5_ASAP7_75t_SL g6807 ( 
.A1(n_6717),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.C(n_269),
.Y(n_6807)
);

NAND2xp5_ASAP7_75t_L g6808 ( 
.A(n_6583),
.B(n_267),
.Y(n_6808)
);

NAND3xp33_ASAP7_75t_L g6809 ( 
.A(n_6583),
.B(n_269),
.C(n_270),
.Y(n_6809)
);

NAND3xp33_ASAP7_75t_L g6810 ( 
.A(n_6583),
.B(n_270),
.C(n_271),
.Y(n_6810)
);

OAI22xp5_ASAP7_75t_L g6811 ( 
.A1(n_6708),
.A2(n_274),
.B1(n_271),
.B2(n_273),
.Y(n_6811)
);

NAND3xp33_ASAP7_75t_L g6812 ( 
.A(n_6587),
.B(n_274),
.C(n_275),
.Y(n_6812)
);

NAND2xp5_ASAP7_75t_L g6813 ( 
.A(n_6729),
.B(n_275),
.Y(n_6813)
);

HB1xp67_ASAP7_75t_L g6814 ( 
.A(n_6658),
.Y(n_6814)
);

NAND2xp5_ASAP7_75t_L g6815 ( 
.A(n_6738),
.B(n_276),
.Y(n_6815)
);

OAI21xp5_ASAP7_75t_SL g6816 ( 
.A1(n_6586),
.A2(n_277),
.B(n_278),
.Y(n_6816)
);

OAI21xp5_ASAP7_75t_SL g6817 ( 
.A1(n_6654),
.A2(n_280),
.B(n_282),
.Y(n_6817)
);

NAND2xp5_ASAP7_75t_L g6818 ( 
.A(n_6698),
.B(n_6587),
.Y(n_6818)
);

NAND2xp5_ASAP7_75t_L g6819 ( 
.A(n_6694),
.B(n_280),
.Y(n_6819)
);

OAI21xp5_ASAP7_75t_L g6820 ( 
.A1(n_6723),
.A2(n_282),
.B(n_283),
.Y(n_6820)
);

NAND2xp5_ASAP7_75t_L g6821 ( 
.A(n_6694),
.B(n_283),
.Y(n_6821)
);

NAND2xp5_ASAP7_75t_L g6822 ( 
.A(n_6681),
.B(n_284),
.Y(n_6822)
);

NOR2xp33_ASAP7_75t_SL g6823 ( 
.A(n_6679),
.B(n_284),
.Y(n_6823)
);

OAI21xp5_ASAP7_75t_SL g6824 ( 
.A1(n_6654),
.A2(n_285),
.B(n_286),
.Y(n_6824)
);

AOI221xp5_ASAP7_75t_L g6825 ( 
.A1(n_6672),
.A2(n_289),
.B1(n_285),
.B2(n_288),
.C(n_290),
.Y(n_6825)
);

AND2x2_ASAP7_75t_L g6826 ( 
.A(n_6710),
.B(n_288),
.Y(n_6826)
);

NAND2xp5_ASAP7_75t_L g6827 ( 
.A(n_6617),
.B(n_291),
.Y(n_6827)
);

OAI22xp5_ASAP7_75t_L g6828 ( 
.A1(n_6658),
.A2(n_295),
.B1(n_292),
.B2(n_294),
.Y(n_6828)
);

AND2x2_ASAP7_75t_L g6829 ( 
.A(n_6710),
.B(n_294),
.Y(n_6829)
);

NAND2xp5_ASAP7_75t_L g6830 ( 
.A(n_6531),
.B(n_296),
.Y(n_6830)
);

OAI21xp33_ASAP7_75t_SL g6831 ( 
.A1(n_6542),
.A2(n_296),
.B(n_297),
.Y(n_6831)
);

NAND2xp5_ASAP7_75t_L g6832 ( 
.A(n_6674),
.B(n_297),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_L g6833 ( 
.A(n_6674),
.B(n_298),
.Y(n_6833)
);

AOI22xp5_ASAP7_75t_L g6834 ( 
.A1(n_6689),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_6834)
);

AND2x2_ASAP7_75t_L g6835 ( 
.A(n_6535),
.B(n_301),
.Y(n_6835)
);

OA21x2_ASAP7_75t_L g6836 ( 
.A1(n_6605),
.A2(n_302),
.B(n_303),
.Y(n_6836)
);

OAI22xp5_ASAP7_75t_L g6837 ( 
.A1(n_6542),
.A2(n_305),
.B1(n_302),
.B2(n_304),
.Y(n_6837)
);

INVx1_ASAP7_75t_L g6838 ( 
.A(n_6554),
.Y(n_6838)
);

AND2x2_ASAP7_75t_L g6839 ( 
.A(n_6535),
.B(n_306),
.Y(n_6839)
);

AND2x2_ASAP7_75t_L g6840 ( 
.A(n_6548),
.B(n_308),
.Y(n_6840)
);

NAND2xp5_ASAP7_75t_L g6841 ( 
.A(n_6554),
.B(n_309),
.Y(n_6841)
);

NAND2xp5_ASAP7_75t_L g6842 ( 
.A(n_6549),
.B(n_309),
.Y(n_6842)
);

OAI21xp5_ASAP7_75t_SL g6843 ( 
.A1(n_6725),
.A2(n_311),
.B(n_312),
.Y(n_6843)
);

NAND2xp5_ASAP7_75t_L g6844 ( 
.A(n_6549),
.B(n_312),
.Y(n_6844)
);

NAND3xp33_ASAP7_75t_L g6845 ( 
.A(n_6600),
.B(n_313),
.C(n_314),
.Y(n_6845)
);

NAND2xp5_ASAP7_75t_L g6846 ( 
.A(n_6734),
.B(n_313),
.Y(n_6846)
);

AND2x2_ASAP7_75t_L g6847 ( 
.A(n_6548),
.B(n_315),
.Y(n_6847)
);

OAI21xp33_ASAP7_75t_L g6848 ( 
.A1(n_6596),
.A2(n_6541),
.B(n_6693),
.Y(n_6848)
);

AOI221xp5_ASAP7_75t_L g6849 ( 
.A1(n_6600),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.C(n_320),
.Y(n_6849)
);

NAND2xp5_ASAP7_75t_SL g6850 ( 
.A(n_6715),
.B(n_317),
.Y(n_6850)
);

OAI22xp5_ASAP7_75t_L g6851 ( 
.A1(n_6691),
.A2(n_6542),
.B1(n_6607),
.B2(n_6695),
.Y(n_6851)
);

OAI221xp5_ASAP7_75t_SL g6852 ( 
.A1(n_6659),
.A2(n_324),
.B1(n_320),
.B2(n_322),
.C(n_325),
.Y(n_6852)
);

OA21x2_ASAP7_75t_L g6853 ( 
.A1(n_6544),
.A2(n_322),
.B(n_326),
.Y(n_6853)
);

NAND2xp5_ASAP7_75t_L g6854 ( 
.A(n_6637),
.B(n_326),
.Y(n_6854)
);

AND2x2_ASAP7_75t_L g6855 ( 
.A(n_6596),
.B(n_327),
.Y(n_6855)
);

AOI22xp33_ASAP7_75t_SL g6856 ( 
.A1(n_6691),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_6856)
);

NAND2xp5_ASAP7_75t_L g6857 ( 
.A(n_6697),
.B(n_330),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_L g6858 ( 
.A(n_6670),
.B(n_332),
.Y(n_6858)
);

NAND4xp25_ASAP7_75t_L g6859 ( 
.A(n_6584),
.B(n_335),
.C(n_333),
.D(n_334),
.Y(n_6859)
);

AND2x2_ASAP7_75t_L g6860 ( 
.A(n_6711),
.B(n_6609),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6609),
.B(n_333),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_L g6862 ( 
.A(n_6639),
.B(n_335),
.Y(n_6862)
);

OAI22xp5_ASAP7_75t_L g6863 ( 
.A1(n_6631),
.A2(n_339),
.B1(n_336),
.B2(n_337),
.Y(n_6863)
);

AND2x2_ASAP7_75t_L g6864 ( 
.A(n_6641),
.B(n_336),
.Y(n_6864)
);

NAND3xp33_ASAP7_75t_L g6865 ( 
.A(n_6603),
.B(n_337),
.C(n_339),
.Y(n_6865)
);

OAI21xp5_ASAP7_75t_L g6866 ( 
.A1(n_6696),
.A2(n_341),
.B(n_342),
.Y(n_6866)
);

OAI221xp5_ASAP7_75t_L g6867 ( 
.A1(n_6657),
.A2(n_344),
.B1(n_341),
.B2(n_342),
.C(n_345),
.Y(n_6867)
);

NAND3xp33_ASAP7_75t_L g6868 ( 
.A(n_6603),
.B(n_344),
.C(n_345),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_SL g6869 ( 
.A(n_6715),
.B(n_347),
.Y(n_6869)
);

NOR2xp33_ASAP7_75t_L g6870 ( 
.A(n_6571),
.B(n_348),
.Y(n_6870)
);

NAND2xp5_ASAP7_75t_L g6871 ( 
.A(n_6639),
.B(n_348),
.Y(n_6871)
);

NOR2xp33_ASAP7_75t_L g6872 ( 
.A(n_6571),
.B(n_349),
.Y(n_6872)
);

NOR2xp33_ASAP7_75t_L g6873 ( 
.A(n_6538),
.B(n_350),
.Y(n_6873)
);

NAND2xp5_ASAP7_75t_L g6874 ( 
.A(n_6639),
.B(n_351),
.Y(n_6874)
);

NAND2xp5_ASAP7_75t_L g6875 ( 
.A(n_6643),
.B(n_6620),
.Y(n_6875)
);

NAND2xp5_ASAP7_75t_L g6876 ( 
.A(n_6651),
.B(n_351),
.Y(n_6876)
);

OAI21xp5_ASAP7_75t_SL g6877 ( 
.A1(n_6566),
.A2(n_352),
.B(n_353),
.Y(n_6877)
);

AND2x2_ASAP7_75t_L g6878 ( 
.A(n_6601),
.B(n_353),
.Y(n_6878)
);

NAND2xp5_ASAP7_75t_L g6879 ( 
.A(n_6651),
.B(n_354),
.Y(n_6879)
);

NAND2xp5_ASAP7_75t_L g6880 ( 
.A(n_6651),
.B(n_354),
.Y(n_6880)
);

AND2x2_ASAP7_75t_L g6881 ( 
.A(n_6566),
.B(n_355),
.Y(n_6881)
);

NAND2xp5_ASAP7_75t_SL g6882 ( 
.A(n_6715),
.B(n_355),
.Y(n_6882)
);

OAI221xp5_ASAP7_75t_SL g6883 ( 
.A1(n_6659),
.A2(n_6687),
.B1(n_6657),
.B2(n_6677),
.C(n_6663),
.Y(n_6883)
);

NAND2xp5_ASAP7_75t_L g6884 ( 
.A(n_6652),
.B(n_356),
.Y(n_6884)
);

NAND2xp5_ASAP7_75t_L g6885 ( 
.A(n_6652),
.B(n_356),
.Y(n_6885)
);

NAND2xp5_ASAP7_75t_L g6886 ( 
.A(n_6652),
.B(n_357),
.Y(n_6886)
);

NAND2xp5_ASAP7_75t_L g6887 ( 
.A(n_6665),
.B(n_357),
.Y(n_6887)
);

NAND2xp5_ASAP7_75t_L g6888 ( 
.A(n_6665),
.B(n_358),
.Y(n_6888)
);

OAI22xp5_ASAP7_75t_L g6889 ( 
.A1(n_6630),
.A2(n_363),
.B1(n_359),
.B2(n_360),
.Y(n_6889)
);

NAND2xp5_ASAP7_75t_L g6890 ( 
.A(n_6706),
.B(n_360),
.Y(n_6890)
);

NAND3xp33_ASAP7_75t_L g6891 ( 
.A(n_6687),
.B(n_364),
.C(n_365),
.Y(n_6891)
);

NOR2xp33_ASAP7_75t_R g6892 ( 
.A(n_6538),
.B(n_6584),
.Y(n_6892)
);

OAI21xp33_ASAP7_75t_L g6893 ( 
.A1(n_6612),
.A2(n_364),
.B(n_366),
.Y(n_6893)
);

AND2x2_ASAP7_75t_L g6894 ( 
.A(n_6598),
.B(n_366),
.Y(n_6894)
);

NAND2xp5_ASAP7_75t_L g6895 ( 
.A(n_6706),
.B(n_368),
.Y(n_6895)
);

AND2x2_ASAP7_75t_L g6896 ( 
.A(n_6537),
.B(n_369),
.Y(n_6896)
);

OAI22xp5_ASAP7_75t_L g6897 ( 
.A1(n_6630),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_6897)
);

NAND2xp5_ASAP7_75t_L g6898 ( 
.A(n_6662),
.B(n_371),
.Y(n_6898)
);

NAND2xp5_ASAP7_75t_L g6899 ( 
.A(n_6553),
.B(n_373),
.Y(n_6899)
);

OAI21xp33_ASAP7_75t_SL g6900 ( 
.A1(n_6525),
.A2(n_373),
.B(n_374),
.Y(n_6900)
);

AND2x2_ASAP7_75t_L g6901 ( 
.A(n_6631),
.B(n_374),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_6649),
.B(n_375),
.Y(n_6902)
);

AND2x2_ASAP7_75t_L g6903 ( 
.A(n_6649),
.B(n_375),
.Y(n_6903)
);

NAND2xp5_ASAP7_75t_L g6904 ( 
.A(n_6553),
.B(n_377),
.Y(n_6904)
);

NAND3xp33_ASAP7_75t_L g6905 ( 
.A(n_6688),
.B(n_378),
.C(n_379),
.Y(n_6905)
);

OAI221xp5_ASAP7_75t_SL g6906 ( 
.A1(n_6677),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.C(n_382),
.Y(n_6906)
);

AND2x2_ASAP7_75t_L g6907 ( 
.A(n_6550),
.B(n_380),
.Y(n_6907)
);

NAND2xp5_ASAP7_75t_L g6908 ( 
.A(n_6555),
.B(n_383),
.Y(n_6908)
);

NAND2xp5_ASAP7_75t_SL g6909 ( 
.A(n_6578),
.B(n_6614),
.Y(n_6909)
);

NAND2xp5_ASAP7_75t_L g6910 ( 
.A(n_6555),
.B(n_384),
.Y(n_6910)
);

NAND2xp5_ASAP7_75t_L g6911 ( 
.A(n_6644),
.B(n_385),
.Y(n_6911)
);

OAI21xp33_ASAP7_75t_SL g6912 ( 
.A1(n_6642),
.A2(n_385),
.B(n_386),
.Y(n_6912)
);

AOI21xp33_ASAP7_75t_L g6913 ( 
.A1(n_6626),
.A2(n_387),
.B(n_388),
.Y(n_6913)
);

NAND2xp5_ASAP7_75t_L g6914 ( 
.A(n_6614),
.B(n_388),
.Y(n_6914)
);

NOR3xp33_ASAP7_75t_SL g6915 ( 
.A(n_6580),
.B(n_389),
.C(n_390),
.Y(n_6915)
);

OAI221xp5_ASAP7_75t_SL g6916 ( 
.A1(n_6663),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.C(n_393),
.Y(n_6916)
);

AND2x2_ASAP7_75t_L g6917 ( 
.A(n_6682),
.B(n_393),
.Y(n_6917)
);

AND2x2_ASAP7_75t_L g6918 ( 
.A(n_6524),
.B(n_6707),
.Y(n_6918)
);

OAI21xp33_ASAP7_75t_L g6919 ( 
.A1(n_6522),
.A2(n_394),
.B(n_395),
.Y(n_6919)
);

OAI22xp5_ASAP7_75t_L g6920 ( 
.A1(n_6688),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_6920)
);

NAND2xp5_ASAP7_75t_L g6921 ( 
.A(n_6614),
.B(n_396),
.Y(n_6921)
);

AND2x2_ASAP7_75t_L g6922 ( 
.A(n_6716),
.B(n_398),
.Y(n_6922)
);

NAND4xp25_ASAP7_75t_L g6923 ( 
.A(n_6655),
.B(n_400),
.C(n_398),
.D(n_399),
.Y(n_6923)
);

AND2x2_ASAP7_75t_L g6924 ( 
.A(n_6629),
.B(n_399),
.Y(n_6924)
);

NAND2xp5_ASAP7_75t_L g6925 ( 
.A(n_6627),
.B(n_400),
.Y(n_6925)
);

NAND3xp33_ASAP7_75t_L g6926 ( 
.A(n_6688),
.B(n_401),
.C(n_402),
.Y(n_6926)
);

NAND3xp33_ASAP7_75t_L g6927 ( 
.A(n_6688),
.B(n_401),
.C(n_403),
.Y(n_6927)
);

NAND2xp5_ASAP7_75t_SL g6928 ( 
.A(n_6578),
.B(n_404),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_L g6929 ( 
.A(n_6633),
.B(n_405),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6646),
.Y(n_6930)
);

OAI22xp5_ASAP7_75t_SL g6931 ( 
.A1(n_6714),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_6931)
);

INVx1_ASAP7_75t_SL g6932 ( 
.A(n_6752),
.Y(n_6932)
);

BUFx2_ASAP7_75t_L g6933 ( 
.A(n_6762),
.Y(n_6933)
);

BUFx3_ASAP7_75t_L g6934 ( 
.A(n_6759),
.Y(n_6934)
);

INVx1_ASAP7_75t_L g6935 ( 
.A(n_6841),
.Y(n_6935)
);

INVx2_ASAP7_75t_L g6936 ( 
.A(n_6763),
.Y(n_6936)
);

NAND2xp5_ASAP7_75t_L g6937 ( 
.A(n_6791),
.B(n_6692),
.Y(n_6937)
);

AND2x2_ASAP7_75t_L g6938 ( 
.A(n_6860),
.B(n_6608),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6838),
.Y(n_6939)
);

AND2x2_ASAP7_75t_L g6940 ( 
.A(n_6758),
.B(n_6699),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_6819),
.Y(n_6941)
);

NAND2xp5_ASAP7_75t_L g6942 ( 
.A(n_6912),
.B(n_6692),
.Y(n_6942)
);

INVx5_ASAP7_75t_SL g6943 ( 
.A(n_6892),
.Y(n_6943)
);

INVx2_ASAP7_75t_L g6944 ( 
.A(n_6765),
.Y(n_6944)
);

HB1xp67_ASAP7_75t_L g6945 ( 
.A(n_6814),
.Y(n_6945)
);

INVx1_ASAP7_75t_L g6946 ( 
.A(n_6821),
.Y(n_6946)
);

BUFx2_ASAP7_75t_L g6947 ( 
.A(n_6918),
.Y(n_6947)
);

AND2x2_ASAP7_75t_L g6948 ( 
.A(n_6778),
.B(n_6699),
.Y(n_6948)
);

AND2x2_ASAP7_75t_L g6949 ( 
.A(n_6780),
.B(n_6611),
.Y(n_6949)
);

AND2x2_ASAP7_75t_L g6950 ( 
.A(n_6784),
.B(n_6616),
.Y(n_6950)
);

INVx2_ASAP7_75t_L g6951 ( 
.A(n_6768),
.Y(n_6951)
);

OAI22xp5_ASAP7_75t_L g6952 ( 
.A1(n_6749),
.A2(n_6915),
.B1(n_6761),
.B2(n_6843),
.Y(n_6952)
);

INVx3_ASAP7_75t_L g6953 ( 
.A(n_6826),
.Y(n_6953)
);

NAND2xp5_ASAP7_75t_L g6954 ( 
.A(n_6877),
.B(n_6642),
.Y(n_6954)
);

OAI21xp33_ASAP7_75t_L g6955 ( 
.A1(n_6848),
.A2(n_6588),
.B(n_6604),
.Y(n_6955)
);

NOR2xp33_ASAP7_75t_L g6956 ( 
.A(n_6767),
.B(n_6653),
.Y(n_6956)
);

AND2x2_ASAP7_75t_L g6957 ( 
.A(n_6788),
.B(n_6632),
.Y(n_6957)
);

INVx1_ASAP7_75t_L g6958 ( 
.A(n_6914),
.Y(n_6958)
);

AND2x2_ASAP7_75t_L g6959 ( 
.A(n_6795),
.B(n_6622),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_6921),
.Y(n_6960)
);

BUFx3_ASAP7_75t_L g6961 ( 
.A(n_6829),
.Y(n_6961)
);

INVx2_ASAP7_75t_L g6962 ( 
.A(n_6853),
.Y(n_6962)
);

BUFx2_ASAP7_75t_L g6963 ( 
.A(n_6754),
.Y(n_6963)
);

AND2x4_ASAP7_75t_L g6964 ( 
.A(n_6861),
.B(n_6727),
.Y(n_6964)
);

OR2x2_ASAP7_75t_L g6965 ( 
.A(n_6875),
.B(n_6523),
.Y(n_6965)
);

INVx2_ASAP7_75t_L g6966 ( 
.A(n_6853),
.Y(n_6966)
);

OAI21xp33_ASAP7_75t_L g6967 ( 
.A1(n_6769),
.A2(n_6529),
.B(n_6606),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6835),
.B(n_6839),
.Y(n_6968)
);

AOI22xp5_ASAP7_75t_L g6969 ( 
.A1(n_6764),
.A2(n_6709),
.B1(n_6645),
.B2(n_6556),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6777),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6781),
.Y(n_6971)
);

NOR2xp33_ASAP7_75t_L g6972 ( 
.A(n_6767),
.B(n_6746),
.Y(n_6972)
);

NAND2xp5_ASAP7_75t_L g6973 ( 
.A(n_6889),
.B(n_6645),
.Y(n_6973)
);

AOI31xp33_ASAP7_75t_SL g6974 ( 
.A1(n_6753),
.A2(n_6552),
.A3(n_6573),
.B(n_6532),
.Y(n_6974)
);

NAND2xp5_ASAP7_75t_L g6975 ( 
.A(n_6889),
.B(n_6645),
.Y(n_6975)
);

AND2x4_ASAP7_75t_L g6976 ( 
.A(n_6878),
.B(n_6736),
.Y(n_6976)
);

AOI221xp5_ASAP7_75t_L g6977 ( 
.A1(n_6751),
.A2(n_6640),
.B1(n_6635),
.B2(n_6573),
.C(n_6615),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6842),
.Y(n_6978)
);

BUFx2_ASAP7_75t_L g6979 ( 
.A(n_6900),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_6844),
.Y(n_6980)
);

AND2x2_ASAP7_75t_L g6981 ( 
.A(n_6840),
.B(n_6592),
.Y(n_6981)
);

OAI221xp5_ASAP7_75t_L g6982 ( 
.A1(n_6816),
.A2(n_6673),
.B1(n_6669),
.B2(n_6732),
.C(n_6701),
.Y(n_6982)
);

NAND2xp5_ASAP7_75t_L g6983 ( 
.A(n_6897),
.B(n_6615),
.Y(n_6983)
);

OR2x2_ASAP7_75t_L g6984 ( 
.A(n_6818),
.B(n_6813),
.Y(n_6984)
);

NOR2xp67_ASAP7_75t_L g6985 ( 
.A(n_6831),
.B(n_6736),
.Y(n_6985)
);

INVx2_ASAP7_75t_L g6986 ( 
.A(n_6917),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6792),
.Y(n_6987)
);

NOR3xp33_ASAP7_75t_L g6988 ( 
.A(n_6931),
.B(n_6685),
.C(n_6668),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6887),
.Y(n_6989)
);

OAI21x1_ASAP7_75t_L g6990 ( 
.A1(n_6909),
.A2(n_6547),
.B(n_6544),
.Y(n_6990)
);

NAND3xp33_ASAP7_75t_L g6991 ( 
.A(n_6770),
.B(n_6547),
.C(n_6551),
.Y(n_6991)
);

BUFx2_ASAP7_75t_L g6992 ( 
.A(n_6881),
.Y(n_6992)
);

OR2x2_ASAP7_75t_L g6993 ( 
.A(n_6815),
.B(n_6597),
.Y(n_6993)
);

INVx2_ASAP7_75t_L g6994 ( 
.A(n_6864),
.Y(n_6994)
);

INVx2_ASAP7_75t_L g6995 ( 
.A(n_6922),
.Y(n_6995)
);

AND2x2_ASAP7_75t_L g6996 ( 
.A(n_6847),
.B(n_6718),
.Y(n_6996)
);

AND2x2_ASAP7_75t_L g6997 ( 
.A(n_6855),
.B(n_6718),
.Y(n_6997)
);

INVx2_ASAP7_75t_L g6998 ( 
.A(n_6896),
.Y(n_6998)
);

INVx1_ASAP7_75t_L g6999 ( 
.A(n_6888),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6890),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6895),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6873),
.B(n_6870),
.Y(n_7002)
);

NAND3xp33_ASAP7_75t_L g7003 ( 
.A(n_6897),
.B(n_6636),
.C(n_6551),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6782),
.Y(n_7004)
);

AND2x2_ASAP7_75t_L g7005 ( 
.A(n_6872),
.B(n_6557),
.Y(n_7005)
);

INVx1_ASAP7_75t_L g7006 ( 
.A(n_6898),
.Y(n_7006)
);

OAI33xp33_ASAP7_75t_L g7007 ( 
.A1(n_6851),
.A2(n_6741),
.A3(n_6636),
.B1(n_6648),
.B2(n_6532),
.B3(n_6539),
.Y(n_7007)
);

OAI33xp33_ASAP7_75t_L g7008 ( 
.A1(n_6851),
.A2(n_6648),
.A3(n_6539),
.B1(n_6528),
.B2(n_6562),
.B3(n_6567),
.Y(n_7008)
);

HB1xp67_ASAP7_75t_L g7009 ( 
.A(n_6836),
.Y(n_7009)
);

AOI33xp33_ASAP7_75t_L g7010 ( 
.A1(n_6856),
.A2(n_6528),
.A3(n_6702),
.B1(n_6569),
.B2(n_6574),
.B3(n_6564),
.Y(n_7010)
);

AND2x2_ASAP7_75t_L g7011 ( 
.A(n_6832),
.B(n_6740),
.Y(n_7011)
);

HB1xp67_ASAP7_75t_L g7012 ( 
.A(n_6836),
.Y(n_7012)
);

INVx2_ASAP7_75t_L g7013 ( 
.A(n_6894),
.Y(n_7013)
);

INVx4_ASAP7_75t_L g7014 ( 
.A(n_6901),
.Y(n_7014)
);

AND2x2_ASAP7_75t_L g7015 ( 
.A(n_6833),
.B(n_6740),
.Y(n_7015)
);

INVx1_ASAP7_75t_L g7016 ( 
.A(n_6930),
.Y(n_7016)
);

AND2x2_ASAP7_75t_L g7017 ( 
.A(n_6757),
.B(n_6728),
.Y(n_7017)
);

OR2x2_ASAP7_75t_L g7018 ( 
.A(n_6857),
.B(n_6613),
.Y(n_7018)
);

OAI21xp33_ASAP7_75t_SL g7019 ( 
.A1(n_6760),
.A2(n_6619),
.B(n_6579),
.Y(n_7019)
);

OAI211xp5_ASAP7_75t_SL g7020 ( 
.A1(n_6817),
.A2(n_6552),
.B(n_6747),
.C(n_6666),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6854),
.Y(n_7021)
);

INVx2_ASAP7_75t_L g7022 ( 
.A(n_6907),
.Y(n_7022)
);

AND2x2_ASAP7_75t_L g7023 ( 
.A(n_6902),
.B(n_6543),
.Y(n_7023)
);

INVx2_ASAP7_75t_L g7024 ( 
.A(n_6903),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6808),
.Y(n_7025)
);

INVx2_ASAP7_75t_SL g7026 ( 
.A(n_6924),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6899),
.Y(n_7027)
);

AND2x2_ASAP7_75t_L g7028 ( 
.A(n_6824),
.B(n_6543),
.Y(n_7028)
);

NOR2xp33_ASAP7_75t_L g7029 ( 
.A(n_6823),
.B(n_6683),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_6804),
.B(n_6543),
.Y(n_7030)
);

NAND2xp5_ASAP7_75t_SL g7031 ( 
.A(n_6837),
.B(n_6578),
.Y(n_7031)
);

AND2x2_ASAP7_75t_L g7032 ( 
.A(n_6806),
.B(n_6624),
.Y(n_7032)
);

AOI211xp5_ASAP7_75t_SL g7033 ( 
.A1(n_6802),
.A2(n_6720),
.B(n_6686),
.C(n_6731),
.Y(n_7033)
);

AND2x2_ASAP7_75t_L g7034 ( 
.A(n_6793),
.B(n_6625),
.Y(n_7034)
);

INVx2_ASAP7_75t_L g7035 ( 
.A(n_6776),
.Y(n_7035)
);

HB1xp67_ASAP7_75t_L g7036 ( 
.A(n_6793),
.Y(n_7036)
);

NAND2xp5_ASAP7_75t_L g7037 ( 
.A(n_6794),
.B(n_6830),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6904),
.Y(n_7038)
);

OAI221xp5_ASAP7_75t_L g7039 ( 
.A1(n_6794),
.A2(n_6673),
.B1(n_6669),
.B2(n_6721),
.C(n_6719),
.Y(n_7039)
);

AND2x2_ASAP7_75t_L g7040 ( 
.A(n_6925),
.B(n_6561),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6908),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_6910),
.Y(n_7042)
);

NAND2xp5_ASAP7_75t_L g7043 ( 
.A(n_6799),
.B(n_6667),
.Y(n_7043)
);

AND2x2_ASAP7_75t_L g7044 ( 
.A(n_6929),
.B(n_6556),
.Y(n_7044)
);

AND2x2_ASAP7_75t_L g7045 ( 
.A(n_6775),
.B(n_6556),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6911),
.Y(n_7046)
);

NOR2xp33_ASAP7_75t_L g7047 ( 
.A(n_6823),
.B(n_6683),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6797),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6796),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6858),
.Y(n_7050)
);

AND2x2_ASAP7_75t_L g7051 ( 
.A(n_6928),
.B(n_6589),
.Y(n_7051)
);

HB1xp67_ASAP7_75t_L g7052 ( 
.A(n_6805),
.Y(n_7052)
);

AND2x2_ASAP7_75t_L g7053 ( 
.A(n_6750),
.B(n_6559),
.Y(n_7053)
);

NAND2xp5_ASAP7_75t_SL g7054 ( 
.A(n_6785),
.B(n_6540),
.Y(n_7054)
);

AND2x2_ASAP7_75t_L g7055 ( 
.A(n_6827),
.B(n_6559),
.Y(n_7055)
);

INVx5_ASAP7_75t_L g7056 ( 
.A(n_6790),
.Y(n_7056)
);

NAND2xp5_ASAP7_75t_L g7057 ( 
.A(n_6789),
.B(n_6676),
.Y(n_7057)
);

INVx2_ASAP7_75t_L g7058 ( 
.A(n_6779),
.Y(n_7058)
);

AO21x2_ASAP7_75t_L g7059 ( 
.A1(n_6913),
.A2(n_6666),
.B(n_6664),
.Y(n_7059)
);

OR2x2_ASAP7_75t_L g7060 ( 
.A(n_6787),
.B(n_6766),
.Y(n_7060)
);

AND2x2_ASAP7_75t_L g7061 ( 
.A(n_6801),
.B(n_6811),
.Y(n_7061)
);

AND2x2_ASAP7_75t_L g7062 ( 
.A(n_6822),
.B(n_6560),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_L g7063 ( 
.A(n_6805),
.B(n_6680),
.Y(n_7063)
);

BUFx2_ASAP7_75t_L g7064 ( 
.A(n_6866),
.Y(n_7064)
);

OAI21xp5_ASAP7_75t_L g7065 ( 
.A1(n_6786),
.A2(n_6926),
.B(n_6905),
.Y(n_7065)
);

AOI211xp5_ASAP7_75t_L g7066 ( 
.A1(n_6883),
.A2(n_6575),
.B(n_6540),
.C(n_6618),
.Y(n_7066)
);

OAI221xp5_ASAP7_75t_L g7067 ( 
.A1(n_6786),
.A2(n_6748),
.B1(n_6739),
.B2(n_6705),
.C(n_6703),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_6876),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6879),
.Y(n_7069)
);

INVx1_ASAP7_75t_SL g7070 ( 
.A(n_6798),
.Y(n_7070)
);

AND2x2_ASAP7_75t_L g7071 ( 
.A(n_6850),
.B(n_6560),
.Y(n_7071)
);

AND2x2_ASAP7_75t_L g7072 ( 
.A(n_6869),
.B(n_6581),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6880),
.Y(n_7073)
);

NAND2xp5_ASAP7_75t_L g7074 ( 
.A(n_6845),
.B(n_6664),
.Y(n_7074)
);

AND2x2_ASAP7_75t_L g7075 ( 
.A(n_6940),
.B(n_6581),
.Y(n_7075)
);

NAND2xp5_ASAP7_75t_L g7076 ( 
.A(n_7036),
.B(n_6865),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_6945),
.Y(n_7077)
);

INVx2_ASAP7_75t_L g7078 ( 
.A(n_6934),
.Y(n_7078)
);

NOR2xp33_ASAP7_75t_L g7079 ( 
.A(n_7056),
.B(n_6771),
.Y(n_7079)
);

INVx2_ASAP7_75t_L g7080 ( 
.A(n_6961),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_7056),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_7036),
.B(n_6868),
.Y(n_7082)
);

AND2x2_ASAP7_75t_L g7083 ( 
.A(n_6933),
.B(n_6594),
.Y(n_7083)
);

OR2x2_ASAP7_75t_L g7084 ( 
.A(n_6932),
.B(n_6923),
.Y(n_7084)
);

AND2x2_ASAP7_75t_L g7085 ( 
.A(n_6943),
.B(n_6932),
.Y(n_7085)
);

INVx1_ASAP7_75t_SL g7086 ( 
.A(n_7056),
.Y(n_7086)
);

BUFx2_ASAP7_75t_L g7087 ( 
.A(n_6947),
.Y(n_7087)
);

NOR2xp33_ASAP7_75t_L g7088 ( 
.A(n_7056),
.B(n_6773),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_7064),
.B(n_6755),
.Y(n_7089)
);

NAND2x1p5_ASAP7_75t_L g7090 ( 
.A(n_6938),
.B(n_6882),
.Y(n_7090)
);

AND2x2_ASAP7_75t_L g7091 ( 
.A(n_6943),
.B(n_6594),
.Y(n_7091)
);

INVx1_ASAP7_75t_SL g7092 ( 
.A(n_6949),
.Y(n_7092)
);

AND2x4_ASAP7_75t_L g7093 ( 
.A(n_6964),
.B(n_6634),
.Y(n_7093)
);

HB1xp67_ASAP7_75t_L g7094 ( 
.A(n_6945),
.Y(n_7094)
);

INVx1_ASAP7_75t_SL g7095 ( 
.A(n_6950),
.Y(n_7095)
);

AND2x2_ASAP7_75t_L g7096 ( 
.A(n_6943),
.B(n_6602),
.Y(n_7096)
);

NAND2xp5_ASAP7_75t_L g7097 ( 
.A(n_7052),
.B(n_6979),
.Y(n_7097)
);

INVx2_ASAP7_75t_L g7098 ( 
.A(n_7052),
.Y(n_7098)
);

BUFx2_ASAP7_75t_L g7099 ( 
.A(n_6964),
.Y(n_7099)
);

NAND2xp5_ASAP7_75t_L g7100 ( 
.A(n_7009),
.B(n_6755),
.Y(n_7100)
);

OR2x2_ASAP7_75t_L g7101 ( 
.A(n_6942),
.B(n_6812),
.Y(n_7101)
);

INVx2_ASAP7_75t_L g7102 ( 
.A(n_6953),
.Y(n_7102)
);

AND2x2_ASAP7_75t_L g7103 ( 
.A(n_6948),
.B(n_6968),
.Y(n_7103)
);

INVx1_ASAP7_75t_SL g7104 ( 
.A(n_6992),
.Y(n_7104)
);

AND2x4_ASAP7_75t_L g7105 ( 
.A(n_6996),
.B(n_6884),
.Y(n_7105)
);

INVx2_ASAP7_75t_L g7106 ( 
.A(n_6953),
.Y(n_7106)
);

AND2x4_ASAP7_75t_L g7107 ( 
.A(n_6997),
.B(n_6885),
.Y(n_7107)
);

NAND2xp5_ASAP7_75t_L g7108 ( 
.A(n_7009),
.B(n_6893),
.Y(n_7108)
);

AND2x2_ASAP7_75t_L g7109 ( 
.A(n_7017),
.B(n_6602),
.Y(n_7109)
);

AND2x2_ASAP7_75t_L g7110 ( 
.A(n_6981),
.B(n_7028),
.Y(n_7110)
);

HB1xp67_ASAP7_75t_L g7111 ( 
.A(n_7012),
.Y(n_7111)
);

INVx1_ASAP7_75t_L g7112 ( 
.A(n_7012),
.Y(n_7112)
);

NAND2x1p5_ASAP7_75t_L g7113 ( 
.A(n_7054),
.B(n_6683),
.Y(n_7113)
);

INVx2_ASAP7_75t_L g7114 ( 
.A(n_6990),
.Y(n_7114)
);

NAND2xp5_ASAP7_75t_L g7115 ( 
.A(n_6983),
.B(n_6849),
.Y(n_7115)
);

AND3x2_ASAP7_75t_L g7116 ( 
.A(n_6972),
.B(n_6820),
.C(n_6800),
.Y(n_7116)
);

AND2x4_ASAP7_75t_L g7117 ( 
.A(n_7023),
.B(n_6886),
.Y(n_7117)
);

AND2x2_ASAP7_75t_L g7118 ( 
.A(n_7030),
.B(n_6610),
.Y(n_7118)
);

OR2x2_ASAP7_75t_SL g7119 ( 
.A(n_6942),
.B(n_6772),
.Y(n_7119)
);

AND2x2_ASAP7_75t_L g7120 ( 
.A(n_6963),
.B(n_6610),
.Y(n_7120)
);

AND2x2_ASAP7_75t_L g7121 ( 
.A(n_6936),
.B(n_6623),
.Y(n_7121)
);

INVx2_ASAP7_75t_L g7122 ( 
.A(n_6957),
.Y(n_7122)
);

BUFx2_ASAP7_75t_L g7123 ( 
.A(n_6976),
.Y(n_7123)
);

AND2x2_ASAP7_75t_L g7124 ( 
.A(n_6944),
.B(n_6623),
.Y(n_7124)
);

AND2x2_ASAP7_75t_L g7125 ( 
.A(n_6951),
.B(n_6540),
.Y(n_7125)
);

INVx1_ASAP7_75t_SL g7126 ( 
.A(n_7002),
.Y(n_7126)
);

AND2x4_ASAP7_75t_L g7127 ( 
.A(n_6976),
.B(n_6862),
.Y(n_7127)
);

INVx2_ASAP7_75t_SL g7128 ( 
.A(n_7026),
.Y(n_7128)
);

INVx2_ASAP7_75t_L g7129 ( 
.A(n_7014),
.Y(n_7129)
);

OR2x2_ASAP7_75t_L g7130 ( 
.A(n_6937),
.B(n_6859),
.Y(n_7130)
);

AND2x2_ASAP7_75t_L g7131 ( 
.A(n_7005),
.B(n_6733),
.Y(n_7131)
);

INVx2_ASAP7_75t_SL g7132 ( 
.A(n_7014),
.Y(n_7132)
);

BUFx2_ASAP7_75t_L g7133 ( 
.A(n_7035),
.Y(n_7133)
);

AND2x2_ASAP7_75t_L g7134 ( 
.A(n_7011),
.B(n_6565),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_7048),
.Y(n_7135)
);

NOR2xp67_ASAP7_75t_L g7136 ( 
.A(n_6956),
.B(n_6783),
.Y(n_7136)
);

OR2x2_ASAP7_75t_L g7137 ( 
.A(n_6937),
.B(n_6807),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_7004),
.Y(n_7138)
);

NOR2xp33_ASAP7_75t_L g7139 ( 
.A(n_7007),
.B(n_7008),
.Y(n_7139)
);

OR2x2_ASAP7_75t_L g7140 ( 
.A(n_6965),
.B(n_6828),
.Y(n_7140)
);

AND2x2_ASAP7_75t_L g7141 ( 
.A(n_7015),
.B(n_6846),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6998),
.Y(n_7142)
);

INVx2_ASAP7_75t_L g7143 ( 
.A(n_7013),
.Y(n_7143)
);

INVx3_ASAP7_75t_L g7144 ( 
.A(n_6994),
.Y(n_7144)
);

OR2x2_ASAP7_75t_L g7145 ( 
.A(n_6954),
.B(n_7060),
.Y(n_7145)
);

AND2x2_ASAP7_75t_L g7146 ( 
.A(n_7032),
.B(n_6730),
.Y(n_7146)
);

OR2x2_ASAP7_75t_L g7147 ( 
.A(n_6954),
.B(n_6828),
.Y(n_7147)
);

OR2x2_ASAP7_75t_L g7148 ( 
.A(n_6993),
.B(n_6871),
.Y(n_7148)
);

AND2x2_ASAP7_75t_L g7149 ( 
.A(n_7058),
.B(n_6730),
.Y(n_7149)
);

INVx2_ASAP7_75t_SL g7150 ( 
.A(n_7053),
.Y(n_7150)
);

AND2x2_ASAP7_75t_L g7151 ( 
.A(n_6956),
.B(n_6737),
.Y(n_7151)
);

NAND2xp5_ASAP7_75t_SL g7152 ( 
.A(n_7066),
.B(n_6920),
.Y(n_7152)
);

AND2x2_ASAP7_75t_L g7153 ( 
.A(n_6984),
.B(n_6737),
.Y(n_7153)
);

AND2x2_ASAP7_75t_L g7154 ( 
.A(n_7045),
.B(n_6618),
.Y(n_7154)
);

NAND2xp5_ASAP7_75t_L g7155 ( 
.A(n_6983),
.B(n_6920),
.Y(n_7155)
);

INVx3_ASAP7_75t_L g7156 ( 
.A(n_6986),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_L g7157 ( 
.A(n_6988),
.B(n_6874),
.Y(n_7157)
);

AND2x2_ASAP7_75t_L g7158 ( 
.A(n_7034),
.B(n_6618),
.Y(n_7158)
);

OR2x2_ASAP7_75t_L g7159 ( 
.A(n_7018),
.B(n_6852),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_7006),
.Y(n_7160)
);

AND2x2_ASAP7_75t_L g7161 ( 
.A(n_7061),
.B(n_7070),
.Y(n_7161)
);

AND2x2_ASAP7_75t_L g7162 ( 
.A(n_7070),
.B(n_6661),
.Y(n_7162)
);

HB1xp67_ASAP7_75t_L g7163 ( 
.A(n_6952),
.Y(n_7163)
);

INVx1_ASAP7_75t_SL g7164 ( 
.A(n_6972),
.Y(n_7164)
);

AND2x2_ASAP7_75t_SL g7165 ( 
.A(n_7037),
.B(n_6774),
.Y(n_7165)
);

INVx1_ASAP7_75t_L g7166 ( 
.A(n_7046),
.Y(n_7166)
);

OR2x2_ASAP7_75t_L g7167 ( 
.A(n_6935),
.B(n_6941),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6958),
.Y(n_7168)
);

AND2x2_ASAP7_75t_L g7169 ( 
.A(n_6959),
.B(n_6661),
.Y(n_7169)
);

AND2x2_ASAP7_75t_L g7170 ( 
.A(n_6995),
.B(n_6756),
.Y(n_7170)
);

AND2x2_ASAP7_75t_L g7171 ( 
.A(n_7010),
.B(n_6756),
.Y(n_7171)
);

AND2x2_ASAP7_75t_L g7172 ( 
.A(n_6985),
.B(n_6577),
.Y(n_7172)
);

NAND2xp5_ASAP7_75t_L g7173 ( 
.A(n_6988),
.B(n_6866),
.Y(n_7173)
);

AND2x2_ASAP7_75t_L g7174 ( 
.A(n_7071),
.B(n_6834),
.Y(n_7174)
);

CKINVDCx20_ASAP7_75t_R g7175 ( 
.A(n_7062),
.Y(n_7175)
);

AND2x2_ASAP7_75t_L g7176 ( 
.A(n_7072),
.B(n_6739),
.Y(n_7176)
);

NAND2x1p5_ASAP7_75t_L g7177 ( 
.A(n_6969),
.B(n_6575),
.Y(n_7177)
);

NAND2xp5_ASAP7_75t_SL g7178 ( 
.A(n_6952),
.B(n_7037),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_6960),
.Y(n_7179)
);

OR2x2_ASAP7_75t_L g7180 ( 
.A(n_6946),
.B(n_6546),
.Y(n_7180)
);

AND2x2_ASAP7_75t_L g7181 ( 
.A(n_6970),
.B(n_6748),
.Y(n_7181)
);

OR2x6_ASAP7_75t_L g7182 ( 
.A(n_7065),
.B(n_6800),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_L g7183 ( 
.A(n_7063),
.B(n_6919),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_7068),
.Y(n_7184)
);

NOR2x1p5_ASAP7_75t_L g7185 ( 
.A(n_7022),
.B(n_6927),
.Y(n_7185)
);

AND2x2_ASAP7_75t_L g7186 ( 
.A(n_6971),
.B(n_6595),
.Y(n_7186)
);

INVx2_ASAP7_75t_L g7187 ( 
.A(n_6962),
.Y(n_7187)
);

INVx1_ASAP7_75t_L g7188 ( 
.A(n_7069),
.Y(n_7188)
);

OR2x2_ASAP7_75t_L g7189 ( 
.A(n_7073),
.B(n_6939),
.Y(n_7189)
);

AND2x2_ASAP7_75t_L g7190 ( 
.A(n_7019),
.B(n_6595),
.Y(n_7190)
);

INVxp67_ASAP7_75t_L g7191 ( 
.A(n_7029),
.Y(n_7191)
);

INVx2_ASAP7_75t_L g7192 ( 
.A(n_6966),
.Y(n_7192)
);

INVxp67_ASAP7_75t_L g7193 ( 
.A(n_7047),
.Y(n_7193)
);

AND2x4_ASAP7_75t_L g7194 ( 
.A(n_7024),
.B(n_6684),
.Y(n_7194)
);

AND2x4_ASAP7_75t_L g7195 ( 
.A(n_7055),
.B(n_6684),
.Y(n_7195)
);

BUFx2_ASAP7_75t_L g7196 ( 
.A(n_7044),
.Y(n_7196)
);

INVx2_ASAP7_75t_L g7197 ( 
.A(n_7051),
.Y(n_7197)
);

AND2x2_ASAP7_75t_L g7198 ( 
.A(n_7040),
.B(n_6700),
.Y(n_7198)
);

HB1xp67_ASAP7_75t_L g7199 ( 
.A(n_7063),
.Y(n_7199)
);

INVx2_ASAP7_75t_L g7200 ( 
.A(n_7050),
.Y(n_7200)
);

AND2x2_ASAP7_75t_L g7201 ( 
.A(n_7033),
.B(n_7016),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6987),
.Y(n_7202)
);

AND2x2_ASAP7_75t_L g7203 ( 
.A(n_7033),
.B(n_6700),
.Y(n_7203)
);

AND2x4_ASAP7_75t_L g7204 ( 
.A(n_6989),
.B(n_6575),
.Y(n_7204)
);

AND2x2_ASAP7_75t_L g7205 ( 
.A(n_6999),
.B(n_6820),
.Y(n_7205)
);

OR2x2_ASAP7_75t_L g7206 ( 
.A(n_7000),
.B(n_6563),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_6978),
.Y(n_7207)
);

OR2x2_ASAP7_75t_L g7208 ( 
.A(n_7001),
.B(n_6980),
.Y(n_7208)
);

AND2x2_ASAP7_75t_L g7209 ( 
.A(n_7031),
.B(n_6621),
.Y(n_7209)
);

INVx6_ASAP7_75t_L g7210 ( 
.A(n_6974),
.Y(n_7210)
);

HB1xp67_ASAP7_75t_L g7211 ( 
.A(n_7043),
.Y(n_7211)
);

HB1xp67_ASAP7_75t_L g7212 ( 
.A(n_7043),
.Y(n_7212)
);

HB1xp67_ASAP7_75t_L g7213 ( 
.A(n_7111),
.Y(n_7213)
);

AND2x2_ASAP7_75t_L g7214 ( 
.A(n_7085),
.B(n_6955),
.Y(n_7214)
);

AND2x2_ASAP7_75t_L g7215 ( 
.A(n_7092),
.B(n_7027),
.Y(n_7215)
);

AND2x2_ASAP7_75t_L g7216 ( 
.A(n_7092),
.B(n_7038),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_7111),
.Y(n_7217)
);

AND2x2_ASAP7_75t_L g7218 ( 
.A(n_7095),
.B(n_7041),
.Y(n_7218)
);

INVx2_ASAP7_75t_SL g7219 ( 
.A(n_7083),
.Y(n_7219)
);

INVx2_ASAP7_75t_L g7220 ( 
.A(n_7175),
.Y(n_7220)
);

INVx1_ASAP7_75t_L g7221 ( 
.A(n_7087),
.Y(n_7221)
);

INVx2_ASAP7_75t_L g7222 ( 
.A(n_7175),
.Y(n_7222)
);

OR2x2_ASAP7_75t_L g7223 ( 
.A(n_7126),
.B(n_6991),
.Y(n_7223)
);

AND2x2_ASAP7_75t_L g7224 ( 
.A(n_7095),
.B(n_7042),
.Y(n_7224)
);

NAND2xp5_ASAP7_75t_L g7225 ( 
.A(n_7139),
.B(n_6977),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_7094),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_7094),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_7196),
.Y(n_7228)
);

INVx1_ASAP7_75t_L g7229 ( 
.A(n_7098),
.Y(n_7229)
);

NAND2xp5_ASAP7_75t_L g7230 ( 
.A(n_7139),
.B(n_6977),
.Y(n_7230)
);

NOR2xp33_ASAP7_75t_L g7231 ( 
.A(n_7086),
.B(n_7020),
.Y(n_7231)
);

NAND2xp5_ASAP7_75t_L g7232 ( 
.A(n_7199),
.B(n_7098),
.Y(n_7232)
);

NOR2xp33_ASAP7_75t_L g7233 ( 
.A(n_7086),
.B(n_7020),
.Y(n_7233)
);

NAND4xp25_ASAP7_75t_L g7234 ( 
.A(n_7097),
.B(n_6967),
.C(n_7067),
.D(n_6974),
.Y(n_7234)
);

INVx1_ASAP7_75t_SL g7235 ( 
.A(n_7210),
.Y(n_7235)
);

AND2x2_ASAP7_75t_L g7236 ( 
.A(n_7103),
.B(n_7099),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_7162),
.Y(n_7237)
);

NAND2xp5_ASAP7_75t_L g7238 ( 
.A(n_7199),
.B(n_6973),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_7123),
.B(n_7021),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_7120),
.Y(n_7240)
);

NOR2xp33_ASAP7_75t_L g7241 ( 
.A(n_7081),
.B(n_7007),
.Y(n_7241)
);

HB1xp67_ASAP7_75t_L g7242 ( 
.A(n_7081),
.Y(n_7242)
);

OAI221xp5_ASAP7_75t_L g7243 ( 
.A1(n_7100),
.A2(n_6975),
.B1(n_6973),
.B2(n_7065),
.C(n_7039),
.Y(n_7243)
);

OAI22xp33_ASAP7_75t_L g7244 ( 
.A1(n_7089),
.A2(n_6975),
.B1(n_7039),
.B2(n_6982),
.Y(n_7244)
);

INVx2_ASAP7_75t_L g7245 ( 
.A(n_7169),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_7126),
.Y(n_7246)
);

BUFx2_ASAP7_75t_L g7247 ( 
.A(n_7090),
.Y(n_7247)
);

BUFx2_ASAP7_75t_L g7248 ( 
.A(n_7090),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_7100),
.Y(n_7249)
);

INVx1_ASAP7_75t_SL g7250 ( 
.A(n_7210),
.Y(n_7250)
);

INVx1_ASAP7_75t_SL g7251 ( 
.A(n_7210),
.Y(n_7251)
);

NAND2xp5_ASAP7_75t_L g7252 ( 
.A(n_7163),
.B(n_7057),
.Y(n_7252)
);

AND2x2_ASAP7_75t_L g7253 ( 
.A(n_7075),
.B(n_7025),
.Y(n_7253)
);

BUFx2_ASAP7_75t_L g7254 ( 
.A(n_7113),
.Y(n_7254)
);

AND2x2_ASAP7_75t_L g7255 ( 
.A(n_7091),
.B(n_7096),
.Y(n_7255)
);

AND2x2_ASAP7_75t_L g7256 ( 
.A(n_7110),
.B(n_7049),
.Y(n_7256)
);

OR2x2_ASAP7_75t_L g7257 ( 
.A(n_7104),
.B(n_7057),
.Y(n_7257)
);

AND2x2_ASAP7_75t_L g7258 ( 
.A(n_7150),
.B(n_7074),
.Y(n_7258)
);

AND2x4_ASAP7_75t_L g7259 ( 
.A(n_7093),
.B(n_7003),
.Y(n_7259)
);

NAND2xp5_ASAP7_75t_L g7260 ( 
.A(n_7163),
.B(n_7074),
.Y(n_7260)
);

INVxp67_ASAP7_75t_L g7261 ( 
.A(n_7088),
.Y(n_7261)
);

OR2x2_ASAP7_75t_L g7262 ( 
.A(n_7104),
.B(n_7067),
.Y(n_7262)
);

NAND4xp25_ASAP7_75t_SL g7263 ( 
.A(n_7173),
.B(n_6982),
.C(n_6825),
.D(n_7008),
.Y(n_7263)
);

INVx1_ASAP7_75t_SL g7264 ( 
.A(n_7097),
.Y(n_7264)
);

AND2x2_ASAP7_75t_L g7265 ( 
.A(n_7133),
.B(n_7059),
.Y(n_7265)
);

INVx1_ASAP7_75t_SL g7266 ( 
.A(n_7164),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_7113),
.Y(n_7267)
);

NOR2xp33_ASAP7_75t_L g7268 ( 
.A(n_7164),
.B(n_7154),
.Y(n_7268)
);

CKINVDCx5p33_ASAP7_75t_R g7269 ( 
.A(n_7088),
.Y(n_7269)
);

AND2x2_ASAP7_75t_L g7270 ( 
.A(n_7078),
.B(n_7059),
.Y(n_7270)
);

OR2x2_ASAP7_75t_L g7271 ( 
.A(n_7178),
.B(n_6724),
.Y(n_7271)
);

INVx3_ASAP7_75t_L g7272 ( 
.A(n_7093),
.Y(n_7272)
);

AND2x4_ASAP7_75t_SL g7273 ( 
.A(n_7080),
.B(n_6704),
.Y(n_7273)
);

NAND2xp5_ASAP7_75t_L g7274 ( 
.A(n_7178),
.B(n_6724),
.Y(n_7274)
);

AND2x2_ASAP7_75t_L g7275 ( 
.A(n_7122),
.B(n_6724),
.Y(n_7275)
);

INVx2_ASAP7_75t_L g7276 ( 
.A(n_7151),
.Y(n_7276)
);

INVx2_ASAP7_75t_L g7277 ( 
.A(n_7131),
.Y(n_7277)
);

AND2x4_ASAP7_75t_L g7278 ( 
.A(n_7124),
.B(n_6712),
.Y(n_7278)
);

HB1xp67_ASAP7_75t_L g7279 ( 
.A(n_7136),
.Y(n_7279)
);

NAND2xp5_ASAP7_75t_L g7280 ( 
.A(n_7165),
.B(n_6803),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_7153),
.Y(n_7281)
);

INVx1_ASAP7_75t_L g7282 ( 
.A(n_7112),
.Y(n_7282)
);

AND2x2_ASAP7_75t_L g7283 ( 
.A(n_7190),
.B(n_6621),
.Y(n_7283)
);

NAND2xp5_ASAP7_75t_L g7284 ( 
.A(n_7173),
.B(n_6809),
.Y(n_7284)
);

INVx2_ASAP7_75t_L g7285 ( 
.A(n_7141),
.Y(n_7285)
);

AND2x4_ASAP7_75t_L g7286 ( 
.A(n_7121),
.B(n_7144),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_7176),
.Y(n_7287)
);

NAND2xp5_ASAP7_75t_L g7288 ( 
.A(n_7211),
.B(n_6810),
.Y(n_7288)
);

AND2x2_ASAP7_75t_L g7289 ( 
.A(n_7201),
.B(n_7125),
.Y(n_7289)
);

AND2x2_ASAP7_75t_L g7290 ( 
.A(n_7172),
.B(n_7128),
.Y(n_7290)
);

NAND2xp5_ASAP7_75t_L g7291 ( 
.A(n_7211),
.B(n_6863),
.Y(n_7291)
);

AND2x2_ASAP7_75t_L g7292 ( 
.A(n_7109),
.B(n_6621),
.Y(n_7292)
);

NAND2xp5_ASAP7_75t_L g7293 ( 
.A(n_7212),
.B(n_6891),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_7144),
.Y(n_7294)
);

HB1xp67_ASAP7_75t_L g7295 ( 
.A(n_7158),
.Y(n_7295)
);

AND2x2_ASAP7_75t_L g7296 ( 
.A(n_7197),
.B(n_6712),
.Y(n_7296)
);

AND2x2_ASAP7_75t_L g7297 ( 
.A(n_7132),
.B(n_6722),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_7156),
.Y(n_7298)
);

NAND2xp5_ASAP7_75t_L g7299 ( 
.A(n_7165),
.B(n_6722),
.Y(n_7299)
);

NAND2xp5_ASAP7_75t_L g7300 ( 
.A(n_7212),
.B(n_6626),
.Y(n_7300)
);

INVx2_ASAP7_75t_L g7301 ( 
.A(n_7134),
.Y(n_7301)
);

AND2x2_ASAP7_75t_L g7302 ( 
.A(n_7102),
.B(n_6675),
.Y(n_7302)
);

AND2x2_ASAP7_75t_L g7303 ( 
.A(n_7106),
.B(n_6534),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_7156),
.Y(n_7304)
);

AND2x2_ASAP7_75t_L g7305 ( 
.A(n_7129),
.B(n_6534),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_7089),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7148),
.Y(n_7307)
);

AND2x4_ASAP7_75t_L g7308 ( 
.A(n_7127),
.B(n_6534),
.Y(n_7308)
);

INVxp67_ASAP7_75t_L g7309 ( 
.A(n_7079),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_7187),
.Y(n_7310)
);

AND2x4_ASAP7_75t_L g7311 ( 
.A(n_7127),
.B(n_6916),
.Y(n_7311)
);

INVx2_ASAP7_75t_SL g7312 ( 
.A(n_7149),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_7192),
.Y(n_7313)
);

AND2x4_ASAP7_75t_L g7314 ( 
.A(n_7195),
.B(n_406),
.Y(n_7314)
);

INVx5_ASAP7_75t_L g7315 ( 
.A(n_7182),
.Y(n_7315)
);

AND2x4_ASAP7_75t_L g7316 ( 
.A(n_7195),
.B(n_407),
.Y(n_7316)
);

INVx1_ASAP7_75t_SL g7317 ( 
.A(n_7161),
.Y(n_7317)
);

INVxp67_ASAP7_75t_SL g7318 ( 
.A(n_7177),
.Y(n_7318)
);

INVx1_ASAP7_75t_SL g7319 ( 
.A(n_7119),
.Y(n_7319)
);

AND2x2_ASAP7_75t_L g7320 ( 
.A(n_7118),
.B(n_408),
.Y(n_7320)
);

INVx2_ASAP7_75t_L g7321 ( 
.A(n_7198),
.Y(n_7321)
);

OR2x2_ASAP7_75t_L g7322 ( 
.A(n_7145),
.B(n_6906),
.Y(n_7322)
);

AND2x2_ASAP7_75t_L g7323 ( 
.A(n_7186),
.B(n_409),
.Y(n_7323)
);

NAND2xp5_ASAP7_75t_L g7324 ( 
.A(n_7116),
.B(n_6867),
.Y(n_7324)
);

AND2x2_ASAP7_75t_L g7325 ( 
.A(n_7105),
.B(n_409),
.Y(n_7325)
);

INVx2_ASAP7_75t_SL g7326 ( 
.A(n_7105),
.Y(n_7326)
);

AND2x2_ASAP7_75t_L g7327 ( 
.A(n_7107),
.B(n_410),
.Y(n_7327)
);

AND2x2_ASAP7_75t_L g7328 ( 
.A(n_7107),
.B(n_410),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_7182),
.Y(n_7329)
);

INVx1_ASAP7_75t_L g7330 ( 
.A(n_7182),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_7077),
.Y(n_7331)
);

AND2x4_ASAP7_75t_L g7332 ( 
.A(n_7220),
.B(n_7117),
.Y(n_7332)
);

AO221x2_ASAP7_75t_L g7333 ( 
.A1(n_7222),
.A2(n_7157),
.B1(n_7155),
.B2(n_7115),
.C(n_7135),
.Y(n_7333)
);

OAI22xp33_ASAP7_75t_L g7334 ( 
.A1(n_7225),
.A2(n_7108),
.B1(n_7177),
.B2(n_7101),
.Y(n_7334)
);

NAND2xp5_ASAP7_75t_SL g7335 ( 
.A(n_7286),
.B(n_7117),
.Y(n_7335)
);

NAND2xp33_ASAP7_75t_SL g7336 ( 
.A(n_7236),
.B(n_7130),
.Y(n_7336)
);

AO221x2_ASAP7_75t_L g7337 ( 
.A1(n_7228),
.A2(n_7157),
.B1(n_7155),
.B2(n_7115),
.C(n_7138),
.Y(n_7337)
);

NAND2xp5_ASAP7_75t_L g7338 ( 
.A(n_7317),
.B(n_7116),
.Y(n_7338)
);

AO221x2_ASAP7_75t_L g7339 ( 
.A1(n_7246),
.A2(n_7166),
.B1(n_7160),
.B2(n_7179),
.C(n_7168),
.Y(n_7339)
);

NAND2xp5_ASAP7_75t_L g7340 ( 
.A(n_7317),
.B(n_7146),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_7295),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7286),
.B(n_7209),
.Y(n_7342)
);

NOR2xp33_ASAP7_75t_L g7343 ( 
.A(n_7269),
.B(n_7191),
.Y(n_7343)
);

NOR2x1_ASAP7_75t_L g7344 ( 
.A(n_7234),
.B(n_7079),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_7255),
.B(n_7203),
.Y(n_7345)
);

CKINVDCx20_ASAP7_75t_R g7346 ( 
.A(n_7273),
.Y(n_7346)
);

AND2x4_ASAP7_75t_L g7347 ( 
.A(n_7326),
.B(n_7142),
.Y(n_7347)
);

AND2x4_ASAP7_75t_L g7348 ( 
.A(n_7312),
.B(n_7272),
.Y(n_7348)
);

NAND2xp5_ASAP7_75t_L g7349 ( 
.A(n_7315),
.B(n_7292),
.Y(n_7349)
);

AO221x2_ASAP7_75t_L g7350 ( 
.A1(n_7225),
.A2(n_7230),
.B1(n_7221),
.B2(n_7301),
.C(n_7277),
.Y(n_7350)
);

AOI22xp5_ASAP7_75t_L g7351 ( 
.A1(n_7230),
.A2(n_7108),
.B1(n_7183),
.B2(n_7152),
.Y(n_7351)
);

NAND2xp5_ASAP7_75t_L g7352 ( 
.A(n_7315),
.B(n_7205),
.Y(n_7352)
);

INVx2_ASAP7_75t_SL g7353 ( 
.A(n_7272),
.Y(n_7353)
);

NOR4xp25_ASAP7_75t_SL g7354 ( 
.A(n_7247),
.B(n_7152),
.C(n_7188),
.D(n_7184),
.Y(n_7354)
);

CKINVDCx5p33_ASAP7_75t_R g7355 ( 
.A(n_7319),
.Y(n_7355)
);

OAI22xp33_ASAP7_75t_L g7356 ( 
.A1(n_7252),
.A2(n_7183),
.B1(n_7082),
.B2(n_7076),
.Y(n_7356)
);

INVx2_ASAP7_75t_L g7357 ( 
.A(n_7315),
.Y(n_7357)
);

NAND2xp5_ASAP7_75t_L g7358 ( 
.A(n_7268),
.B(n_7170),
.Y(n_7358)
);

INVxp33_ASAP7_75t_SL g7359 ( 
.A(n_7279),
.Y(n_7359)
);

NAND2xp5_ASAP7_75t_L g7360 ( 
.A(n_7319),
.B(n_7174),
.Y(n_7360)
);

OR2x2_ASAP7_75t_L g7361 ( 
.A(n_7266),
.B(n_7084),
.Y(n_7361)
);

NOR2x1_ASAP7_75t_L g7362 ( 
.A(n_7234),
.B(n_7137),
.Y(n_7362)
);

NAND2xp5_ASAP7_75t_L g7363 ( 
.A(n_7266),
.B(n_7181),
.Y(n_7363)
);

INVxp67_ASAP7_75t_L g7364 ( 
.A(n_7248),
.Y(n_7364)
);

OAI22xp33_ASAP7_75t_L g7365 ( 
.A1(n_7252),
.A2(n_7082),
.B1(n_7076),
.B2(n_7147),
.Y(n_7365)
);

NAND2xp5_ASAP7_75t_L g7366 ( 
.A(n_7314),
.B(n_7191),
.Y(n_7366)
);

NOR2xp33_ASAP7_75t_L g7367 ( 
.A(n_7280),
.B(n_7193),
.Y(n_7367)
);

NAND2xp33_ASAP7_75t_SL g7368 ( 
.A(n_7219),
.B(n_7189),
.Y(n_7368)
);

NAND2xp5_ASAP7_75t_L g7369 ( 
.A(n_7314),
.B(n_7193),
.Y(n_7369)
);

OR2x2_ASAP7_75t_L g7370 ( 
.A(n_7262),
.B(n_7140),
.Y(n_7370)
);

AO221x2_ASAP7_75t_L g7371 ( 
.A1(n_7240),
.A2(n_7207),
.B1(n_7202),
.B2(n_7143),
.C(n_7200),
.Y(n_7371)
);

AND2x4_ASAP7_75t_L g7372 ( 
.A(n_7245),
.B(n_7204),
.Y(n_7372)
);

AOI22xp5_ASAP7_75t_L g7373 ( 
.A1(n_7243),
.A2(n_7171),
.B1(n_7114),
.B2(n_7185),
.Y(n_7373)
);

NAND2xp5_ASAP7_75t_L g7374 ( 
.A(n_7316),
.B(n_7204),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_7316),
.B(n_7194),
.Y(n_7375)
);

NAND2xp5_ASAP7_75t_SL g7376 ( 
.A(n_7259),
.B(n_7159),
.Y(n_7376)
);

OR2x2_ASAP7_75t_L g7377 ( 
.A(n_7223),
.B(n_7180),
.Y(n_7377)
);

INVx2_ASAP7_75t_L g7378 ( 
.A(n_7254),
.Y(n_7378)
);

NAND2xp5_ASAP7_75t_L g7379 ( 
.A(n_7320),
.B(n_7285),
.Y(n_7379)
);

AND2x2_ASAP7_75t_L g7380 ( 
.A(n_7289),
.B(n_7194),
.Y(n_7380)
);

AO221x2_ASAP7_75t_L g7381 ( 
.A1(n_7237),
.A2(n_7114),
.B1(n_7167),
.B2(n_7208),
.C(n_7206),
.Y(n_7381)
);

NAND2xp5_ASAP7_75t_L g7382 ( 
.A(n_7325),
.B(n_7327),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_7242),
.Y(n_7383)
);

NOR2x1_ASAP7_75t_L g7384 ( 
.A(n_7260),
.B(n_411),
.Y(n_7384)
);

NAND2xp5_ASAP7_75t_L g7385 ( 
.A(n_7328),
.B(n_412),
.Y(n_7385)
);

AND2x2_ASAP7_75t_L g7386 ( 
.A(n_7290),
.B(n_412),
.Y(n_7386)
);

AOI22xp5_ASAP7_75t_L g7387 ( 
.A1(n_7263),
.A2(n_7241),
.B1(n_7244),
.B2(n_7238),
.Y(n_7387)
);

AND2x4_ASAP7_75t_L g7388 ( 
.A(n_7308),
.B(n_413),
.Y(n_7388)
);

NOR2xp33_ASAP7_75t_L g7389 ( 
.A(n_7261),
.B(n_415),
.Y(n_7389)
);

NOR2xp33_ASAP7_75t_L g7390 ( 
.A(n_7309),
.B(n_417),
.Y(n_7390)
);

INVxp33_ASAP7_75t_SL g7391 ( 
.A(n_7260),
.Y(n_7391)
);

NAND2xp33_ASAP7_75t_L g7392 ( 
.A(n_7257),
.B(n_417),
.Y(n_7392)
);

INVx2_ASAP7_75t_SL g7393 ( 
.A(n_7308),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_7311),
.B(n_418),
.Y(n_7394)
);

CKINVDCx5p33_ASAP7_75t_R g7395 ( 
.A(n_7323),
.Y(n_7395)
);

INVx2_ASAP7_75t_SL g7396 ( 
.A(n_7303),
.Y(n_7396)
);

INVxp33_ASAP7_75t_SL g7397 ( 
.A(n_7231),
.Y(n_7397)
);

NAND2xp33_ASAP7_75t_SL g7398 ( 
.A(n_7239),
.B(n_419),
.Y(n_7398)
);

NAND2xp33_ASAP7_75t_SL g7399 ( 
.A(n_7215),
.B(n_7216),
.Y(n_7399)
);

NOR2xp33_ASAP7_75t_SL g7400 ( 
.A(n_7287),
.B(n_419),
.Y(n_7400)
);

AO221x2_ASAP7_75t_L g7401 ( 
.A1(n_7232),
.A2(n_420),
.B1(n_421),
.B2(n_422),
.C(n_423),
.Y(n_7401)
);

AOI22xp5_ASAP7_75t_L g7402 ( 
.A1(n_7238),
.A2(n_425),
.B1(n_421),
.B2(n_423),
.Y(n_7402)
);

OAI221xp5_ASAP7_75t_L g7403 ( 
.A1(n_7274),
.A2(n_425),
.B1(n_426),
.B2(n_427),
.C(n_430),
.Y(n_7403)
);

NOR2xp33_ASAP7_75t_L g7404 ( 
.A(n_7271),
.B(n_426),
.Y(n_7404)
);

NAND2xp5_ASAP7_75t_L g7405 ( 
.A(n_7311),
.B(n_427),
.Y(n_7405)
);

OAI221xp5_ASAP7_75t_L g7406 ( 
.A1(n_7274),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.C(n_434),
.Y(n_7406)
);

AO221x2_ASAP7_75t_L g7407 ( 
.A1(n_7232),
.A2(n_431),
.B1(n_433),
.B2(n_434),
.C(n_438),
.Y(n_7407)
);

NAND2xp33_ASAP7_75t_SL g7408 ( 
.A(n_7218),
.B(n_438),
.Y(n_7408)
);

NOR2x1_ASAP7_75t_L g7409 ( 
.A(n_7264),
.B(n_439),
.Y(n_7409)
);

NAND2xp5_ASAP7_75t_L g7410 ( 
.A(n_7253),
.B(n_439),
.Y(n_7410)
);

NAND2xp5_ASAP7_75t_L g7411 ( 
.A(n_7259),
.B(n_440),
.Y(n_7411)
);

AOI22xp5_ASAP7_75t_L g7412 ( 
.A1(n_7306),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_7412)
);

NOR2x1_ASAP7_75t_L g7413 ( 
.A(n_7264),
.B(n_441),
.Y(n_7413)
);

NAND2xp33_ASAP7_75t_SL g7414 ( 
.A(n_7224),
.B(n_443),
.Y(n_7414)
);

AO221x2_ASAP7_75t_L g7415 ( 
.A1(n_7249),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.C(n_447),
.Y(n_7415)
);

NAND2xp5_ASAP7_75t_L g7416 ( 
.A(n_7256),
.B(n_444),
.Y(n_7416)
);

AND2x2_ASAP7_75t_L g7417 ( 
.A(n_7321),
.B(n_445),
.Y(n_7417)
);

CKINVDCx20_ASAP7_75t_R g7418 ( 
.A(n_7283),
.Y(n_7418)
);

NAND2xp5_ASAP7_75t_L g7419 ( 
.A(n_7278),
.B(n_449),
.Y(n_7419)
);

AND2x2_ASAP7_75t_L g7420 ( 
.A(n_7380),
.B(n_7258),
.Y(n_7420)
);

INVx5_ASAP7_75t_SL g7421 ( 
.A(n_7357),
.Y(n_7421)
);

HB1xp67_ASAP7_75t_L g7422 ( 
.A(n_7355),
.Y(n_7422)
);

INVx2_ASAP7_75t_L g7423 ( 
.A(n_7418),
.Y(n_7423)
);

AND2x2_ASAP7_75t_L g7424 ( 
.A(n_7345),
.B(n_7318),
.Y(n_7424)
);

OAI22xp5_ASAP7_75t_L g7425 ( 
.A1(n_7387),
.A2(n_7250),
.B1(n_7251),
.B2(n_7235),
.Y(n_7425)
);

NAND2xp5_ASAP7_75t_L g7426 ( 
.A(n_7333),
.B(n_7265),
.Y(n_7426)
);

INVxp67_ASAP7_75t_L g7427 ( 
.A(n_7409),
.Y(n_7427)
);

AND2x2_ASAP7_75t_L g7428 ( 
.A(n_7386),
.B(n_7214),
.Y(n_7428)
);

INVx1_ASAP7_75t_L g7429 ( 
.A(n_7340),
.Y(n_7429)
);

INVx1_ASAP7_75t_SL g7430 ( 
.A(n_7346),
.Y(n_7430)
);

INVx2_ASAP7_75t_L g7431 ( 
.A(n_7395),
.Y(n_7431)
);

OR2x2_ASAP7_75t_L g7432 ( 
.A(n_7350),
.B(n_7281),
.Y(n_7432)
);

AND2x2_ASAP7_75t_L g7433 ( 
.A(n_7350),
.B(n_7305),
.Y(n_7433)
);

OR2x2_ASAP7_75t_L g7434 ( 
.A(n_7333),
.B(n_7294),
.Y(n_7434)
);

OAI21xp33_ASAP7_75t_L g7435 ( 
.A1(n_7362),
.A2(n_7233),
.B(n_7324),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_7363),
.Y(n_7436)
);

INVxp67_ASAP7_75t_L g7437 ( 
.A(n_7413),
.Y(n_7437)
);

INVx2_ASAP7_75t_SL g7438 ( 
.A(n_7348),
.Y(n_7438)
);

NOR2xp33_ASAP7_75t_L g7439 ( 
.A(n_7391),
.B(n_7299),
.Y(n_7439)
);

OR2x2_ASAP7_75t_L g7440 ( 
.A(n_7337),
.B(n_7298),
.Y(n_7440)
);

OR2x2_ASAP7_75t_L g7441 ( 
.A(n_7337),
.B(n_7304),
.Y(n_7441)
);

INVx2_ASAP7_75t_SL g7442 ( 
.A(n_7347),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_7360),
.Y(n_7443)
);

AND2x2_ASAP7_75t_L g7444 ( 
.A(n_7396),
.B(n_7267),
.Y(n_7444)
);

NAND2xp5_ASAP7_75t_L g7445 ( 
.A(n_7351),
.B(n_7213),
.Y(n_7445)
);

AND2x2_ASAP7_75t_L g7446 ( 
.A(n_7332),
.B(n_7297),
.Y(n_7446)
);

INVx3_ASAP7_75t_L g7447 ( 
.A(n_7372),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_7338),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_7377),
.Y(n_7449)
);

NAND2xp5_ASAP7_75t_L g7450 ( 
.A(n_7401),
.B(n_7235),
.Y(n_7450)
);

INVx1_ASAP7_75t_L g7451 ( 
.A(n_7352),
.Y(n_7451)
);

INVx1_ASAP7_75t_L g7452 ( 
.A(n_7401),
.Y(n_7452)
);

INVx2_ASAP7_75t_L g7453 ( 
.A(n_7407),
.Y(n_7453)
);

AND2x2_ASAP7_75t_L g7454 ( 
.A(n_7341),
.B(n_7307),
.Y(n_7454)
);

INVx1_ASAP7_75t_L g7455 ( 
.A(n_7407),
.Y(n_7455)
);

OR2x2_ASAP7_75t_L g7456 ( 
.A(n_7358),
.B(n_7381),
.Y(n_7456)
);

OR2x2_ASAP7_75t_L g7457 ( 
.A(n_7381),
.B(n_7250),
.Y(n_7457)
);

OR2x2_ASAP7_75t_L g7458 ( 
.A(n_7353),
.B(n_7251),
.Y(n_7458)
);

AND2x2_ASAP7_75t_L g7459 ( 
.A(n_7354),
.B(n_7378),
.Y(n_7459)
);

AND2x2_ASAP7_75t_L g7460 ( 
.A(n_7393),
.B(n_7276),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_7415),
.Y(n_7461)
);

INVx1_ASAP7_75t_L g7462 ( 
.A(n_7415),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_7384),
.Y(n_7463)
);

INVx2_ASAP7_75t_L g7464 ( 
.A(n_7388),
.Y(n_7464)
);

AND2x2_ASAP7_75t_L g7465 ( 
.A(n_7344),
.B(n_7296),
.Y(n_7465)
);

INVx2_ASAP7_75t_L g7466 ( 
.A(n_7417),
.Y(n_7466)
);

AND2x2_ASAP7_75t_L g7467 ( 
.A(n_7342),
.B(n_7229),
.Y(n_7467)
);

BUFx2_ASAP7_75t_L g7468 ( 
.A(n_7368),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_7370),
.Y(n_7469)
);

NAND2xp5_ASAP7_75t_L g7470 ( 
.A(n_7356),
.B(n_7217),
.Y(n_7470)
);

NOR2x1p5_ASAP7_75t_L g7471 ( 
.A(n_7374),
.B(n_7322),
.Y(n_7471)
);

INVx1_ASAP7_75t_L g7472 ( 
.A(n_7416),
.Y(n_7472)
);

NAND2xp5_ASAP7_75t_L g7473 ( 
.A(n_7365),
.B(n_7226),
.Y(n_7473)
);

NAND2xp5_ASAP7_75t_L g7474 ( 
.A(n_7383),
.B(n_7227),
.Y(n_7474)
);

AND2x2_ASAP7_75t_L g7475 ( 
.A(n_7335),
.B(n_7302),
.Y(n_7475)
);

INVx1_ASAP7_75t_SL g7476 ( 
.A(n_7399),
.Y(n_7476)
);

OR2x2_ASAP7_75t_L g7477 ( 
.A(n_7376),
.B(n_7291),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7410),
.Y(n_7478)
);

INVx1_ASAP7_75t_L g7479 ( 
.A(n_7379),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_7371),
.Y(n_7480)
);

HB1xp67_ASAP7_75t_L g7481 ( 
.A(n_7371),
.Y(n_7481)
);

NAND2xp33_ASAP7_75t_L g7482 ( 
.A(n_7361),
.B(n_7291),
.Y(n_7482)
);

AND2x2_ASAP7_75t_L g7483 ( 
.A(n_7364),
.B(n_7331),
.Y(n_7483)
);

AND2x4_ASAP7_75t_L g7484 ( 
.A(n_7375),
.B(n_7310),
.Y(n_7484)
);

NAND4xp25_ASAP7_75t_L g7485 ( 
.A(n_7373),
.B(n_7282),
.C(n_7324),
.D(n_7293),
.Y(n_7485)
);

INVx1_ASAP7_75t_L g7486 ( 
.A(n_7366),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_L g7487 ( 
.A(n_7359),
.B(n_7275),
.Y(n_7487)
);

NAND2xp5_ASAP7_75t_L g7488 ( 
.A(n_7339),
.B(n_7270),
.Y(n_7488)
);

AND2x2_ASAP7_75t_L g7489 ( 
.A(n_7343),
.B(n_7278),
.Y(n_7489)
);

INVx1_ASAP7_75t_SL g7490 ( 
.A(n_7336),
.Y(n_7490)
);

AND2x2_ASAP7_75t_L g7491 ( 
.A(n_7339),
.B(n_7313),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_7369),
.Y(n_7492)
);

INVx1_ASAP7_75t_L g7493 ( 
.A(n_7411),
.Y(n_7493)
);

INVx2_ASAP7_75t_L g7494 ( 
.A(n_7382),
.Y(n_7494)
);

INVxp67_ASAP7_75t_SL g7495 ( 
.A(n_7334),
.Y(n_7495)
);

NAND3xp33_ASAP7_75t_SL g7496 ( 
.A(n_7349),
.B(n_7300),
.C(n_7293),
.Y(n_7496)
);

INVx2_ASAP7_75t_L g7497 ( 
.A(n_7423),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_7422),
.Y(n_7498)
);

AND2x2_ASAP7_75t_L g7499 ( 
.A(n_7430),
.B(n_7424),
.Y(n_7499)
);

OAI21xp5_ASAP7_75t_L g7500 ( 
.A1(n_7481),
.A2(n_7300),
.B(n_7394),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_7469),
.Y(n_7501)
);

INVx1_ASAP7_75t_L g7502 ( 
.A(n_7477),
.Y(n_7502)
);

INVx2_ASAP7_75t_L g7503 ( 
.A(n_7447),
.Y(n_7503)
);

OR2x2_ASAP7_75t_L g7504 ( 
.A(n_7490),
.B(n_7405),
.Y(n_7504)
);

AND2x2_ASAP7_75t_L g7505 ( 
.A(n_7430),
.B(n_7367),
.Y(n_7505)
);

NAND2xp5_ASAP7_75t_L g7506 ( 
.A(n_7490),
.B(n_7329),
.Y(n_7506)
);

NAND2xp5_ASAP7_75t_L g7507 ( 
.A(n_7447),
.B(n_7330),
.Y(n_7507)
);

NAND2xp5_ASAP7_75t_L g7508 ( 
.A(n_7495),
.B(n_7404),
.Y(n_7508)
);

AOI221xp5_ASAP7_75t_L g7509 ( 
.A1(n_7435),
.A2(n_7288),
.B1(n_7284),
.B2(n_7397),
.C(n_7398),
.Y(n_7509)
);

INVx2_ASAP7_75t_L g7510 ( 
.A(n_7428),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_7482),
.Y(n_7511)
);

AND2x2_ASAP7_75t_L g7512 ( 
.A(n_7446),
.B(n_7390),
.Y(n_7512)
);

INVxp33_ASAP7_75t_L g7513 ( 
.A(n_7465),
.Y(n_7513)
);

OAI22xp33_ASAP7_75t_L g7514 ( 
.A1(n_7426),
.A2(n_7288),
.B1(n_7284),
.B2(n_7400),
.Y(n_7514)
);

AND2x2_ASAP7_75t_L g7515 ( 
.A(n_7420),
.B(n_7389),
.Y(n_7515)
);

NOR2xp33_ASAP7_75t_L g7516 ( 
.A(n_7463),
.B(n_7408),
.Y(n_7516)
);

AOI21xp33_ASAP7_75t_SL g7517 ( 
.A1(n_7425),
.A2(n_7406),
.B(n_7403),
.Y(n_7517)
);

OR2x2_ASAP7_75t_L g7518 ( 
.A(n_7445),
.B(n_7419),
.Y(n_7518)
);

INVx2_ASAP7_75t_L g7519 ( 
.A(n_7458),
.Y(n_7519)
);

NAND2xp5_ASAP7_75t_L g7520 ( 
.A(n_7449),
.B(n_7412),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7457),
.Y(n_7521)
);

NAND2xp5_ASAP7_75t_L g7522 ( 
.A(n_7433),
.B(n_7385),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7467),
.Y(n_7523)
);

NAND2xp5_ASAP7_75t_L g7524 ( 
.A(n_7442),
.B(n_7392),
.Y(n_7524)
);

INVx1_ASAP7_75t_L g7525 ( 
.A(n_7460),
.Y(n_7525)
);

NAND2xp5_ASAP7_75t_L g7526 ( 
.A(n_7491),
.B(n_7402),
.Y(n_7526)
);

NOR2xp67_ASAP7_75t_L g7527 ( 
.A(n_7438),
.B(n_7414),
.Y(n_7527)
);

INVx2_ASAP7_75t_L g7528 ( 
.A(n_7453),
.Y(n_7528)
);

AND2x2_ASAP7_75t_L g7529 ( 
.A(n_7468),
.B(n_449),
.Y(n_7529)
);

INVx2_ASAP7_75t_L g7530 ( 
.A(n_7471),
.Y(n_7530)
);

NOR2x1_ASAP7_75t_L g7531 ( 
.A(n_7445),
.B(n_450),
.Y(n_7531)
);

AND2x2_ASAP7_75t_L g7532 ( 
.A(n_7489),
.B(n_450),
.Y(n_7532)
);

INVx1_ASAP7_75t_L g7533 ( 
.A(n_7450),
.Y(n_7533)
);

NAND2xp33_ASAP7_75t_SL g7534 ( 
.A(n_7456),
.B(n_451),
.Y(n_7534)
);

NAND2xp5_ASAP7_75t_L g7535 ( 
.A(n_7476),
.B(n_451),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7427),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7437),
.Y(n_7537)
);

OAI21xp33_ASAP7_75t_L g7538 ( 
.A1(n_7435),
.A2(n_452),
.B(n_453),
.Y(n_7538)
);

INVxp67_ASAP7_75t_SL g7539 ( 
.A(n_7439),
.Y(n_7539)
);

AND2x2_ASAP7_75t_L g7540 ( 
.A(n_7444),
.B(n_453),
.Y(n_7540)
);

NAND2xp5_ASAP7_75t_L g7541 ( 
.A(n_7476),
.B(n_454),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7452),
.Y(n_7542)
);

AND2x2_ASAP7_75t_L g7543 ( 
.A(n_7454),
.B(n_7459),
.Y(n_7543)
);

INVx2_ASAP7_75t_L g7544 ( 
.A(n_7455),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_7432),
.Y(n_7545)
);

INVx1_ASAP7_75t_L g7546 ( 
.A(n_7461),
.Y(n_7546)
);

OAI22xp5_ASAP7_75t_L g7547 ( 
.A1(n_7426),
.A2(n_7480),
.B1(n_7434),
.B2(n_7473),
.Y(n_7547)
);

INVx1_ASAP7_75t_L g7548 ( 
.A(n_7462),
.Y(n_7548)
);

INVx1_ASAP7_75t_L g7549 ( 
.A(n_7443),
.Y(n_7549)
);

INVx2_ASAP7_75t_SL g7550 ( 
.A(n_7484),
.Y(n_7550)
);

OR2x2_ASAP7_75t_L g7551 ( 
.A(n_7425),
.B(n_455),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7487),
.Y(n_7552)
);

NAND2xp5_ASAP7_75t_L g7553 ( 
.A(n_7421),
.B(n_455),
.Y(n_7553)
);

AO21x1_ASAP7_75t_SL g7554 ( 
.A1(n_7487),
.A2(n_456),
.B(n_458),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_L g7555 ( 
.A(n_7421),
.B(n_456),
.Y(n_7555)
);

OR2x2_ASAP7_75t_L g7556 ( 
.A(n_7473),
.B(n_459),
.Y(n_7556)
);

INVxp67_ASAP7_75t_L g7557 ( 
.A(n_7488),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_7440),
.Y(n_7558)
);

AND2x2_ASAP7_75t_L g7559 ( 
.A(n_7475),
.B(n_461),
.Y(n_7559)
);

AND2x2_ASAP7_75t_L g7560 ( 
.A(n_7431),
.B(n_461),
.Y(n_7560)
);

AND2x4_ASAP7_75t_L g7561 ( 
.A(n_7550),
.B(n_7484),
.Y(n_7561)
);

AOI22xp5_ASAP7_75t_L g7562 ( 
.A1(n_7557),
.A2(n_7485),
.B1(n_7496),
.B2(n_7448),
.Y(n_7562)
);

AOI22xp33_ASAP7_75t_L g7563 ( 
.A1(n_7531),
.A2(n_7485),
.B1(n_7493),
.B2(n_7466),
.Y(n_7563)
);

INVx2_ASAP7_75t_L g7564 ( 
.A(n_7499),
.Y(n_7564)
);

INVx1_ASAP7_75t_L g7565 ( 
.A(n_7505),
.Y(n_7565)
);

NOR2xp33_ASAP7_75t_L g7566 ( 
.A(n_7513),
.B(n_7464),
.Y(n_7566)
);

INVxp67_ASAP7_75t_L g7567 ( 
.A(n_7554),
.Y(n_7567)
);

NOR2x1p5_ASAP7_75t_L g7568 ( 
.A(n_7539),
.B(n_7494),
.Y(n_7568)
);

OAI22xp33_ASAP7_75t_L g7569 ( 
.A1(n_7504),
.A2(n_7488),
.B1(n_7441),
.B2(n_7470),
.Y(n_7569)
);

OAI22xp33_ASAP7_75t_L g7570 ( 
.A1(n_7522),
.A2(n_7470),
.B1(n_7478),
.B2(n_7472),
.Y(n_7570)
);

INVx1_ASAP7_75t_L g7571 ( 
.A(n_7553),
.Y(n_7571)
);

NAND2xp5_ASAP7_75t_L g7572 ( 
.A(n_7559),
.B(n_7421),
.Y(n_7572)
);

AND2x2_ASAP7_75t_L g7573 ( 
.A(n_7510),
.B(n_7515),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_7553),
.Y(n_7574)
);

OAI22xp5_ASAP7_75t_L g7575 ( 
.A1(n_7502),
.A2(n_7429),
.B1(n_7436),
.B2(n_7479),
.Y(n_7575)
);

OAI21xp5_ASAP7_75t_SL g7576 ( 
.A1(n_7511),
.A2(n_7483),
.B(n_7451),
.Y(n_7576)
);

NAND2xp5_ASAP7_75t_L g7577 ( 
.A(n_7532),
.B(n_7486),
.Y(n_7577)
);

INVx2_ASAP7_75t_L g7578 ( 
.A(n_7540),
.Y(n_7578)
);

OA21x2_ASAP7_75t_L g7579 ( 
.A1(n_7500),
.A2(n_7474),
.B(n_7492),
.Y(n_7579)
);

INVx2_ASAP7_75t_L g7580 ( 
.A(n_7530),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7555),
.Y(n_7581)
);

NAND2xp5_ASAP7_75t_L g7582 ( 
.A(n_7527),
.B(n_7474),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_7555),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_7508),
.Y(n_7584)
);

AND2x2_ASAP7_75t_L g7585 ( 
.A(n_7519),
.B(n_462),
.Y(n_7585)
);

INVx1_ASAP7_75t_SL g7586 ( 
.A(n_7508),
.Y(n_7586)
);

INVxp67_ASAP7_75t_L g7587 ( 
.A(n_7516),
.Y(n_7587)
);

AOI21xp5_ASAP7_75t_L g7588 ( 
.A1(n_7534),
.A2(n_462),
.B(n_464),
.Y(n_7588)
);

INVx1_ASAP7_75t_L g7589 ( 
.A(n_7551),
.Y(n_7589)
);

INVx1_ASAP7_75t_L g7590 ( 
.A(n_7503),
.Y(n_7590)
);

AND2x2_ASAP7_75t_L g7591 ( 
.A(n_7543),
.B(n_464),
.Y(n_7591)
);

NAND2xp5_ASAP7_75t_L g7592 ( 
.A(n_7523),
.B(n_465),
.Y(n_7592)
);

AOI221xp5_ASAP7_75t_L g7593 ( 
.A1(n_7547),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.C(n_472),
.Y(n_7593)
);

INVx2_ASAP7_75t_L g7594 ( 
.A(n_7512),
.Y(n_7594)
);

INVx1_ASAP7_75t_L g7595 ( 
.A(n_7529),
.Y(n_7595)
);

INVx2_ASAP7_75t_L g7596 ( 
.A(n_7556),
.Y(n_7596)
);

NOR2xp67_ASAP7_75t_L g7597 ( 
.A(n_7525),
.B(n_473),
.Y(n_7597)
);

AND2x2_ASAP7_75t_L g7598 ( 
.A(n_7497),
.B(n_474),
.Y(n_7598)
);

AND2x2_ASAP7_75t_L g7599 ( 
.A(n_7501),
.B(n_474),
.Y(n_7599)
);

INVx1_ASAP7_75t_L g7600 ( 
.A(n_7507),
.Y(n_7600)
);

AOI22xp5_ASAP7_75t_L g7601 ( 
.A1(n_7522),
.A2(n_478),
.B1(n_475),
.B2(n_476),
.Y(n_7601)
);

OAI22xp5_ASAP7_75t_L g7602 ( 
.A1(n_7506),
.A2(n_7545),
.B1(n_7552),
.B2(n_7521),
.Y(n_7602)
);

NAND2xp5_ASAP7_75t_L g7603 ( 
.A(n_7560),
.B(n_475),
.Y(n_7603)
);

AOI221xp5_ASAP7_75t_L g7604 ( 
.A1(n_7547),
.A2(n_7500),
.B1(n_7514),
.B2(n_7526),
.C(n_7558),
.Y(n_7604)
);

INVx1_ASAP7_75t_L g7605 ( 
.A(n_7507),
.Y(n_7605)
);

AOI22xp5_ASAP7_75t_L g7606 ( 
.A1(n_7526),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_7606)
);

INVx1_ASAP7_75t_L g7607 ( 
.A(n_7506),
.Y(n_7607)
);

INVx1_ASAP7_75t_SL g7608 ( 
.A(n_7524),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_7561),
.Y(n_7609)
);

AOI322xp5_ASAP7_75t_L g7610 ( 
.A1(n_7569),
.A2(n_7509),
.A3(n_7537),
.B1(n_7536),
.B2(n_7533),
.C1(n_7520),
.C2(n_7528),
.Y(n_7610)
);

XOR2x2_ASAP7_75t_L g7611 ( 
.A(n_7604),
.B(n_7524),
.Y(n_7611)
);

INVx1_ASAP7_75t_L g7612 ( 
.A(n_7561),
.Y(n_7612)
);

INVx1_ASAP7_75t_L g7613 ( 
.A(n_7573),
.Y(n_7613)
);

INVxp67_ASAP7_75t_L g7614 ( 
.A(n_7579),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_7579),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_7597),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_7597),
.Y(n_7617)
);

NAND2xp33_ASAP7_75t_SL g7618 ( 
.A(n_7568),
.B(n_7498),
.Y(n_7618)
);

OAI22xp5_ASAP7_75t_L g7619 ( 
.A1(n_7562),
.A2(n_7535),
.B1(n_7541),
.B2(n_7549),
.Y(n_7619)
);

AND2x2_ASAP7_75t_L g7620 ( 
.A(n_7564),
.B(n_7544),
.Y(n_7620)
);

INVx1_ASAP7_75t_L g7621 ( 
.A(n_7565),
.Y(n_7621)
);

AOI22xp5_ASAP7_75t_L g7622 ( 
.A1(n_7567),
.A2(n_7538),
.B1(n_7520),
.B2(n_7518),
.Y(n_7622)
);

INVx1_ASAP7_75t_L g7623 ( 
.A(n_7586),
.Y(n_7623)
);

NOR2xp67_ASAP7_75t_L g7624 ( 
.A(n_7607),
.B(n_7541),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7591),
.Y(n_7625)
);

AOI21xp33_ASAP7_75t_SL g7626 ( 
.A1(n_7602),
.A2(n_7570),
.B(n_7572),
.Y(n_7626)
);

INVx2_ASAP7_75t_L g7627 ( 
.A(n_7578),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7577),
.Y(n_7628)
);

AOI221xp5_ASAP7_75t_L g7629 ( 
.A1(n_7600),
.A2(n_7517),
.B1(n_7542),
.B2(n_7546),
.C(n_7548),
.Y(n_7629)
);

INVx1_ASAP7_75t_SL g7630 ( 
.A(n_7608),
.Y(n_7630)
);

OR2x2_ASAP7_75t_L g7631 ( 
.A(n_7594),
.B(n_479),
.Y(n_7631)
);

INVx1_ASAP7_75t_SL g7632 ( 
.A(n_7585),
.Y(n_7632)
);

AND2x2_ASAP7_75t_L g7633 ( 
.A(n_7590),
.B(n_481),
.Y(n_7633)
);

HB1xp67_ASAP7_75t_L g7634 ( 
.A(n_7584),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_7582),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7605),
.Y(n_7636)
);

NAND2xp5_ASAP7_75t_L g7637 ( 
.A(n_7588),
.B(n_482),
.Y(n_7637)
);

NAND2xp5_ASAP7_75t_L g7638 ( 
.A(n_7598),
.B(n_483),
.Y(n_7638)
);

NAND2xp5_ASAP7_75t_L g7639 ( 
.A(n_7562),
.B(n_483),
.Y(n_7639)
);

OAI21xp33_ASAP7_75t_L g7640 ( 
.A1(n_7630),
.A2(n_7566),
.B(n_7576),
.Y(n_7640)
);

INVx1_ASAP7_75t_L g7641 ( 
.A(n_7615),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_7634),
.Y(n_7642)
);

XOR2xp5_ASAP7_75t_L g7643 ( 
.A(n_7611),
.B(n_7595),
.Y(n_7643)
);

NAND2xp5_ASAP7_75t_L g7644 ( 
.A(n_7609),
.B(n_7563),
.Y(n_7644)
);

NAND2xp5_ASAP7_75t_SL g7645 ( 
.A(n_7626),
.B(n_7593),
.Y(n_7645)
);

INVxp67_ASAP7_75t_L g7646 ( 
.A(n_7612),
.Y(n_7646)
);

O2A1O1Ixp33_ASAP7_75t_SL g7647 ( 
.A1(n_7614),
.A2(n_7575),
.B(n_7587),
.C(n_7592),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_7613),
.Y(n_7648)
);

XOR2x2_ASAP7_75t_L g7649 ( 
.A(n_7622),
.B(n_7603),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7620),
.Y(n_7650)
);

XNOR2xp5_ASAP7_75t_L g7651 ( 
.A(n_7622),
.B(n_7632),
.Y(n_7651)
);

NAND2xp5_ASAP7_75t_L g7652 ( 
.A(n_7624),
.B(n_7625),
.Y(n_7652)
);

INVx1_ASAP7_75t_L g7653 ( 
.A(n_7616),
.Y(n_7653)
);

OAI22xp5_ASAP7_75t_L g7654 ( 
.A1(n_7623),
.A2(n_7580),
.B1(n_7601),
.B2(n_7574),
.Y(n_7654)
);

OAI211xp5_ASAP7_75t_L g7655 ( 
.A1(n_7610),
.A2(n_7581),
.B(n_7583),
.C(n_7571),
.Y(n_7655)
);

INVx1_ASAP7_75t_L g7656 ( 
.A(n_7617),
.Y(n_7656)
);

INVxp67_ASAP7_75t_L g7657 ( 
.A(n_7618),
.Y(n_7657)
);

XNOR2xp5_ASAP7_75t_L g7658 ( 
.A(n_7619),
.B(n_7596),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_7633),
.Y(n_7659)
);

INVx2_ASAP7_75t_L g7660 ( 
.A(n_7631),
.Y(n_7660)
);

INVx1_ASAP7_75t_SL g7661 ( 
.A(n_7638),
.Y(n_7661)
);

AOI21xp33_ASAP7_75t_SL g7662 ( 
.A1(n_7639),
.A2(n_7589),
.B(n_7599),
.Y(n_7662)
);

OAI21xp5_ASAP7_75t_L g7663 ( 
.A1(n_7610),
.A2(n_7601),
.B(n_7606),
.Y(n_7663)
);

OAI21xp33_ASAP7_75t_L g7664 ( 
.A1(n_7621),
.A2(n_7606),
.B(n_484),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_7627),
.Y(n_7665)
);

AOI21xp33_ASAP7_75t_L g7666 ( 
.A1(n_7636),
.A2(n_484),
.B(n_485),
.Y(n_7666)
);

NAND2xp5_ASAP7_75t_L g7667 ( 
.A(n_7628),
.B(n_485),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_7651),
.Y(n_7668)
);

INVx2_ASAP7_75t_L g7669 ( 
.A(n_7649),
.Y(n_7669)
);

AND2x2_ASAP7_75t_L g7670 ( 
.A(n_7650),
.B(n_7665),
.Y(n_7670)
);

INVx1_ASAP7_75t_L g7671 ( 
.A(n_7643),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_7658),
.Y(n_7672)
);

INVx2_ASAP7_75t_L g7673 ( 
.A(n_7660),
.Y(n_7673)
);

INVxp67_ASAP7_75t_L g7674 ( 
.A(n_7642),
.Y(n_7674)
);

INVx1_ASAP7_75t_SL g7675 ( 
.A(n_7644),
.Y(n_7675)
);

INVx8_ASAP7_75t_L g7676 ( 
.A(n_7646),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_7647),
.Y(n_7677)
);

INVx2_ASAP7_75t_L g7678 ( 
.A(n_7659),
.Y(n_7678)
);

INVxp67_ASAP7_75t_L g7679 ( 
.A(n_7652),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_7640),
.Y(n_7680)
);

INVx2_ASAP7_75t_L g7681 ( 
.A(n_7661),
.Y(n_7681)
);

INVx1_ASAP7_75t_L g7682 ( 
.A(n_7640),
.Y(n_7682)
);

INVx2_ASAP7_75t_L g7683 ( 
.A(n_7648),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_7663),
.Y(n_7684)
);

BUFx4f_ASAP7_75t_SL g7685 ( 
.A(n_7645),
.Y(n_7685)
);

INVx1_ASAP7_75t_L g7686 ( 
.A(n_7641),
.Y(n_7686)
);

INVx1_ASAP7_75t_L g7687 ( 
.A(n_7655),
.Y(n_7687)
);

NOR2xp33_ASAP7_75t_L g7688 ( 
.A(n_7662),
.B(n_7635),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_7667),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_7654),
.Y(n_7690)
);

INVxp67_ASAP7_75t_L g7691 ( 
.A(n_7653),
.Y(n_7691)
);

BUFx2_ASAP7_75t_L g7692 ( 
.A(n_7657),
.Y(n_7692)
);

INVx1_ASAP7_75t_L g7693 ( 
.A(n_7656),
.Y(n_7693)
);

INVx1_ASAP7_75t_L g7694 ( 
.A(n_7664),
.Y(n_7694)
);

INVx1_ASAP7_75t_L g7695 ( 
.A(n_7666),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_7651),
.Y(n_7696)
);

INVx1_ASAP7_75t_SL g7697 ( 
.A(n_7643),
.Y(n_7697)
);

INVx1_ASAP7_75t_SL g7698 ( 
.A(n_7643),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7651),
.Y(n_7699)
);

OAI21xp5_ASAP7_75t_SL g7700 ( 
.A1(n_7697),
.A2(n_7629),
.B(n_7637),
.Y(n_7700)
);

INVxp67_ASAP7_75t_L g7701 ( 
.A(n_7684),
.Y(n_7701)
);

AO22x2_ASAP7_75t_L g7702 ( 
.A1(n_7687),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_7702)
);

AOI22xp5_ASAP7_75t_L g7703 ( 
.A1(n_7697),
.A2(n_7698),
.B1(n_7683),
.B2(n_7676),
.Y(n_7703)
);

OAI21xp5_ASAP7_75t_L g7704 ( 
.A1(n_7698),
.A2(n_486),
.B(n_487),
.Y(n_7704)
);

BUFx6f_ASAP7_75t_L g7705 ( 
.A(n_7676),
.Y(n_7705)
);

AOI21xp5_ASAP7_75t_L g7706 ( 
.A1(n_7688),
.A2(n_489),
.B(n_490),
.Y(n_7706)
);

AOI221xp5_ASAP7_75t_L g7707 ( 
.A1(n_7676),
.A2(n_489),
.B1(n_492),
.B2(n_493),
.C(n_494),
.Y(n_7707)
);

AO22x1_ASAP7_75t_L g7708 ( 
.A1(n_7677),
.A2(n_494),
.B1(n_495),
.B2(n_497),
.Y(n_7708)
);

OAI221xp5_ASAP7_75t_L g7709 ( 
.A1(n_7692),
.A2(n_497),
.B1(n_498),
.B2(n_499),
.C(n_500),
.Y(n_7709)
);

NAND4xp25_ASAP7_75t_L g7710 ( 
.A(n_7675),
.B(n_498),
.C(n_500),
.D(n_501),
.Y(n_7710)
);

INVx1_ASAP7_75t_L g7711 ( 
.A(n_7675),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7685),
.Y(n_7712)
);

OAI211xp5_ASAP7_75t_SL g7713 ( 
.A1(n_7671),
.A2(n_504),
.B(n_505),
.C(n_507),
.Y(n_7713)
);

AOI22xp33_ASAP7_75t_L g7714 ( 
.A1(n_7689),
.A2(n_7686),
.B1(n_7673),
.B2(n_7695),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_7670),
.Y(n_7715)
);

A2O1A1Ixp33_ASAP7_75t_L g7716 ( 
.A1(n_7674),
.A2(n_507),
.B(n_508),
.C(n_509),
.Y(n_7716)
);

OAI221xp5_ASAP7_75t_L g7717 ( 
.A1(n_7691),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.C(n_511),
.Y(n_7717)
);

OAI211xp5_ASAP7_75t_L g7718 ( 
.A1(n_7680),
.A2(n_510),
.B(n_511),
.C(n_512),
.Y(n_7718)
);

AOI211xp5_ASAP7_75t_SL g7719 ( 
.A1(n_7679),
.A2(n_512),
.B(n_513),
.C(n_514),
.Y(n_7719)
);

AOI21xp5_ASAP7_75t_SL g7720 ( 
.A1(n_7682),
.A2(n_513),
.B(n_514),
.Y(n_7720)
);

OAI22xp33_ASAP7_75t_L g7721 ( 
.A1(n_7693),
.A2(n_7681),
.B1(n_7678),
.B2(n_7699),
.Y(n_7721)
);

HB1xp67_ASAP7_75t_L g7722 ( 
.A(n_7690),
.Y(n_7722)
);

OAI21xp5_ASAP7_75t_SL g7723 ( 
.A1(n_7668),
.A2(n_515),
.B(n_516),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7669),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_L g7725 ( 
.A(n_7696),
.B(n_516),
.Y(n_7725)
);

AOI221xp5_ASAP7_75t_L g7726 ( 
.A1(n_7672),
.A2(n_518),
.B1(n_519),
.B2(n_521),
.C(n_523),
.Y(n_7726)
);

OAI22xp5_ASAP7_75t_L g7727 ( 
.A1(n_7694),
.A2(n_518),
.B1(n_519),
.B2(n_521),
.Y(n_7727)
);

OAI22xp5_ASAP7_75t_L g7728 ( 
.A1(n_7691),
.A2(n_525),
.B1(n_526),
.B2(n_527),
.Y(n_7728)
);

NOR3xp33_ASAP7_75t_L g7729 ( 
.A(n_7697),
.B(n_526),
.C(n_527),
.Y(n_7729)
);

INVxp67_ASAP7_75t_L g7730 ( 
.A(n_7684),
.Y(n_7730)
);

AOI22xp5_ASAP7_75t_L g7731 ( 
.A1(n_7697),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_7731)
);

AOI22xp5_ASAP7_75t_L g7732 ( 
.A1(n_7703),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.Y(n_7732)
);

NAND4xp25_ASAP7_75t_L g7733 ( 
.A(n_7714),
.B(n_532),
.C(n_533),
.D(n_534),
.Y(n_7733)
);

AOI221xp5_ASAP7_75t_SL g7734 ( 
.A1(n_7721),
.A2(n_532),
.B1(n_535),
.B2(n_537),
.C(n_538),
.Y(n_7734)
);

NAND2xp33_ASAP7_75t_R g7735 ( 
.A(n_7711),
.B(n_535),
.Y(n_7735)
);

NOR2x1_ASAP7_75t_L g7736 ( 
.A(n_7715),
.B(n_537),
.Y(n_7736)
);

AOI222xp33_ASAP7_75t_L g7737 ( 
.A1(n_7701),
.A2(n_7730),
.B1(n_7705),
.B2(n_7722),
.C1(n_7724),
.C2(n_7700),
.Y(n_7737)
);

AOI221xp5_ASAP7_75t_L g7738 ( 
.A1(n_7705),
.A2(n_539),
.B1(n_540),
.B2(n_541),
.C(n_542),
.Y(n_7738)
);

NOR2xp33_ASAP7_75t_L g7739 ( 
.A(n_7705),
.B(n_539),
.Y(n_7739)
);

OAI21xp33_ASAP7_75t_SL g7740 ( 
.A1(n_7712),
.A2(n_540),
.B(n_541),
.Y(n_7740)
);

OAI211xp5_ASAP7_75t_L g7741 ( 
.A1(n_7723),
.A2(n_544),
.B(n_545),
.C(n_547),
.Y(n_7741)
);

O2A1O1Ixp33_ASAP7_75t_L g7742 ( 
.A1(n_7725),
.A2(n_544),
.B(n_545),
.C(n_549),
.Y(n_7742)
);

AOI22xp5_ASAP7_75t_L g7743 ( 
.A1(n_7729),
.A2(n_7710),
.B1(n_7702),
.B2(n_7713),
.Y(n_7743)
);

OAI22xp5_ASAP7_75t_L g7744 ( 
.A1(n_7731),
.A2(n_550),
.B1(n_551),
.B2(n_552),
.Y(n_7744)
);

AOI322xp5_ASAP7_75t_L g7745 ( 
.A1(n_7726),
.A2(n_550),
.A3(n_551),
.B1(n_552),
.B2(n_553),
.C1(n_555),
.C2(n_556),
.Y(n_7745)
);

INVx1_ASAP7_75t_SL g7746 ( 
.A(n_7708),
.Y(n_7746)
);

AOI211xp5_ASAP7_75t_L g7747 ( 
.A1(n_7720),
.A2(n_556),
.B(n_557),
.C(n_558),
.Y(n_7747)
);

AOI21xp5_ASAP7_75t_L g7748 ( 
.A1(n_7702),
.A2(n_557),
.B(n_559),
.Y(n_7748)
);

OAI21xp33_ASAP7_75t_L g7749 ( 
.A1(n_7704),
.A2(n_560),
.B(n_561),
.Y(n_7749)
);

NAND3xp33_ASAP7_75t_L g7750 ( 
.A(n_7719),
.B(n_560),
.C(n_562),
.Y(n_7750)
);

AOI211xp5_ASAP7_75t_L g7751 ( 
.A1(n_7718),
.A2(n_564),
.B(n_565),
.C(n_567),
.Y(n_7751)
);

OAI211xp5_ASAP7_75t_L g7752 ( 
.A1(n_7706),
.A2(n_564),
.B(n_568),
.C(n_569),
.Y(n_7752)
);

A2O1A1Ixp33_ASAP7_75t_L g7753 ( 
.A1(n_7716),
.A2(n_568),
.B(n_570),
.C(n_571),
.Y(n_7753)
);

AOI221xp5_ASAP7_75t_L g7754 ( 
.A1(n_7728),
.A2(n_571),
.B1(n_573),
.B2(n_574),
.C(n_575),
.Y(n_7754)
);

OAI211xp5_ASAP7_75t_L g7755 ( 
.A1(n_7707),
.A2(n_574),
.B(n_575),
.C(n_576),
.Y(n_7755)
);

AOI22xp5_ASAP7_75t_L g7756 ( 
.A1(n_7727),
.A2(n_576),
.B1(n_577),
.B2(n_578),
.Y(n_7756)
);

NAND2xp5_ASAP7_75t_L g7757 ( 
.A(n_7709),
.B(n_578),
.Y(n_7757)
);

NAND4xp25_ASAP7_75t_L g7758 ( 
.A(n_7717),
.B(n_579),
.C(n_580),
.D(n_581),
.Y(n_7758)
);

AOI211xp5_ASAP7_75t_L g7759 ( 
.A1(n_7721),
.A2(n_579),
.B(n_580),
.C(n_582),
.Y(n_7759)
);

A2O1A1Ixp33_ASAP7_75t_L g7760 ( 
.A1(n_7703),
.A2(n_583),
.B(n_584),
.C(n_585),
.Y(n_7760)
);

AOI21xp33_ASAP7_75t_L g7761 ( 
.A1(n_7737),
.A2(n_583),
.B(n_584),
.Y(n_7761)
);

NOR4xp25_ASAP7_75t_L g7762 ( 
.A(n_7746),
.B(n_586),
.C(n_587),
.D(n_588),
.Y(n_7762)
);

AOI221xp5_ASAP7_75t_L g7763 ( 
.A1(n_7740),
.A2(n_589),
.B1(n_590),
.B2(n_591),
.C(n_593),
.Y(n_7763)
);

NAND2xp5_ASAP7_75t_L g7764 ( 
.A(n_7736),
.B(n_589),
.Y(n_7764)
);

O2A1O1Ixp33_ASAP7_75t_L g7765 ( 
.A1(n_7760),
.A2(n_593),
.B(n_594),
.C(n_595),
.Y(n_7765)
);

NOR2x1_ASAP7_75t_SL g7766 ( 
.A(n_7741),
.B(n_594),
.Y(n_7766)
);

AOI221xp5_ASAP7_75t_L g7767 ( 
.A1(n_7750),
.A2(n_596),
.B1(n_597),
.B2(n_598),
.C(n_599),
.Y(n_7767)
);

AOI22xp5_ASAP7_75t_L g7768 ( 
.A1(n_7735),
.A2(n_596),
.B1(n_597),
.B2(n_598),
.Y(n_7768)
);

OAI21xp33_ASAP7_75t_L g7769 ( 
.A1(n_7749),
.A2(n_600),
.B(n_601),
.Y(n_7769)
);

AOI21xp5_ASAP7_75t_L g7770 ( 
.A1(n_7757),
.A2(n_600),
.B(n_601),
.Y(n_7770)
);

AOI22xp5_ASAP7_75t_L g7771 ( 
.A1(n_7743),
.A2(n_7744),
.B1(n_7758),
.B2(n_7733),
.Y(n_7771)
);

AOI211xp5_ASAP7_75t_L g7772 ( 
.A1(n_7755),
.A2(n_602),
.B(n_603),
.C(n_604),
.Y(n_7772)
);

OAI211xp5_ASAP7_75t_SL g7773 ( 
.A1(n_7747),
.A2(n_602),
.B(n_603),
.C(n_605),
.Y(n_7773)
);

AND2x2_ASAP7_75t_L g7774 ( 
.A(n_7734),
.B(n_7751),
.Y(n_7774)
);

INVx1_ASAP7_75t_SL g7775 ( 
.A(n_7748),
.Y(n_7775)
);

NAND3xp33_ASAP7_75t_SL g7776 ( 
.A(n_7759),
.B(n_606),
.C(n_607),
.Y(n_7776)
);

OAI21xp5_ASAP7_75t_SL g7777 ( 
.A1(n_7742),
.A2(n_608),
.B(n_609),
.Y(n_7777)
);

O2A1O1Ixp33_ASAP7_75t_L g7778 ( 
.A1(n_7753),
.A2(n_7739),
.B(n_7752),
.C(n_7754),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7732),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_7766),
.Y(n_7780)
);

INVx1_ASAP7_75t_L g7781 ( 
.A(n_7764),
.Y(n_7781)
);

AOI22xp5_ASAP7_75t_L g7782 ( 
.A1(n_7774),
.A2(n_7756),
.B1(n_7738),
.B2(n_7745),
.Y(n_7782)
);

INVx1_ASAP7_75t_L g7783 ( 
.A(n_7768),
.Y(n_7783)
);

INVx1_ASAP7_75t_L g7784 ( 
.A(n_7775),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_7773),
.Y(n_7785)
);

NOR2x1_ASAP7_75t_L g7786 ( 
.A(n_7776),
.B(n_609),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_7771),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7765),
.Y(n_7788)
);

INVx3_ASAP7_75t_L g7789 ( 
.A(n_7779),
.Y(n_7789)
);

INVx1_ASAP7_75t_L g7790 ( 
.A(n_7777),
.Y(n_7790)
);

INVxp67_ASAP7_75t_SL g7791 ( 
.A(n_7761),
.Y(n_7791)
);

INVx1_ASAP7_75t_L g7792 ( 
.A(n_7778),
.Y(n_7792)
);

INVx2_ASAP7_75t_L g7793 ( 
.A(n_7762),
.Y(n_7793)
);

INVx2_ASAP7_75t_L g7794 ( 
.A(n_7772),
.Y(n_7794)
);

INVx1_ASAP7_75t_L g7795 ( 
.A(n_7769),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_7770),
.Y(n_7796)
);

NOR3xp33_ASAP7_75t_L g7797 ( 
.A(n_7784),
.B(n_7763),
.C(n_7767),
.Y(n_7797)
);

INVxp67_ASAP7_75t_L g7798 ( 
.A(n_7780),
.Y(n_7798)
);

INVx1_ASAP7_75t_L g7799 ( 
.A(n_7789),
.Y(n_7799)
);

INVxp67_ASAP7_75t_L g7800 ( 
.A(n_7789),
.Y(n_7800)
);

OAI22xp5_ASAP7_75t_SL g7801 ( 
.A1(n_7793),
.A2(n_610),
.B1(n_611),
.B2(n_612),
.Y(n_7801)
);

INVx2_ASAP7_75t_L g7802 ( 
.A(n_7786),
.Y(n_7802)
);

NAND2xp5_ASAP7_75t_L g7803 ( 
.A(n_7792),
.B(n_610),
.Y(n_7803)
);

XNOR2xp5_ASAP7_75t_L g7804 ( 
.A(n_7787),
.B(n_612),
.Y(n_7804)
);

NOR3xp33_ASAP7_75t_L g7805 ( 
.A(n_7781),
.B(n_614),
.C(n_616),
.Y(n_7805)
);

NAND2xp5_ASAP7_75t_L g7806 ( 
.A(n_7796),
.B(n_614),
.Y(n_7806)
);

NAND4xp75_ASAP7_75t_L g7807 ( 
.A(n_7790),
.B(n_618),
.C(n_619),
.D(n_620),
.Y(n_7807)
);

O2A1O1Ixp33_ASAP7_75t_L g7808 ( 
.A1(n_7791),
.A2(n_621),
.B(n_624),
.C(n_625),
.Y(n_7808)
);

OR2x2_ASAP7_75t_L g7809 ( 
.A(n_7785),
.B(n_621),
.Y(n_7809)
);

AND2x4_ASAP7_75t_L g7810 ( 
.A(n_7783),
.B(n_624),
.Y(n_7810)
);

XNOR2x1_ASAP7_75t_L g7811 ( 
.A(n_7782),
.B(n_625),
.Y(n_7811)
);

NAND3xp33_ASAP7_75t_L g7812 ( 
.A(n_7788),
.B(n_626),
.C(n_627),
.Y(n_7812)
);

NAND4xp75_ASAP7_75t_L g7813 ( 
.A(n_7795),
.B(n_626),
.C(n_627),
.D(n_628),
.Y(n_7813)
);

CKINVDCx6p67_ASAP7_75t_R g7814 ( 
.A(n_7794),
.Y(n_7814)
);

AOI221xp5_ASAP7_75t_L g7815 ( 
.A1(n_7792),
.A2(n_628),
.B1(n_629),
.B2(n_631),
.C(n_632),
.Y(n_7815)
);

NAND2xp33_ASAP7_75t_L g7816 ( 
.A(n_7805),
.B(n_629),
.Y(n_7816)
);

NOR2xp33_ASAP7_75t_R g7817 ( 
.A(n_7814),
.B(n_632),
.Y(n_7817)
);

NOR2xp33_ASAP7_75t_R g7818 ( 
.A(n_7799),
.B(n_635),
.Y(n_7818)
);

NAND2xp33_ASAP7_75t_SL g7819 ( 
.A(n_7801),
.B(n_635),
.Y(n_7819)
);

NAND3xp33_ASAP7_75t_L g7820 ( 
.A(n_7800),
.B(n_1330),
.C(n_1328),
.Y(n_7820)
);

NOR2xp33_ASAP7_75t_R g7821 ( 
.A(n_7804),
.B(n_636),
.Y(n_7821)
);

NOR2xp33_ASAP7_75t_R g7822 ( 
.A(n_7803),
.B(n_637),
.Y(n_7822)
);

NAND2xp5_ASAP7_75t_SL g7823 ( 
.A(n_7798),
.B(n_638),
.Y(n_7823)
);

NAND3xp33_ASAP7_75t_L g7824 ( 
.A(n_7802),
.B(n_1330),
.C(n_1328),
.Y(n_7824)
);

NOR2xp33_ASAP7_75t_R g7825 ( 
.A(n_7806),
.B(n_638),
.Y(n_7825)
);

NOR2xp33_ASAP7_75t_R g7826 ( 
.A(n_7809),
.B(n_639),
.Y(n_7826)
);

NOR2xp33_ASAP7_75t_R g7827 ( 
.A(n_7810),
.B(n_639),
.Y(n_7827)
);

NOR2xp33_ASAP7_75t_R g7828 ( 
.A(n_7810),
.B(n_640),
.Y(n_7828)
);

NAND2xp5_ASAP7_75t_SL g7829 ( 
.A(n_7815),
.B(n_641),
.Y(n_7829)
);

NOR2xp33_ASAP7_75t_R g7830 ( 
.A(n_7811),
.B(n_642),
.Y(n_7830)
);

NAND2xp5_ASAP7_75t_L g7831 ( 
.A(n_7797),
.B(n_642),
.Y(n_7831)
);

XNOR2xp5_ASAP7_75t_L g7832 ( 
.A(n_7807),
.B(n_643),
.Y(n_7832)
);

NOR2xp33_ASAP7_75t_R g7833 ( 
.A(n_7813),
.B(n_643),
.Y(n_7833)
);

OR4x1_ASAP7_75t_L g7834 ( 
.A(n_7831),
.B(n_7808),
.C(n_7812),
.D(n_646),
.Y(n_7834)
);

NAND4xp25_ASAP7_75t_L g7835 ( 
.A(n_7819),
.B(n_644),
.C(n_645),
.D(n_647),
.Y(n_7835)
);

INVx2_ASAP7_75t_L g7836 ( 
.A(n_7832),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_7827),
.Y(n_7837)
);

NAND5xp2_ASAP7_75t_L g7838 ( 
.A(n_7830),
.B(n_644),
.C(n_645),
.D(n_647),
.E(n_648),
.Y(n_7838)
);

NAND3xp33_ASAP7_75t_SL g7839 ( 
.A(n_7817),
.B(n_650),
.C(n_651),
.Y(n_7839)
);

NOR3xp33_ASAP7_75t_SL g7840 ( 
.A(n_7820),
.B(n_651),
.C(n_652),
.Y(n_7840)
);

AND5x1_ASAP7_75t_L g7841 ( 
.A(n_7833),
.B(n_654),
.C(n_655),
.D(n_656),
.E(n_657),
.Y(n_7841)
);

OR4x2_ASAP7_75t_L g7842 ( 
.A(n_7821),
.B(n_655),
.C(n_656),
.D(n_657),
.Y(n_7842)
);

HB1xp67_ASAP7_75t_L g7843 ( 
.A(n_7828),
.Y(n_7843)
);

OAI22x1_ASAP7_75t_L g7844 ( 
.A1(n_7823),
.A2(n_658),
.B1(n_660),
.B2(n_661),
.Y(n_7844)
);

AND2x4_ASAP7_75t_L g7845 ( 
.A(n_7829),
.B(n_7824),
.Y(n_7845)
);

INVx2_ASAP7_75t_SL g7846 ( 
.A(n_7843),
.Y(n_7846)
);

CKINVDCx5p33_ASAP7_75t_R g7847 ( 
.A(n_7837),
.Y(n_7847)
);

INVx2_ASAP7_75t_L g7848 ( 
.A(n_7842),
.Y(n_7848)
);

NAND2xp5_ASAP7_75t_L g7849 ( 
.A(n_7836),
.B(n_7826),
.Y(n_7849)
);

BUFx6f_ASAP7_75t_L g7850 ( 
.A(n_7845),
.Y(n_7850)
);

NOR2xp33_ASAP7_75t_L g7851 ( 
.A(n_7838),
.B(n_7816),
.Y(n_7851)
);

NAND3x1_ASAP7_75t_L g7852 ( 
.A(n_7841),
.B(n_7818),
.C(n_7825),
.Y(n_7852)
);

INVx1_ASAP7_75t_L g7853 ( 
.A(n_7852),
.Y(n_7853)
);

XNOR2xp5_ASAP7_75t_L g7854 ( 
.A(n_7846),
.B(n_7839),
.Y(n_7854)
);

NAND2xp33_ASAP7_75t_SL g7855 ( 
.A(n_7848),
.B(n_7822),
.Y(n_7855)
);

AOI22xp33_ASAP7_75t_L g7856 ( 
.A1(n_7850),
.A2(n_7835),
.B1(n_7844),
.B2(n_7834),
.Y(n_7856)
);

AOI22xp5_ASAP7_75t_L g7857 ( 
.A1(n_7853),
.A2(n_7855),
.B1(n_7850),
.B2(n_7851),
.Y(n_7857)
);

AND2x4_ASAP7_75t_L g7858 ( 
.A(n_7856),
.B(n_7849),
.Y(n_7858)
);

AOI22xp5_ASAP7_75t_L g7859 ( 
.A1(n_7854),
.A2(n_7847),
.B1(n_7840),
.B2(n_663),
.Y(n_7859)
);

XNOR2xp5_ASAP7_75t_L g7860 ( 
.A(n_7857),
.B(n_658),
.Y(n_7860)
);

AOI22xp33_ASAP7_75t_L g7861 ( 
.A1(n_7860),
.A2(n_7858),
.B1(n_7859),
.B2(n_664),
.Y(n_7861)
);

OAI22xp5_ASAP7_75t_SL g7862 ( 
.A1(n_7861),
.A2(n_662),
.B1(n_663),
.B2(n_665),
.Y(n_7862)
);

AOI22xp33_ASAP7_75t_L g7863 ( 
.A1(n_7862),
.A2(n_666),
.B1(n_667),
.B2(n_668),
.Y(n_7863)
);

XNOR2xp5_ASAP7_75t_L g7864 ( 
.A(n_7863),
.B(n_667),
.Y(n_7864)
);

INVx1_ASAP7_75t_L g7865 ( 
.A(n_7864),
.Y(n_7865)
);

AOI22xp33_ASAP7_75t_SL g7866 ( 
.A1(n_7865),
.A2(n_668),
.B1(n_670),
.B2(n_671),
.Y(n_7866)
);

OAI221xp5_ASAP7_75t_R g7867 ( 
.A1(n_7866),
.A2(n_671),
.B1(n_672),
.B2(n_673),
.C(n_674),
.Y(n_7867)
);

AOI21xp33_ASAP7_75t_L g7868 ( 
.A1(n_7867),
.A2(n_673),
.B(n_675),
.Y(n_7868)
);

AOI211xp5_ASAP7_75t_L g7869 ( 
.A1(n_7868),
.A2(n_677),
.B(n_678),
.C(n_679),
.Y(n_7869)
);


endmodule