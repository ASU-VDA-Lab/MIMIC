module fake_jpeg_169_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_10),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_72),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_55),
.B1(n_53),
.B2(n_42),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_45),
.B1(n_43),
.B2(n_47),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_52),
.B1(n_44),
.B2(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_54),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_1),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_71),
.Y(n_88)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_85),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_102),
.C(n_9),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_3),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_51),
.B1(n_42),
.B2(n_52),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_76),
.C(n_84),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_16),
.C(n_38),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_23),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_18),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_2),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_116),
.B1(n_11),
.B2(n_13),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_105),
.B(n_100),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_119),
.B(n_112),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_7),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_120),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_9),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_11),
.C(n_12),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_120),
.C(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_129),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_26),
.B1(n_35),
.B2(n_30),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_131),
.B1(n_24),
.B2(n_25),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_10),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_130),
.C(n_28),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_133),
.B(n_127),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_139),
.B(n_144),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_125),
.C(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_146),
.B(n_149),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_132),
.B1(n_131),
.B2(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_146),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_150),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_148),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_151),
.B(n_140),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_27),
.Y(n_158)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_158),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_29),
.Y(n_160)
);


endmodule