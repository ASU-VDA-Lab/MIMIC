module fake_aes_8385_n_10 (n_3, n_1, n_2, n_0, n_10);
input n_3;
input n_1;
input n_2;
input n_0;
output n_10;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_7;
wire n_8;
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_1), .B(n_3), .Y(n_4) );
AO21x1_ASAP7_75t_L g5 ( .A1(n_2), .A2(n_1), .B(n_0), .Y(n_5) );
OR2x2_ASAP7_75t_L g6 ( .A(n_5), .B(n_0), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_4), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_7), .B(n_6), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
endmodule