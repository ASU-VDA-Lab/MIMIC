module fake_netlist_6_1830_n_5264 (n_992, n_1, n_801, n_1234, n_1458, n_1199, n_741, n_1027, n_1351, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_212, n_700, n_50, n_1307, n_1038, n_578, n_1581, n_1003, n_365, n_168, n_1237, n_1061, n_1357, n_77, n_783, n_798, n_188, n_1575, n_509, n_1342, n_245, n_1209, n_1348, n_1387, n_677, n_805, n_1151, n_396, n_350, n_78, n_1380, n_442, n_480, n_142, n_1402, n_1009, n_62, n_1160, n_883, n_1238, n_1032, n_1247, n_1547, n_1553, n_893, n_1099, n_1264, n_1192, n_471, n_424, n_1555, n_1415, n_1370, n_369, n_287, n_415, n_830, n_65, n_230, n_461, n_873, n_141, n_383, n_1285, n_1371, n_200, n_447, n_1172, n_852, n_71, n_229, n_1532, n_1393, n_1517, n_1078, n_250, n_544, n_1140, n_1444, n_1579, n_35, n_1263, n_836, n_375, n_522, n_1261, n_945, n_1511, n_1143, n_1422, n_1232, n_1572, n_616, n_658, n_1119, n_428, n_1433, n_1541, n_1300, n_641, n_822, n_693, n_1313, n_1056, n_758, n_516, n_1455, n_1163, n_1180, n_943, n_1550, n_491, n_42, n_772, n_1344, n_666, n_371, n_940, n_770, n_567, n_405, n_213, n_538, n_1106, n_886, n_1471, n_343, n_953, n_1094, n_1345, n_494, n_539, n_493, n_155, n_45, n_454, n_1421, n_638, n_1404, n_1211, n_381, n_887, n_112, n_1280, n_713, n_1400, n_126, n_1467, n_58, n_976, n_224, n_48, n_1445, n_1526, n_1560, n_734, n_1088, n_196, n_1231, n_917, n_574, n_9, n_907, n_6, n_1446, n_14, n_659, n_407, n_913, n_808, n_867, n_1230, n_473, n_1193, n_1054, n_559, n_1333, n_44, n_163, n_1558, n_281, n_551, n_699, n_564, n_451, n_824, n_279, n_686, n_757, n_594, n_577, n_166, n_619, n_1367, n_1336, n_521, n_572, n_395, n_813, n_1481, n_323, n_606, n_1441, n_818, n_1123, n_1309, n_92, n_513, n_645, n_1381, n_331, n_916, n_483, n_102, n_608, n_261, n_630, n_32, n_541, n_512, n_121, n_433, n_792, n_476, n_2, n_1328, n_219, n_264, n_263, n_1162, n_860, n_1530, n_788, n_939, n_1543, n_821, n_938, n_1302, n_1068, n_329, n_982, n_549, n_1075, n_408, n_932, n_61, n_237, n_243, n_979, n_905, n_117, n_175, n_322, n_993, n_689, n_354, n_1330, n_1413, n_134, n_1278, n_547, n_558, n_1064, n_1396, n_634, n_136, n_966, n_764, n_692, n_733, n_1233, n_1289, n_487, n_241, n_30, n_1107, n_1014, n_1290, n_882, n_1354, n_586, n_423, n_318, n_1111, n_715, n_1251, n_1265, n_88, n_530, n_1563, n_277, n_618, n_1297, n_1312, n_199, n_1167, n_1359, n_674, n_871, n_922, n_268, n_1335, n_210, n_1069, n_5, n_612, n_178, n_247, n_1165, n_355, n_702, n_347, n_1175, n_328, n_1386, n_429, n_1012, n_195, n_780, n_675, n_903, n_1540, n_1504, n_286, n_254, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_816, n_1157, n_1462, n_1188, n_877, n_604, n_825, n_728, n_1063, n_26, n_55, n_267, n_1124, n_515, n_598, n_696, n_1515, n_961, n_437, n_1082, n_1317, n_593, n_514, n_687, n_697, n_890, n_637, n_295, n_701, n_950, n_388, n_190, n_484, n_170, n_891, n_1412, n_949, n_678, n_283, n_91, n_507, n_968, n_909, n_1369, n_881, n_1008, n_760, n_1546, n_590, n_63, n_362, n_148, n_161, n_22, n_462, n_1033, n_1052, n_1296, n_304, n_694, n_1294, n_1420, n_125, n_297, n_595, n_627, n_524, n_1465, n_342, n_1044, n_1391, n_449, n_131, n_1523, n_1208, n_1164, n_1295, n_1072, n_1527, n_1495, n_1438, n_495, n_815, n_1100, n_585, n_1487, n_840, n_874, n_1128, n_382, n_673, n_1071, n_1067, n_1565, n_1493, n_898, n_255, n_284, n_865, n_925, n_1101, n_15, n_1026, n_38, n_289, n_1364, n_615, n_1249, n_59, n_1293, n_1127, n_1512, n_1451, n_320, n_108, n_639, n_963, n_794, n_727, n_894, n_685, n_353, n_605, n_1514, n_826, n_872, n_1139, n_86, n_104, n_718, n_1018, n_1521, n_1366, n_542, n_847, n_644, n_682, n_851, n_305, n_72, n_996, n_532, n_173, n_1308, n_1376, n_1513, n_413, n_791, n_510, n_837, n_79, n_1488, n_948, n_704, n_977, n_1005, n_536, n_622, n_147, n_1469, n_581, n_765, n_432, n_987, n_1492, n_1340, n_631, n_720, n_153, n_842, n_1432, n_156, n_145, n_843, n_656, n_989, n_1277, n_797, n_1473, n_1246, n_899, n_189, n_738, n_1304, n_1035, n_294, n_499, n_1426, n_705, n_11, n_1004, n_1176, n_1529, n_1022, n_614, n_529, n_425, n_684, n_1431, n_1474, n_1571, n_1577, n_1181, n_37, n_486, n_947, n_1117, n_1087, n_1448, n_648, n_657, n_1049, n_1505, n_803, n_290, n_118, n_926, n_927, n_919, n_478, n_929, n_107, n_1228, n_417, n_446, n_89, n_1568, n_1490, n_777, n_1299, n_272, n_526, n_1183, n_1436, n_1384, n_69, n_293, n_53, n_458, n_1070, n_998, n_16, n_717, n_18, n_154, n_1383, n_1178, n_98, n_1424, n_1073, n_1000, n_796, n_252, n_1195, n_1507, n_184, n_552, n_1358, n_1388, n_216, n_912, n_1519, n_745, n_1284, n_1142, n_716, n_1475, n_623, n_1048, n_1201, n_1398, n_884, n_1395, n_731, n_1502, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_312, n_1368, n_66, n_1418, n_958, n_292, n_1250, n_100, n_1137, n_880, n_889, n_150, n_1478, n_589, n_1310, n_819, n_1363, n_1334, n_767, n_1314, n_600, n_964, n_831, n_477, n_954, n_864, n_1110, n_1410, n_399, n_1440, n_124, n_1382, n_1534, n_1564, n_211, n_1483, n_1372, n_231, n_40, n_1457, n_505, n_319, n_1339, n_537, n_1427, n_311, n_1466, n_10, n_403, n_1080, n_723, n_596, n_123, n_546, n_562, n_1141, n_1268, n_386, n_1220, n_556, n_162, n_1136, n_128, n_1125, n_970, n_642, n_995, n_276, n_1159, n_1092, n_441, n_221, n_1060, n_444, n_146, n_1252, n_1223, n_303, n_511, n_193, n_1286, n_1053, n_416, n_520, n_418, n_1093, n_113, n_1533, n_4, n_266, n_296, n_775, n_651, n_1153, n_439, n_217, n_518, n_1531, n_1185, n_453, n_215, n_914, n_759, n_426, n_317, n_90, n_54, n_1453, n_488, n_497, n_773, n_920, n_99, n_1374, n_1315, n_13, n_1224, n_1459, n_1135, n_1169, n_1179, n_401, n_324, n_335, n_1470, n_463, n_1243, n_848, n_120, n_301, n_274, n_1096, n_1091, n_1580, n_1425, n_36, n_1267, n_1281, n_983, n_427, n_1520, n_496, n_906, n_1390, n_688, n_1077, n_1419, n_351, n_259, n_177, n_1437, n_385, n_1439, n_1323, n_858, n_1331, n_613, n_736, n_501, n_956, n_960, n_663, n_856, n_379, n_778, n_1134, n_410, n_1129, n_554, n_602, n_664, n_171, n_169, n_1429, n_435, n_793, n_326, n_587, n_580, n_762, n_1030, n_1202, n_465, n_1079, n_341, n_828, n_607, n_316, n_419, n_28, n_1551, n_1103, n_144, n_1203, n_820, n_951, n_106, n_725, n_952, n_999, n_358, n_1254, n_160, n_186, n_0, n_368, n_575, n_994, n_1508, n_732, n_974, n_392, n_724, n_1020, n_1042, n_628, n_1273, n_1434, n_1573, n_557, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_1275, n_485, n_1549, n_67, n_443, n_1510, n_892, n_768, n_421, n_1468, n_238, n_1095, n_202, n_597, n_280, n_1270, n_1187, n_610, n_1403, n_1024, n_198, n_179, n_248, n_517, n_667, n_1206, n_621, n_1037, n_1397, n_1279, n_1115, n_750, n_901, n_1499, n_468, n_923, n_504, n_1409, n_183, n_1015, n_1503, n_466, n_1057, n_603, n_991, n_235, n_1126, n_340, n_710, n_1108, n_1182, n_1298, n_39, n_73, n_785, n_746, n_609, n_101, n_167, n_1356, n_127, n_1497, n_1168, n_1216, n_133, n_1320, n_96, n_1430, n_1316, n_1287, n_1452, n_1586, n_302, n_380, n_1535, n_137, n_20, n_1190, n_397, n_122, n_34, n_1262, n_218, n_1213, n_70, n_1350, n_172, n_1443, n_1272, n_239, n_97, n_782, n_1539, n_490, n_220, n_809, n_1043, n_986, n_80, n_1472, n_1081, n_402, n_352, n_800, n_1084, n_1171, n_460, n_1361, n_1491, n_662, n_374, n_1152, n_450, n_921, n_1346, n_711, n_579, n_1352, n_937, n_370, n_650, n_1046, n_1145, n_330, n_1121, n_1102, n_972, n_1405, n_258, n_1406, n_456, n_1332, n_260, n_313, n_624, n_962, n_1041, n_565, n_356, n_1569, n_936, n_1288, n_1186, n_1062, n_885, n_896, n_83, n_654, n_411, n_152, n_1222, n_599, n_776, n_321, n_105, n_227, n_204, n_482, n_934, n_1407, n_420, n_1341, n_394, n_1456, n_1489, n_164, n_23, n_942, n_1524, n_543, n_1496, n_1271, n_1545, n_1355, n_1225, n_1544, n_1485, n_325, n_804, n_464, n_533, n_806, n_879, n_959, n_584, n_244, n_1343, n_1522, n_76, n_548, n_94, n_282, n_833, n_1567, n_523, n_1319, n_707, n_345, n_799, n_1548, n_1155, n_139, n_41, n_273, n_787, n_1416, n_1528, n_1146, n_159, n_1086, n_1066, n_157, n_1282, n_550, n_275, n_652, n_560, n_1484, n_1241, n_1321, n_569, n_737, n_1318, n_1235, n_1229, n_306, n_1292, n_1373, n_21, n_346, n_3, n_1029, n_1447, n_790, n_138, n_1498, n_1210, n_49, n_299, n_1248, n_1556, n_902, n_333, n_1047, n_1385, n_431, n_24, n_459, n_1269, n_502, n_672, n_1257, n_285, n_1375, n_85, n_655, n_706, n_1045, n_786, n_1236, n_1559, n_834, n_19, n_29, n_75, n_743, n_766, n_430, n_1325, n_1002, n_545, n_489, n_251, n_1019, n_636, n_729, n_110, n_151, n_876, n_774, n_1337, n_660, n_438, n_1477, n_1360, n_1200, n_479, n_1353, n_1454, n_869, n_1154, n_1113, n_646, n_528, n_391, n_1098, n_1329, n_817, n_262, n_187, n_897, n_846, n_841, n_1476, n_1001, n_508, n_1050, n_1411, n_1463, n_1177, n_332, n_1150, n_1562, n_398, n_1191, n_566, n_1023, n_1076, n_1118, n_194, n_57, n_1007, n_1378, n_855, n_52, n_591, n_1377, n_256, n_853, n_440, n_695, n_1542, n_875, n_209, n_367, n_680, n_661, n_278, n_1256, n_671, n_7, n_933, n_740, n_703, n_978, n_384, n_1291, n_1217, n_751, n_749, n_310, n_1324, n_1399, n_1435, n_969, n_988, n_1065, n_84, n_1401, n_1255, n_568, n_1516, n_143, n_1536, n_180, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_1394, n_1327, n_1326, n_739, n_400, n_955, n_337, n_1379, n_214, n_246, n_1338, n_1097, n_935, n_781, n_789, n_1554, n_1130, n_181, n_182, n_573, n_769, n_676, n_327, n_1120, n_832, n_1583, n_555, n_389, n_814, n_669, n_176, n_114, n_300, n_222, n_747, n_74, n_1389, n_1105, n_721, n_1461, n_742, n_535, n_691, n_372, n_111, n_314, n_1408, n_378, n_1196, n_377, n_863, n_601, n_338, n_1283, n_918, n_748, n_506, n_1114, n_56, n_763, n_1147, n_360, n_1506, n_119, n_957, n_895, n_866, n_1227, n_191, n_387, n_452, n_744, n_971, n_946, n_344, n_761, n_1303, n_1205, n_1258, n_1392, n_174, n_1173, n_525, n_1116, n_611, n_1570, n_1219, n_8, n_1174, n_1016, n_1347, n_795, n_1501, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_1083, n_109, n_445, n_1561, n_930, n_888, n_1112, n_234, n_910, n_1460, n_911, n_82, n_1464, n_27, n_236, n_653, n_1414, n_752, n_908, n_944, n_576, n_1028, n_472, n_270, n_414, n_563, n_1011, n_1566, n_1215, n_25, n_93, n_839, n_708, n_668, n_626, n_990, n_1500, n_779, n_1537, n_1104, n_854, n_1058, n_498, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_1509, n_103, n_1109, n_185, n_712, n_348, n_1276, n_376, n_390, n_1148, n_31, n_334, n_1161, n_1085, n_232, n_46, n_1239, n_771, n_1584, n_470, n_475, n_924, n_298, n_1582, n_492, n_1149, n_265, n_1184, n_228, n_719, n_1525, n_455, n_1585, n_363, n_1090, n_592, n_1518, n_829, n_1156, n_1362, n_393, n_984, n_503, n_1450, n_132, n_868, n_570, n_859, n_406, n_735, n_878, n_620, n_130, n_519, n_307, n_469, n_1218, n_500, n_1482, n_981, n_714, n_1349, n_291, n_1144, n_357, n_985, n_481, n_997, n_1301, n_802, n_561, n_33, n_980, n_1306, n_1198, n_436, n_116, n_409, n_1244, n_1574, n_240, n_756, n_810, n_1133, n_635, n_95, n_1194, n_1051, n_253, n_1552, n_583, n_249, n_201, n_1039, n_1442, n_1034, n_1480, n_1158, n_754, n_941, n_975, n_1031, n_115, n_1305, n_553, n_43, n_849, n_753, n_467, n_269, n_359, n_973, n_1479, n_1055, n_582, n_861, n_857, n_967, n_571, n_271, n_404, n_158, n_206, n_679, n_633, n_1170, n_665, n_588, n_225, n_1260, n_308, n_309, n_1010, n_149, n_1040, n_915, n_632, n_1166, n_812, n_1131, n_534, n_1578, n_1006, n_373, n_87, n_257, n_1557, n_730, n_1311, n_1494, n_670, n_203, n_207, n_1089, n_1365, n_1417, n_205, n_1242, n_681, n_1226, n_1274, n_1486, n_412, n_640, n_1322, n_81, n_965, n_1428, n_1576, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_422, n_722, n_862, n_135, n_165, n_540, n_1423, n_457, n_364, n_629, n_900, n_1449, n_531, n_827, n_60, n_361, n_1025, n_336, n_12, n_1013, n_1259, n_192, n_1538, n_51, n_649, n_1240, n_5264);

input n_992;
input n_1;
input n_801;
input n_1234;
input n_1458;
input n_1199;
input n_741;
input n_1027;
input n_1351;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_212;
input n_700;
input n_50;
input n_1307;
input n_1038;
input n_578;
input n_1581;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_1357;
input n_77;
input n_783;
input n_798;
input n_188;
input n_1575;
input n_509;
input n_1342;
input n_245;
input n_1209;
input n_1348;
input n_1387;
input n_677;
input n_805;
input n_1151;
input n_396;
input n_350;
input n_78;
input n_1380;
input n_442;
input n_480;
input n_142;
input n_1402;
input n_1009;
input n_62;
input n_1160;
input n_883;
input n_1238;
input n_1032;
input n_1247;
input n_1547;
input n_1553;
input n_893;
input n_1099;
input n_1264;
input n_1192;
input n_471;
input n_424;
input n_1555;
input n_1415;
input n_1370;
input n_369;
input n_287;
input n_415;
input n_830;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_1371;
input n_200;
input n_447;
input n_1172;
input n_852;
input n_71;
input n_229;
input n_1532;
input n_1393;
input n_1517;
input n_1078;
input n_250;
input n_544;
input n_1140;
input n_1444;
input n_1579;
input n_35;
input n_1263;
input n_836;
input n_375;
input n_522;
input n_1261;
input n_945;
input n_1511;
input n_1143;
input n_1422;
input n_1232;
input n_1572;
input n_616;
input n_658;
input n_1119;
input n_428;
input n_1433;
input n_1541;
input n_1300;
input n_641;
input n_822;
input n_693;
input n_1313;
input n_1056;
input n_758;
input n_516;
input n_1455;
input n_1163;
input n_1180;
input n_943;
input n_1550;
input n_491;
input n_42;
input n_772;
input n_1344;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_405;
input n_213;
input n_538;
input n_1106;
input n_886;
input n_1471;
input n_343;
input n_953;
input n_1094;
input n_1345;
input n_494;
input n_539;
input n_493;
input n_155;
input n_45;
input n_454;
input n_1421;
input n_638;
input n_1404;
input n_1211;
input n_381;
input n_887;
input n_112;
input n_1280;
input n_713;
input n_1400;
input n_126;
input n_1467;
input n_58;
input n_976;
input n_224;
input n_48;
input n_1445;
input n_1526;
input n_1560;
input n_734;
input n_1088;
input n_196;
input n_1231;
input n_917;
input n_574;
input n_9;
input n_907;
input n_6;
input n_1446;
input n_14;
input n_659;
input n_407;
input n_913;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1054;
input n_559;
input n_1333;
input n_44;
input n_163;
input n_1558;
input n_281;
input n_551;
input n_699;
input n_564;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_577;
input n_166;
input n_619;
input n_1367;
input n_1336;
input n_521;
input n_572;
input n_395;
input n_813;
input n_1481;
input n_323;
input n_606;
input n_1441;
input n_818;
input n_1123;
input n_1309;
input n_92;
input n_513;
input n_645;
input n_1381;
input n_331;
input n_916;
input n_483;
input n_102;
input n_608;
input n_261;
input n_630;
input n_32;
input n_541;
input n_512;
input n_121;
input n_433;
input n_792;
input n_476;
input n_2;
input n_1328;
input n_219;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_1530;
input n_788;
input n_939;
input n_1543;
input n_821;
input n_938;
input n_1302;
input n_1068;
input n_329;
input n_982;
input n_549;
input n_1075;
input n_408;
input n_932;
input n_61;
input n_237;
input n_243;
input n_979;
input n_905;
input n_117;
input n_175;
input n_322;
input n_993;
input n_689;
input n_354;
input n_1330;
input n_1413;
input n_134;
input n_1278;
input n_547;
input n_558;
input n_1064;
input n_1396;
input n_634;
input n_136;
input n_966;
input n_764;
input n_692;
input n_733;
input n_1233;
input n_1289;
input n_487;
input n_241;
input n_30;
input n_1107;
input n_1014;
input n_1290;
input n_882;
input n_1354;
input n_586;
input n_423;
input n_318;
input n_1111;
input n_715;
input n_1251;
input n_1265;
input n_88;
input n_530;
input n_1563;
input n_277;
input n_618;
input n_1297;
input n_1312;
input n_199;
input n_1167;
input n_1359;
input n_674;
input n_871;
input n_922;
input n_268;
input n_1335;
input n_210;
input n_1069;
input n_5;
input n_612;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_1175;
input n_328;
input n_1386;
input n_429;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_903;
input n_1540;
input n_1504;
input n_286;
input n_254;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_816;
input n_1157;
input n_1462;
input n_1188;
input n_877;
input n_604;
input n_825;
input n_728;
input n_1063;
input n_26;
input n_55;
input n_267;
input n_1124;
input n_515;
input n_598;
input n_696;
input n_1515;
input n_961;
input n_437;
input n_1082;
input n_1317;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_295;
input n_701;
input n_950;
input n_388;
input n_190;
input n_484;
input n_170;
input n_891;
input n_1412;
input n_949;
input n_678;
input n_283;
input n_91;
input n_507;
input n_968;
input n_909;
input n_1369;
input n_881;
input n_1008;
input n_760;
input n_1546;
input n_590;
input n_63;
input n_362;
input n_148;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_1296;
input n_304;
input n_694;
input n_1294;
input n_1420;
input n_125;
input n_297;
input n_595;
input n_627;
input n_524;
input n_1465;
input n_342;
input n_1044;
input n_1391;
input n_449;
input n_131;
input n_1523;
input n_1208;
input n_1164;
input n_1295;
input n_1072;
input n_1527;
input n_1495;
input n_1438;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_1487;
input n_840;
input n_874;
input n_1128;
input n_382;
input n_673;
input n_1071;
input n_1067;
input n_1565;
input n_1493;
input n_898;
input n_255;
input n_284;
input n_865;
input n_925;
input n_1101;
input n_15;
input n_1026;
input n_38;
input n_289;
input n_1364;
input n_615;
input n_1249;
input n_59;
input n_1293;
input n_1127;
input n_1512;
input n_1451;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_605;
input n_1514;
input n_826;
input n_872;
input n_1139;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_1521;
input n_1366;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_305;
input n_72;
input n_996;
input n_532;
input n_173;
input n_1308;
input n_1376;
input n_1513;
input n_413;
input n_791;
input n_510;
input n_837;
input n_79;
input n_1488;
input n_948;
input n_704;
input n_977;
input n_1005;
input n_536;
input n_622;
input n_147;
input n_1469;
input n_581;
input n_765;
input n_432;
input n_987;
input n_1492;
input n_1340;
input n_631;
input n_720;
input n_153;
input n_842;
input n_1432;
input n_156;
input n_145;
input n_843;
input n_656;
input n_989;
input n_1277;
input n_797;
input n_1473;
input n_1246;
input n_899;
input n_189;
input n_738;
input n_1304;
input n_1035;
input n_294;
input n_499;
input n_1426;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_1529;
input n_1022;
input n_614;
input n_529;
input n_425;
input n_684;
input n_1431;
input n_1474;
input n_1571;
input n_1577;
input n_1181;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_1087;
input n_1448;
input n_648;
input n_657;
input n_1049;
input n_1505;
input n_803;
input n_290;
input n_118;
input n_926;
input n_927;
input n_919;
input n_478;
input n_929;
input n_107;
input n_1228;
input n_417;
input n_446;
input n_89;
input n_1568;
input n_1490;
input n_777;
input n_1299;
input n_272;
input n_526;
input n_1183;
input n_1436;
input n_1384;
input n_69;
input n_293;
input n_53;
input n_458;
input n_1070;
input n_998;
input n_16;
input n_717;
input n_18;
input n_154;
input n_1383;
input n_1178;
input n_98;
input n_1424;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_1507;
input n_184;
input n_552;
input n_1358;
input n_1388;
input n_216;
input n_912;
input n_1519;
input n_745;
input n_1284;
input n_1142;
input n_716;
input n_1475;
input n_623;
input n_1048;
input n_1201;
input n_1398;
input n_884;
input n_1395;
input n_731;
input n_1502;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_312;
input n_1368;
input n_66;
input n_1418;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_880;
input n_889;
input n_150;
input n_1478;
input n_589;
input n_1310;
input n_819;
input n_1363;
input n_1334;
input n_767;
input n_1314;
input n_600;
input n_964;
input n_831;
input n_477;
input n_954;
input n_864;
input n_1110;
input n_1410;
input n_399;
input n_1440;
input n_124;
input n_1382;
input n_1534;
input n_1564;
input n_211;
input n_1483;
input n_1372;
input n_231;
input n_40;
input n_1457;
input n_505;
input n_319;
input n_1339;
input n_537;
input n_1427;
input n_311;
input n_1466;
input n_10;
input n_403;
input n_1080;
input n_723;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1220;
input n_556;
input n_162;
input n_1136;
input n_128;
input n_1125;
input n_970;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_1092;
input n_441;
input n_221;
input n_1060;
input n_444;
input n_146;
input n_1252;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1286;
input n_1053;
input n_416;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_1533;
input n_4;
input n_266;
input n_296;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_217;
input n_518;
input n_1531;
input n_1185;
input n_453;
input n_215;
input n_914;
input n_759;
input n_426;
input n_317;
input n_90;
input n_54;
input n_1453;
input n_488;
input n_497;
input n_773;
input n_920;
input n_99;
input n_1374;
input n_1315;
input n_13;
input n_1224;
input n_1459;
input n_1135;
input n_1169;
input n_1179;
input n_401;
input n_324;
input n_335;
input n_1470;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_301;
input n_274;
input n_1096;
input n_1091;
input n_1580;
input n_1425;
input n_36;
input n_1267;
input n_1281;
input n_983;
input n_427;
input n_1520;
input n_496;
input n_906;
input n_1390;
input n_688;
input n_1077;
input n_1419;
input n_351;
input n_259;
input n_177;
input n_1437;
input n_385;
input n_1439;
input n_1323;
input n_858;
input n_1331;
input n_613;
input n_736;
input n_501;
input n_956;
input n_960;
input n_663;
input n_856;
input n_379;
input n_778;
input n_1134;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_664;
input n_171;
input n_169;
input n_1429;
input n_435;
input n_793;
input n_326;
input n_587;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_465;
input n_1079;
input n_341;
input n_828;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1551;
input n_1103;
input n_144;
input n_1203;
input n_820;
input n_951;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_1508;
input n_732;
input n_974;
input n_392;
input n_724;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_1434;
input n_1573;
input n_557;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_1275;
input n_485;
input n_1549;
input n_67;
input n_443;
input n_1510;
input n_892;
input n_768;
input n_421;
input n_1468;
input n_238;
input n_1095;
input n_202;
input n_597;
input n_280;
input n_1270;
input n_1187;
input n_610;
input n_1403;
input n_1024;
input n_198;
input n_179;
input n_248;
input n_517;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1397;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_1499;
input n_468;
input n_923;
input n_504;
input n_1409;
input n_183;
input n_1015;
input n_1503;
input n_466;
input n_1057;
input n_603;
input n_991;
input n_235;
input n_1126;
input n_340;
input n_710;
input n_1108;
input n_1182;
input n_1298;
input n_39;
input n_73;
input n_785;
input n_746;
input n_609;
input n_101;
input n_167;
input n_1356;
input n_127;
input n_1497;
input n_1168;
input n_1216;
input n_133;
input n_1320;
input n_96;
input n_1430;
input n_1316;
input n_1287;
input n_1452;
input n_1586;
input n_302;
input n_380;
input n_1535;
input n_137;
input n_20;
input n_1190;
input n_397;
input n_122;
input n_34;
input n_1262;
input n_218;
input n_1213;
input n_70;
input n_1350;
input n_172;
input n_1443;
input n_1272;
input n_239;
input n_97;
input n_782;
input n_1539;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_986;
input n_80;
input n_1472;
input n_1081;
input n_402;
input n_352;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_1361;
input n_1491;
input n_662;
input n_374;
input n_1152;
input n_450;
input n_921;
input n_1346;
input n_711;
input n_579;
input n_1352;
input n_937;
input n_370;
input n_650;
input n_1046;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_972;
input n_1405;
input n_258;
input n_1406;
input n_456;
input n_1332;
input n_260;
input n_313;
input n_624;
input n_962;
input n_1041;
input n_565;
input n_356;
input n_1569;
input n_936;
input n_1288;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_654;
input n_411;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_105;
input n_227;
input n_204;
input n_482;
input n_934;
input n_1407;
input n_420;
input n_1341;
input n_394;
input n_1456;
input n_1489;
input n_164;
input n_23;
input n_942;
input n_1524;
input n_543;
input n_1496;
input n_1271;
input n_1545;
input n_1355;
input n_1225;
input n_1544;
input n_1485;
input n_325;
input n_804;
input n_464;
input n_533;
input n_806;
input n_879;
input n_959;
input n_584;
input n_244;
input n_1343;
input n_1522;
input n_76;
input n_548;
input n_94;
input n_282;
input n_833;
input n_1567;
input n_523;
input n_1319;
input n_707;
input n_345;
input n_799;
input n_1548;
input n_1155;
input n_139;
input n_41;
input n_273;
input n_787;
input n_1416;
input n_1528;
input n_1146;
input n_159;
input n_1086;
input n_1066;
input n_157;
input n_1282;
input n_550;
input n_275;
input n_652;
input n_560;
input n_1484;
input n_1241;
input n_1321;
input n_569;
input n_737;
input n_1318;
input n_1235;
input n_1229;
input n_306;
input n_1292;
input n_1373;
input n_21;
input n_346;
input n_3;
input n_1029;
input n_1447;
input n_790;
input n_138;
input n_1498;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_1556;
input n_902;
input n_333;
input n_1047;
input n_1385;
input n_431;
input n_24;
input n_459;
input n_1269;
input n_502;
input n_672;
input n_1257;
input n_285;
input n_1375;
input n_85;
input n_655;
input n_706;
input n_1045;
input n_786;
input n_1236;
input n_1559;
input n_834;
input n_19;
input n_29;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1325;
input n_1002;
input n_545;
input n_489;
input n_251;
input n_1019;
input n_636;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_1337;
input n_660;
input n_438;
input n_1477;
input n_1360;
input n_1200;
input n_479;
input n_1353;
input n_1454;
input n_869;
input n_1154;
input n_1113;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_1329;
input n_817;
input n_262;
input n_187;
input n_897;
input n_846;
input n_841;
input n_1476;
input n_1001;
input n_508;
input n_1050;
input n_1411;
input n_1463;
input n_1177;
input n_332;
input n_1150;
input n_1562;
input n_398;
input n_1191;
input n_566;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_1378;
input n_855;
input n_52;
input n_591;
input n_1377;
input n_256;
input n_853;
input n_440;
input n_695;
input n_1542;
input n_875;
input n_209;
input n_367;
input n_680;
input n_661;
input n_278;
input n_1256;
input n_671;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_384;
input n_1291;
input n_1217;
input n_751;
input n_749;
input n_310;
input n_1324;
input n_1399;
input n_1435;
input n_969;
input n_988;
input n_1065;
input n_84;
input n_1401;
input n_1255;
input n_568;
input n_1516;
input n_143;
input n_1536;
input n_180;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_1394;
input n_1327;
input n_1326;
input n_739;
input n_400;
input n_955;
input n_337;
input n_1379;
input n_214;
input n_246;
input n_1338;
input n_1097;
input n_935;
input n_781;
input n_789;
input n_1554;
input n_1130;
input n_181;
input n_182;
input n_573;
input n_769;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_1583;
input n_555;
input n_389;
input n_814;
input n_669;
input n_176;
input n_114;
input n_300;
input n_222;
input n_747;
input n_74;
input n_1389;
input n_1105;
input n_721;
input n_1461;
input n_742;
input n_535;
input n_691;
input n_372;
input n_111;
input n_314;
input n_1408;
input n_378;
input n_1196;
input n_377;
input n_863;
input n_601;
input n_338;
input n_1283;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1147;
input n_360;
input n_1506;
input n_119;
input n_957;
input n_895;
input n_866;
input n_1227;
input n_191;
input n_387;
input n_452;
input n_744;
input n_971;
input n_946;
input n_344;
input n_761;
input n_1303;
input n_1205;
input n_1258;
input n_1392;
input n_174;
input n_1173;
input n_525;
input n_1116;
input n_611;
input n_1570;
input n_1219;
input n_8;
input n_1174;
input n_1016;
input n_1347;
input n_795;
input n_1501;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_1083;
input n_109;
input n_445;
input n_1561;
input n_930;
input n_888;
input n_1112;
input n_234;
input n_910;
input n_1460;
input n_911;
input n_82;
input n_1464;
input n_27;
input n_236;
input n_653;
input n_1414;
input n_752;
input n_908;
input n_944;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_414;
input n_563;
input n_1011;
input n_1566;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_708;
input n_668;
input n_626;
input n_990;
input n_1500;
input n_779;
input n_1537;
input n_1104;
input n_854;
input n_1058;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_1509;
input n_103;
input n_1109;
input n_185;
input n_712;
input n_348;
input n_1276;
input n_376;
input n_390;
input n_1148;
input n_31;
input n_334;
input n_1161;
input n_1085;
input n_232;
input n_46;
input n_1239;
input n_771;
input n_1584;
input n_470;
input n_475;
input n_924;
input n_298;
input n_1582;
input n_492;
input n_1149;
input n_265;
input n_1184;
input n_228;
input n_719;
input n_1525;
input n_455;
input n_1585;
input n_363;
input n_1090;
input n_592;
input n_1518;
input n_829;
input n_1156;
input n_1362;
input n_393;
input n_984;
input n_503;
input n_1450;
input n_132;
input n_868;
input n_570;
input n_859;
input n_406;
input n_735;
input n_878;
input n_620;
input n_130;
input n_519;
input n_307;
input n_469;
input n_1218;
input n_500;
input n_1482;
input n_981;
input n_714;
input n_1349;
input n_291;
input n_1144;
input n_357;
input n_985;
input n_481;
input n_997;
input n_1301;
input n_802;
input n_561;
input n_33;
input n_980;
input n_1306;
input n_1198;
input n_436;
input n_116;
input n_409;
input n_1244;
input n_1574;
input n_240;
input n_756;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_1051;
input n_253;
input n_1552;
input n_583;
input n_249;
input n_201;
input n_1039;
input n_1442;
input n_1034;
input n_1480;
input n_1158;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_1305;
input n_553;
input n_43;
input n_849;
input n_753;
input n_467;
input n_269;
input n_359;
input n_973;
input n_1479;
input n_1055;
input n_582;
input n_861;
input n_857;
input n_967;
input n_571;
input n_271;
input n_404;
input n_158;
input n_206;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1010;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_812;
input n_1131;
input n_534;
input n_1578;
input n_1006;
input n_373;
input n_87;
input n_257;
input n_1557;
input n_730;
input n_1311;
input n_1494;
input n_670;
input n_203;
input n_207;
input n_1089;
input n_1365;
input n_1417;
input n_205;
input n_1242;
input n_681;
input n_1226;
input n_1274;
input n_1486;
input n_412;
input n_640;
input n_1322;
input n_81;
input n_965;
input n_1428;
input n_1576;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_422;
input n_722;
input n_862;
input n_135;
input n_165;
input n_540;
input n_1423;
input n_457;
input n_364;
input n_629;
input n_900;
input n_1449;
input n_531;
input n_827;
input n_60;
input n_361;
input n_1025;
input n_336;
input n_12;
input n_1013;
input n_1259;
input n_192;
input n_1538;
input n_51;
input n_649;
input n_1240;

output n_5264;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5254;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_3089;
wire n_4978;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_4829;
wire n_3222;
wire n_4699;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_3376;
wire n_4868;
wire n_3801;
wire n_4249;
wire n_3564;
wire n_1844;
wire n_5057;
wire n_3030;
wire n_2838;
wire n_5229;
wire n_3427;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_2786;
wire n_5239;
wire n_1971;
wire n_1781;
wire n_2004;
wire n_4814;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_3664;
wire n_1936;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_4262;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_5063;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_2764;
wire n_2895;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_4993;
wire n_2072;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_2514;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_4394;
wire n_2279;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_3696;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_3614;
wire n_5183;
wire n_2145;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_3179;
wire n_3400;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_2239;
wire n_4310;
wire n_5212;
wire n_2689;
wire n_2191;
wire n_4528;
wire n_4914;
wire n_4939;
wire n_3418;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_3631;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_4551;
wire n_2857;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_5035;
wire n_3390;
wire n_3656;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_3006;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_4592;
wire n_2199;
wire n_2661;
wire n_1955;
wire n_1791;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_3606;
wire n_3591;
wire n_2788;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_5176;
wire n_4428;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_2822;
wire n_4180;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_4761;
wire n_2884;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_4189;
wire n_3817;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_4380;
wire n_4996;
wire n_4990;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_3594;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_4601;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_2798;
wire n_2852;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_3375;
wire n_3899;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_4512;
wire n_4081;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_5124;
wire n_3951;
wire n_3569;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_3027;
wire n_4083;
wire n_1810;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_4027;
wire n_3154;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_4095;
wire n_2881;
wire n_1702;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_3697;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_3478;
wire n_3936;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_3101;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_3552;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_3444;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_3017;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_3795;
wire n_3852;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_3266;
wire n_3574;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_4504;
wire n_3844;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_5248;
wire n_1708;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_3275;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_2356;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_3750;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_2058;
wire n_2660;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_4047;
wire n_3413;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_4277;
wire n_4526;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_3725;
wire n_3933;
wire n_2311;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_4146;
wire n_1802;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_2271;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_2954;
wire n_2728;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_3159;
wire n_4701;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_3922;
wire n_5204;
wire n_4991;
wire n_2554;
wire n_1913;
wire n_4934;
wire n_5087;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_2604;
wire n_2407;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_2948;
wire n_2119;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_3837;
wire n_2718;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_3324;
wire n_2338;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_2144;
wire n_1604;
wire n_4487;
wire n_4866;
wire n_4889;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2892;
wire n_2132;
wire n_4120;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1951;
wire n_4362;
wire n_3311;
wire n_3913;
wire n_5121;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_4404;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_4132;
wire n_2995;
wire n_4844;
wire n_4438;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_3250;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_3414;
wire n_4870;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_2598;
wire n_1916;
wire n_1683;
wire n_4304;
wire n_4558;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_4016;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_3730;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2808;
wire n_2037;
wire n_4567;
wire n_5150;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_2970;
wire n_2342;
wire n_2167;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_2258;
wire n_2390;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_2734;
wire n_1782;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_3381;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_4143;
wire n_4170;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_2588;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_5170;
wire n_2827;
wire n_3515;
wire n_2951;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_4543;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_3629;
wire n_3920;
wire n_4892;
wire n_3255;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_4783;
wire n_4910;
wire n_3083;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5203;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_2430;
wire n_2721;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_4521;
wire n_3204;
wire n_4920;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_2726;
wire n_4303;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_1856;
wire n_2077;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_3111;
wire n_1885;
wire n_3054;
wire n_4730;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_3619;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1867;
wire n_2630;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_2256;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_2806;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_3624;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_2378;
wire n_2655;
wire n_4600;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_2593;
wire n_4255;
wire n_4071;
wire n_3568;
wire n_3850;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_2961;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_4745;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_3599;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_3022;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_4800;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_2691;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5168;
wire n_4661;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_3053;
wire n_1808;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_5125;
wire n_2650;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_4097;
wire n_1666;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_3590;
wire n_2435;
wire n_4419;
wire n_5184;
wire n_1736;
wire n_4053;
wire n_3848;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_2745;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5079;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_2783;
wire n_3188;
wire n_2462;
wire n_3243;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_5049;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_4754;
wire n_2993;
wire n_4647;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_4983;
wire n_1778;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_3636;
wire n_2327;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_3637;
wire n_4574;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_3236;
wire n_2755;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_2722;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1692;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_2789;
wire n_5152;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_3134;
wire n_3115;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_4145;
wire n_4901;
wire n_4821;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_2141;
wire n_3930;
wire n_4943;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_2021;
wire n_4942;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_5186;
wire n_2417;
wire n_5093;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1872;
wire n_5040;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_2045;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_2565;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_2566;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_4106;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_3553;
wire n_2465;
wire n_2275;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_3699;
wire n_4913;
wire n_2312;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_2042;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_1770;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_4089;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_3264;
wire n_2010;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_4865;
wire n_2043;
wire n_3206;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1819;
wire n_3555;
wire n_3155;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1958;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_3301;
wire n_4241;
wire n_1853;
wire n_2324;
wire n_2977;
wire n_1739;
wire n_2847;
wire n_2557;
wire n_2405;
wire n_4050;
wire n_2647;
wire n_2336;
wire n_2521;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1985;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2603;
wire n_2090;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_5022;
wire n_3296;
wire n_2551;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_3822;
wire n_4163;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_4372;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_5108;
wire n_4032;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_3419;
wire n_4478;
wire n_1662;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_4673;
wire n_2519;
wire n_3415;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_2165;
wire n_2750;
wire n_2775;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_3953;
wire n_4588;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_4019;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_4330;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_2316;
wire n_1771;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_2771;
wire n_3020;
wire n_4525;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_2372;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_3196;
wire n_2504;
wire n_2623;
wire n_2063;
wire n_5005;
wire n_2475;
wire n_5181;
wire n_3144;
wire n_3244;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2357;
wire n_2025;
wire n_4654;
wire n_3640;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_2648;
wire n_3212;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1806;
wire n_2023;
wire n_2720;
wire n_2204;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_2627;
wire n_4422;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_2278;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_5189;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_3628;
wire n_4734;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_2704;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_2479;
wire n_1823;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_5004;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_2759;
wire n_2361;
wire n_2266;
wire n_4876;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_1794;
wire n_4493;
wire n_4924;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_4953;
wire n_2944;
wire n_2348;
wire n_3831;
wire n_5167;
wire n_3589;
wire n_2066;
wire n_3391;
wire n_1800;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_4494;
wire n_2380;
wire n_4786;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_4282;
wire n_3493;
wire n_3774;
wire n_2910;
wire n_3268;
wire n_1785;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_2287;
wire n_2492;
wire n_3778;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_3334;
wire n_5097;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_4059;
wire n_4121;
wire n_3290;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_2600;
wire n_3508;
wire n_4353;
wire n_4787;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_2440;
wire n_3521;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_2909;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_4210;
wire n_4981;
wire n_2891;
wire n_2709;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_3945;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

CKINVDCx16_ASAP7_75t_R g1587 ( 
.A(n_1086),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1443),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1500),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_59),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1154),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1422),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_259),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1347),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_249),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1462),
.Y(n_1596)
);

BUFx10_ASAP7_75t_L g1597 ( 
.A(n_1052),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_592),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1433),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_66),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1356),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1103),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1518),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_303),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1490),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1461),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1425),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1211),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_188),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_488),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_683),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_645),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1532),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_472),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1480),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_440),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_590),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1125),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_478),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_904),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_223),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1516),
.Y(n_1622)
);

BUFx8_ASAP7_75t_SL g1623 ( 
.A(n_1416),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1361),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_337),
.Y(n_1625)
);

CKINVDCx20_ASAP7_75t_R g1626 ( 
.A(n_1268),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_257),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1166),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_836),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_73),
.Y(n_1630)
);

BUFx10_ASAP7_75t_L g1631 ( 
.A(n_511),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1261),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1173),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_937),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_421),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_501),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_560),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1300),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_799),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1087),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1450),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_184),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1491),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1331),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1470),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1517),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_37),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1497),
.Y(n_1648)
);

BUFx10_ASAP7_75t_L g1649 ( 
.A(n_1526),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_158),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1468),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_355),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_851),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1435),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1148),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_599),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_473),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_780),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1123),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1373),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_699),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1181),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_875),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_454),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_769),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1115),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_701),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_11),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1391),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_380),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_744),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_570),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1494),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_567),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1477),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_923),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_266),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_557),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_107),
.Y(n_1679)
);

BUFx10_ASAP7_75t_L g1680 ( 
.A(n_252),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1337),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1405),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1178),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_263),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1421),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_592),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_682),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1003),
.Y(n_1688)
);

BUFx5_ASAP7_75t_L g1689 ( 
.A(n_1317),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_302),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1227),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_460),
.Y(n_1692)
);

CKINVDCx16_ASAP7_75t_R g1693 ( 
.A(n_171),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1261),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_692),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_845),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_151),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1486),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_229),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1448),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_855),
.Y(n_1701)
);

BUFx8_ASAP7_75t_SL g1702 ( 
.A(n_581),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1392),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_718),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1374),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1134),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_664),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_933),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_638),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_624),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_275),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1453),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1082),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1510),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1122),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_558),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_382),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_270),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1268),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1484),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_56),
.Y(n_1721)
);

CKINVDCx20_ASAP7_75t_R g1722 ( 
.A(n_1458),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1548),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_745),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1506),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_800),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_370),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_524),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1513),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1011),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_995),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_106),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1229),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_136),
.Y(n_1734)
);

CKINVDCx16_ASAP7_75t_R g1735 ( 
.A(n_1372),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1178),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1482),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1547),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_753),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1133),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1446),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1028),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_249),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_187),
.Y(n_1744)
);

CKINVDCx16_ASAP7_75t_R g1745 ( 
.A(n_983),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_54),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_561),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_171),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1216),
.Y(n_1749)
);

BUFx10_ASAP7_75t_L g1750 ( 
.A(n_746),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_135),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_450),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_371),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1437),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_861),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_378),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_635),
.Y(n_1757)
);

BUFx10_ASAP7_75t_L g1758 ( 
.A(n_1157),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1011),
.Y(n_1759)
);

CKINVDCx20_ASAP7_75t_R g1760 ( 
.A(n_839),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_171),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1175),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1584),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_85),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1505),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_116),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_586),
.Y(n_1767)
);

BUFx5_ASAP7_75t_L g1768 ( 
.A(n_923),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1111),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_766),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1395),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1030),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_877),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_765),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_356),
.Y(n_1775)
);

CKINVDCx14_ASAP7_75t_R g1776 ( 
.A(n_1488),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1402),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_798),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_556),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_768),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1447),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_180),
.Y(n_1782)
);

CKINVDCx14_ASAP7_75t_R g1783 ( 
.A(n_837),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1063),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1151),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_614),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1092),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1210),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_345),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1512),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_352),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_425),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1572),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1488),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_535),
.Y(n_1795)
);

CKINVDCx14_ASAP7_75t_R g1796 ( 
.A(n_661),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1180),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1222),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_213),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1537),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1555),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_126),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1144),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_76),
.Y(n_1804)
);

CKINVDCx16_ASAP7_75t_R g1805 ( 
.A(n_686),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_186),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1483),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1529),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1286),
.Y(n_1809)
);

CKINVDCx14_ASAP7_75t_R g1810 ( 
.A(n_1505),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_94),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1293),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_785),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1173),
.Y(n_1814)
);

CKINVDCx20_ASAP7_75t_R g1815 ( 
.A(n_1441),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_228),
.Y(n_1816)
);

BUFx10_ASAP7_75t_L g1817 ( 
.A(n_51),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1474),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1006),
.Y(n_1819)
);

CKINVDCx20_ASAP7_75t_R g1820 ( 
.A(n_976),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1404),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_349),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_829),
.Y(n_1823)
);

CKINVDCx20_ASAP7_75t_R g1824 ( 
.A(n_422),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_561),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_21),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_427),
.Y(n_1827)
);

CKINVDCx16_ASAP7_75t_R g1828 ( 
.A(n_1262),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_388),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_35),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_690),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1182),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_372),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_221),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_990),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_476),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1579),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1525),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1234),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_278),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_392),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1321),
.Y(n_1842)
);

BUFx2_ASAP7_75t_SL g1843 ( 
.A(n_1278),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1524),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1530),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1454),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1457),
.Y(n_1847)
);

BUFx10_ASAP7_75t_L g1848 ( 
.A(n_1209),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_18),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_319),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_791),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1035),
.Y(n_1852)
);

INVx3_ASAP7_75t_L g1853 ( 
.A(n_1131),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1233),
.Y(n_1854)
);

CKINVDCx16_ASAP7_75t_R g1855 ( 
.A(n_335),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_953),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1288),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1567),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_184),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_782),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1348),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_673),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_199),
.Y(n_1863)
);

INVx2_ASAP7_75t_SL g1864 ( 
.A(n_1198),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_567),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1022),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_997),
.Y(n_1867)
);

CKINVDCx20_ASAP7_75t_R g1868 ( 
.A(n_483),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_907),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_56),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_1321),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1477),
.Y(n_1872)
);

BUFx10_ASAP7_75t_L g1873 ( 
.A(n_96),
.Y(n_1873)
);

CKINVDCx20_ASAP7_75t_R g1874 ( 
.A(n_1446),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_386),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1114),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1333),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1514),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1533),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1444),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_191),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_819),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1216),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1078),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_779),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_499),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_501),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1033),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_544),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_712),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1469),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_767),
.Y(n_1892)
);

CKINVDCx16_ASAP7_75t_R g1893 ( 
.A(n_324),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_428),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_776),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_457),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_328),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1310),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_691),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_306),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_938),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_269),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1409),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1272),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1565),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1279),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_442),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1564),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1466),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_256),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1513),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_357),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1023),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1026),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1352),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1517),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_257),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_189),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_62),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_286),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_0),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1149),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1502),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_47),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_784),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_1317),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1164),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1406),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_724),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_621),
.Y(n_1930)
);

CKINVDCx20_ASAP7_75t_R g1931 ( 
.A(n_1353),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_935),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1031),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_227),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1342),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1460),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1116),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1424),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1433),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1253),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1411),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1200),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1071),
.Y(n_1943)
);

CKINVDCx14_ASAP7_75t_R g1944 ( 
.A(n_88),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_414),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1264),
.Y(n_1946)
);

BUFx10_ASAP7_75t_L g1947 ( 
.A(n_768),
.Y(n_1947)
);

BUFx3_ASAP7_75t_L g1948 ( 
.A(n_1463),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_795),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_571),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_367),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1439),
.Y(n_1952)
);

INVx1_ASAP7_75t_SL g1953 ( 
.A(n_493),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_777),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_469),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_117),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1218),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_426),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_61),
.Y(n_1959)
);

CKINVDCx20_ASAP7_75t_R g1960 ( 
.A(n_262),
.Y(n_1960)
);

CKINVDCx20_ASAP7_75t_R g1961 ( 
.A(n_996),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_903),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_521),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_302),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1008),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1501),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_333),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1156),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1438),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_803),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_157),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_314),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_680),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_277),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1155),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_189),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_375),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_674),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_471),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1290),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_596),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_176),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_609),
.Y(n_1983)
);

CKINVDCx14_ASAP7_75t_R g1984 ( 
.A(n_871),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_306),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_797),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1522),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_186),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1456),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_616),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_1311),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_615),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_765),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1201),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1481),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_403),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_420),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_804),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_220),
.Y(n_1999)
);

CKINVDCx20_ASAP7_75t_R g2000 ( 
.A(n_1425),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_979),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1188),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_861),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_11),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_905),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1418),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_93),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1429),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_358),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1143),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1511),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_601),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_488),
.Y(n_2013)
);

CKINVDCx16_ASAP7_75t_R g2014 ( 
.A(n_779),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_58),
.Y(n_2015)
);

BUFx10_ASAP7_75t_L g2016 ( 
.A(n_1487),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1528),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_965),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_433),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1116),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1379),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1213),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1436),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1459),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1540),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_1285),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1434),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_799),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_463),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1187),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_474),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_306),
.Y(n_2032)
);

CKINVDCx20_ASAP7_75t_R g2033 ( 
.A(n_1185),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_534),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_265),
.Y(n_2035)
);

BUFx10_ASAP7_75t_L g2036 ( 
.A(n_256),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1483),
.Y(n_2037)
);

CKINVDCx20_ASAP7_75t_R g2038 ( 
.A(n_1230),
.Y(n_2038)
);

CKINVDCx20_ASAP7_75t_R g2039 ( 
.A(n_812),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_1052),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_719),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1314),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1121),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_645),
.Y(n_2044)
);

CKINVDCx14_ASAP7_75t_R g2045 ( 
.A(n_1523),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_377),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_842),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_738),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_496),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_955),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_487),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1021),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1168),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1476),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1473),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_976),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_172),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1287),
.Y(n_2058)
);

BUFx3_ASAP7_75t_L g2059 ( 
.A(n_1412),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_926),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_1428),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_9),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1289),
.Y(n_2063)
);

INVx2_ASAP7_75t_SL g2064 ( 
.A(n_216),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1464),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1029),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_870),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1509),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_77),
.Y(n_2069)
);

CKINVDCx20_ASAP7_75t_R g2070 ( 
.A(n_1158),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1504),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_83),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1229),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_594),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1410),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1420),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_406),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_109),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_905),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_493),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_290),
.Y(n_2081)
);

CKINVDCx16_ASAP7_75t_R g2082 ( 
.A(n_686),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1143),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_39),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_919),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1032),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1496),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1182),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_228),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_1478),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1256),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_748),
.Y(n_2092)
);

CKINVDCx20_ASAP7_75t_R g2093 ( 
.A(n_1183),
.Y(n_2093)
);

INVx1_ASAP7_75t_SL g2094 ( 
.A(n_448),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_1493),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_364),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_126),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1361),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_917),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1451),
.Y(n_2100)
);

BUFx5_ASAP7_75t_L g2101 ( 
.A(n_223),
.Y(n_2101)
);

INVx2_ASAP7_75t_SL g2102 ( 
.A(n_1414),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_312),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_789),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_778),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1091),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_281),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_989),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_610),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_1471),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_822),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_53),
.Y(n_2112)
);

CKINVDCx20_ASAP7_75t_R g2113 ( 
.A(n_450),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_849),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1308),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_335),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_528),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_856),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1208),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_192),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_1230),
.Y(n_2121)
);

BUFx3_ASAP7_75t_L g2122 ( 
.A(n_739),
.Y(n_2122)
);

BUFx10_ASAP7_75t_L g2123 ( 
.A(n_689),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1401),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_522),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1521),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_869),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_350),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_920),
.Y(n_2129)
);

BUFx3_ASAP7_75t_L g2130 ( 
.A(n_1418),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1282),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_1040),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_1379),
.Y(n_2133)
);

BUFx6f_ASAP7_75t_L g2134 ( 
.A(n_565),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_182),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_537),
.Y(n_2136)
);

BUFx6f_ASAP7_75t_L g2137 ( 
.A(n_415),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1527),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_693),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_646),
.Y(n_2140)
);

BUFx5_ASAP7_75t_L g2141 ( 
.A(n_848),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1174),
.Y(n_2142)
);

CKINVDCx16_ASAP7_75t_R g2143 ( 
.A(n_1076),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_834),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_741),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_217),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1478),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_632),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1378),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1273),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1578),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_998),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1440),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_130),
.Y(n_2154)
);

CKINVDCx20_ASAP7_75t_R g2155 ( 
.A(n_1536),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1495),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1485),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1214),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_648),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1413),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_513),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1239),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1426),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_533),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_18),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_L g2166 ( 
.A(n_346),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1081),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_398),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_573),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1017),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_1124),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_416),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_1489),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1121),
.Y(n_2174)
);

BUFx10_ASAP7_75t_L g2175 ( 
.A(n_1492),
.Y(n_2175)
);

INVx2_ASAP7_75t_SL g2176 ( 
.A(n_468),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_1375),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1549),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1355),
.Y(n_2179)
);

BUFx5_ASAP7_75t_L g2180 ( 
.A(n_85),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1507),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_608),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1427),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1267),
.Y(n_2184)
);

HB1xp67_ASAP7_75t_L g2185 ( 
.A(n_467),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1499),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_911),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1123),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_351),
.Y(n_2189)
);

BUFx3_ASAP7_75t_L g2190 ( 
.A(n_1179),
.Y(n_2190)
);

BUFx6f_ASAP7_75t_L g2191 ( 
.A(n_903),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_649),
.Y(n_2192)
);

BUFx3_ASAP7_75t_L g2193 ( 
.A(n_28),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_262),
.Y(n_2194)
);

BUFx8_ASAP7_75t_SL g2195 ( 
.A(n_668),
.Y(n_2195)
);

BUFx3_ASAP7_75t_L g2196 ( 
.A(n_1531),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1487),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1106),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_206),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_410),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_102),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1105),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_472),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_757),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_274),
.Y(n_2206)
);

CKINVDCx5p33_ASAP7_75t_R g2207 ( 
.A(n_60),
.Y(n_2207)
);

BUFx10_ASAP7_75t_L g2208 ( 
.A(n_412),
.Y(n_2208)
);

CKINVDCx5p33_ASAP7_75t_R g2209 ( 
.A(n_1415),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1442),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_895),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_760),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1394),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1408),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_579),
.Y(n_2215)
);

CKINVDCx16_ASAP7_75t_R g2216 ( 
.A(n_1445),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_436),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1050),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1054),
.Y(n_2219)
);

CKINVDCx20_ASAP7_75t_R g2220 ( 
.A(n_316),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_470),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1579),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1403),
.Y(n_2223)
);

CKINVDCx16_ASAP7_75t_R g2224 ( 
.A(n_816),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_834),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_1498),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_1503),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_310),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_1562),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_1126),
.Y(n_2230)
);

INVxp67_ASAP7_75t_L g2231 ( 
.A(n_712),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_971),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_657),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_243),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_1508),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1452),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_933),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_6),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_416),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1283),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1336),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_272),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_754),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_952),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1467),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_930),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1010),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1423),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1449),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_332),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_560),
.Y(n_2251)
);

CKINVDCx20_ASAP7_75t_R g2252 ( 
.A(n_377),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_110),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1212),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1472),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_1534),
.Y(n_2256)
);

BUFx2_ASAP7_75t_SL g2257 ( 
.A(n_199),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1463),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_1430),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_419),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1455),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_115),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1535),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1432),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_999),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1542),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_558),
.Y(n_2267)
);

CKINVDCx20_ASAP7_75t_R g2268 ( 
.A(n_988),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_945),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_1001),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_423),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_443),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_583),
.Y(n_2273)
);

INVxp33_ASAP7_75t_L g2274 ( 
.A(n_762),
.Y(n_2274)
);

CKINVDCx20_ASAP7_75t_R g2275 ( 
.A(n_562),
.Y(n_2275)
);

CKINVDCx20_ASAP7_75t_R g2276 ( 
.A(n_835),
.Y(n_2276)
);

CKINVDCx20_ASAP7_75t_R g2277 ( 
.A(n_1469),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1550),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_432),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_724),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_1515),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_665),
.Y(n_2282)
);

CKINVDCx20_ASAP7_75t_R g2283 ( 
.A(n_1557),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_563),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1098),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_421),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_1071),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1059),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1291),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_622),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_1129),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_961),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_583),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_703),
.Y(n_2294)
);

BUFx3_ASAP7_75t_L g2295 ( 
.A(n_955),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_837),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_825),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1419),
.Y(n_2298)
);

CKINVDCx16_ASAP7_75t_R g2299 ( 
.A(n_101),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_943),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_824),
.Y(n_2301)
);

BUFx6f_ASAP7_75t_L g2302 ( 
.A(n_1519),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_1256),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_867),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_826),
.Y(n_2305)
);

CKINVDCx20_ASAP7_75t_R g2306 ( 
.A(n_740),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1376),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1404),
.Y(n_2308)
);

CKINVDCx16_ASAP7_75t_R g2309 ( 
.A(n_1180),
.Y(n_2309)
);

INVx3_ASAP7_75t_L g2310 ( 
.A(n_697),
.Y(n_2310)
);

BUFx2_ASAP7_75t_L g2311 ( 
.A(n_1048),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_239),
.Y(n_2312)
);

CKINVDCx20_ASAP7_75t_R g2313 ( 
.A(n_1417),
.Y(n_2313)
);

CKINVDCx20_ASAP7_75t_R g2314 ( 
.A(n_74),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_967),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1050),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_704),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_550),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_879),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1060),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_893),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_56),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_299),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1563),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_784),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_900),
.Y(n_2326)
);

BUFx5_ASAP7_75t_L g2327 ( 
.A(n_671),
.Y(n_2327)
);

BUFx5_ASAP7_75t_L g2328 ( 
.A(n_1313),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_125),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_21),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_132),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_832),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_1465),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_135),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_1528),
.Y(n_2335)
);

CKINVDCx16_ASAP7_75t_R g2336 ( 
.A(n_939),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_545),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_705),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_1174),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_576),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1319),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_251),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1328),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_508),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_1479),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_602),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_1159),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1520),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_357),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1431),
.Y(n_2350)
);

BUFx10_ASAP7_75t_L g2351 ( 
.A(n_356),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_511),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_1085),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_1407),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_625),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1318),
.Y(n_2356)
);

INVxp67_ASAP7_75t_L g2357 ( 
.A(n_94),
.Y(n_2357)
);

CKINVDCx5p33_ASAP7_75t_R g2358 ( 
.A(n_474),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_223),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1475),
.Y(n_2360)
);

BUFx5_ASAP7_75t_L g2361 ( 
.A(n_1585),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_1623),
.Y(n_2362)
);

INVxp33_ASAP7_75t_SL g2363 ( 
.A(n_1610),
.Y(n_2363)
);

INVxp67_ASAP7_75t_SL g2364 ( 
.A(n_1677),
.Y(n_2364)
);

INVxp33_ASAP7_75t_SL g2365 ( 
.A(n_1723),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2101),
.Y(n_2366)
);

INVxp67_ASAP7_75t_SL g2367 ( 
.A(n_1677),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2180),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2180),
.Y(n_2369)
);

INVxp67_ASAP7_75t_SL g2370 ( 
.A(n_1917),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2180),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2180),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_1944),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1689),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_1643),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_1702),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1689),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1689),
.Y(n_2378)
);

CKINVDCx20_ASAP7_75t_R g2379 ( 
.A(n_1776),
.Y(n_2379)
);

INVxp33_ASAP7_75t_L g2380 ( 
.A(n_1832),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_2195),
.Y(n_2381)
);

INVxp67_ASAP7_75t_L g2382 ( 
.A(n_1645),
.Y(n_2382)
);

CKINVDCx16_ASAP7_75t_R g2383 ( 
.A(n_1693),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1689),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1689),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1768),
.Y(n_2386)
);

BUFx3_ASAP7_75t_L g2387 ( 
.A(n_1834),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1768),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2141),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2141),
.Y(n_2390)
);

INVxp33_ASAP7_75t_SL g2391 ( 
.A(n_1833),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2141),
.Y(n_2392)
);

CKINVDCx16_ASAP7_75t_R g2393 ( 
.A(n_1855),
.Y(n_2393)
);

NOR2xp67_ASAP7_75t_L g2394 ( 
.A(n_1615),
.B(n_0),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_1893),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2299),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2141),
.Y(n_2397)
);

INVxp67_ASAP7_75t_L g2398 ( 
.A(n_1737),
.Y(n_2398)
);

CKINVDCx5p33_ASAP7_75t_R g2399 ( 
.A(n_1783),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2141),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2327),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2327),
.Y(n_2402)
);

CKINVDCx20_ASAP7_75t_R g2403 ( 
.A(n_1796),
.Y(n_2403)
);

INVxp33_ASAP7_75t_SL g2404 ( 
.A(n_1845),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_1810),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2327),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2327),
.Y(n_2407)
);

BUFx2_ASAP7_75t_L g2408 ( 
.A(n_1756),
.Y(n_2408)
);

INVxp67_ASAP7_75t_SL g2409 ( 
.A(n_1853),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2328),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2328),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2328),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2361),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2361),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2361),
.Y(n_2415)
);

INVxp67_ASAP7_75t_L g2416 ( 
.A(n_1779),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2361),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2359),
.Y(n_2418)
);

INVx1_ASAP7_75t_SL g2419 ( 
.A(n_1825),
.Y(n_2419)
);

CKINVDCx16_ASAP7_75t_R g2420 ( 
.A(n_1587),
.Y(n_2420)
);

CKINVDCx20_ASAP7_75t_R g2421 ( 
.A(n_1984),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_2045),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1593),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1604),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1609),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1630),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_1642),
.Y(n_2427)
);

INVxp67_ASAP7_75t_L g2428 ( 
.A(n_2049),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1690),
.Y(n_2429)
);

CKINVDCx16_ASAP7_75t_R g2430 ( 
.A(n_1735),
.Y(n_2430)
);

CKINVDCx14_ASAP7_75t_R g2431 ( 
.A(n_2108),
.Y(n_2431)
);

INVxp67_ASAP7_75t_SL g2432 ( 
.A(n_1853),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1697),
.Y(n_2433)
);

INVxp67_ASAP7_75t_SL g2434 ( 
.A(n_2017),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1711),
.Y(n_2435)
);

CKINVDCx20_ASAP7_75t_R g2436 ( 
.A(n_1745),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_1805),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1718),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1744),
.Y(n_2439)
);

INVxp33_ASAP7_75t_SL g2440 ( 
.A(n_1978),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_1746),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_1782),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1799),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1804),
.Y(n_2444)
);

CKINVDCx16_ASAP7_75t_R g2445 ( 
.A(n_1828),
.Y(n_2445)
);

INVxp67_ASAP7_75t_L g2446 ( 
.A(n_2311),
.Y(n_2446)
);

INVxp67_ASAP7_75t_L g2447 ( 
.A(n_2162),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1816),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_1849),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_1850),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_1900),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_1919),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1934),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_1956),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1959),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1964),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1974),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2015),
.Y(n_2458)
);

INVxp33_ASAP7_75t_L g2459 ( 
.A(n_2185),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2035),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_1764),
.Y(n_2461)
);

CKINVDCx16_ASAP7_75t_R g2462 ( 
.A(n_2014),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_1588),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2072),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2078),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2089),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2103),
.Y(n_2467)
);

INVxp67_ASAP7_75t_L g2468 ( 
.A(n_2227),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2146),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2198),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_1764),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2242),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2253),
.Y(n_2473)
);

INVxp33_ASAP7_75t_L g2474 ( 
.A(n_2312),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2322),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2334),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2193),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_1764),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_1811),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_1811),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_1811),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2082),
.Y(n_2482)
);

CKINVDCx20_ASAP7_75t_R g2483 ( 
.A(n_2143),
.Y(n_2483)
);

INVxp67_ASAP7_75t_SL g2484 ( 
.A(n_2310),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2216),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_2224),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_2309),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_1999),
.Y(n_2488)
);

INVxp67_ASAP7_75t_SL g2489 ( 
.A(n_2310),
.Y(n_2489)
);

CKINVDCx16_ASAP7_75t_R g2490 ( 
.A(n_2336),
.Y(n_2490)
);

CKINVDCx16_ASAP7_75t_R g2491 ( 
.A(n_1680),
.Y(n_2491)
);

CKINVDCx20_ASAP7_75t_R g2492 ( 
.A(n_1620),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_L g2493 ( 
.A(n_1999),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_1621),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_1684),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_1721),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_1918),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2004),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2107),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2228),
.Y(n_2500)
);

INVxp67_ASAP7_75t_L g2501 ( 
.A(n_1680),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_1588),
.Y(n_2502)
);

INVxp67_ASAP7_75t_SL g2503 ( 
.A(n_1588),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_1590),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_1589),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_1595),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_1658),
.Y(n_2507)
);

INVxp67_ASAP7_75t_SL g2508 ( 
.A(n_1700),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_1822),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_1822),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_1822),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_1872),
.Y(n_2512)
);

INVxp67_ASAP7_75t_SL g2513 ( 
.A(n_1872),
.Y(n_2513)
);

INVx2_ASAP7_75t_SL g2514 ( 
.A(n_1817),
.Y(n_2514)
);

BUFx2_ASAP7_75t_L g2515 ( 
.A(n_1600),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_1625),
.Y(n_2516)
);

CKINVDCx16_ASAP7_75t_R g2517 ( 
.A(n_1873),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_1907),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_1907),
.Y(n_2519)
);

CKINVDCx20_ASAP7_75t_R g2520 ( 
.A(n_1626),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1981),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_1981),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1981),
.Y(n_2523)
);

INVxp67_ASAP7_75t_L g2524 ( 
.A(n_1873),
.Y(n_2524)
);

INVxp33_ASAP7_75t_L g2525 ( 
.A(n_2274),
.Y(n_2525)
);

INVxp67_ASAP7_75t_L g2526 ( 
.A(n_2036),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2026),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2027),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2086),
.Y(n_2529)
);

INVxp33_ASAP7_75t_SL g2530 ( 
.A(n_1647),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2086),
.Y(n_2531)
);

BUFx2_ASAP7_75t_L g2532 ( 
.A(n_1668),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2134),
.Y(n_2533)
);

INVxp33_ASAP7_75t_SL g2534 ( 
.A(n_1679),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2137),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2137),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_1699),
.Y(n_2537)
);

BUFx3_ASAP7_75t_L g2538 ( 
.A(n_1644),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2166),
.Y(n_2539)
);

INVxp33_ASAP7_75t_L g2540 ( 
.A(n_1591),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2191),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2191),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2191),
.Y(n_2543)
);

INVxp67_ASAP7_75t_L g2544 ( 
.A(n_1597),
.Y(n_2544)
);

INVxp33_ASAP7_75t_L g2545 ( 
.A(n_1594),
.Y(n_2545)
);

CKINVDCx16_ASAP7_75t_R g2546 ( 
.A(n_1631),
.Y(n_2546)
);

INVxp67_ASAP7_75t_L g2547 ( 
.A(n_1649),
.Y(n_2547)
);

BUFx3_ASAP7_75t_L g2548 ( 
.A(n_1736),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2203),
.Y(n_2549)
);

CKINVDCx16_ASAP7_75t_R g2550 ( 
.A(n_1750),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2530),
.B(n_1627),
.Y(n_2551)
);

INVxp33_ASAP7_75t_SL g2552 ( 
.A(n_2362),
.Y(n_2552)
);

BUFx8_ASAP7_75t_SL g2553 ( 
.A(n_2376),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2512),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2533),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2364),
.B(n_2302),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2503),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2363),
.A2(n_1732),
.B1(n_1748),
.B2(n_1734),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2461),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2508),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2513),
.Y(n_2561)
);

INVx4_ASAP7_75t_L g2562 ( 
.A(n_2399),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2367),
.B(n_2302),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2365),
.A2(n_1751),
.B1(n_1766),
.B2(n_1761),
.Y(n_2564)
);

INVx6_ASAP7_75t_L g2565 ( 
.A(n_2387),
.Y(n_2565)
);

XNOR2xp5_ASAP7_75t_L g2566 ( 
.A(n_2492),
.B(n_1650),
.Y(n_2566)
);

INVx3_ASAP7_75t_L g2567 ( 
.A(n_2471),
.Y(n_2567)
);

OAI21x1_ASAP7_75t_L g2568 ( 
.A1(n_2366),
.A2(n_1694),
.B(n_1687),
.Y(n_2568)
);

OAI22x1_ASAP7_75t_SL g2569 ( 
.A1(n_2520),
.A2(n_1897),
.B1(n_1960),
.B2(n_1802),
.Y(n_2569)
);

AND2x4_ASAP7_75t_L g2570 ( 
.A(n_2373),
.B(n_1778),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2471),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2471),
.Y(n_2572)
);

OAI21x1_ASAP7_75t_L g2573 ( 
.A1(n_2368),
.A2(n_2371),
.B(n_2369),
.Y(n_2573)
);

AND2x4_ASAP7_75t_L g2574 ( 
.A(n_2370),
.B(n_1791),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2481),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2534),
.B(n_1743),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2405),
.B(n_2064),
.Y(n_2577)
);

AND2x4_ASAP7_75t_L g2578 ( 
.A(n_2382),
.B(n_1846),
.Y(n_2578)
);

BUFx2_ASAP7_75t_L g2579 ( 
.A(n_2436),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2422),
.B(n_1806),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2372),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2483),
.Y(n_2582)
);

BUFx6f_ASAP7_75t_L g2583 ( 
.A(n_2481),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2409),
.B(n_1753),
.Y(n_2584)
);

INVx4_ASAP7_75t_L g2585 ( 
.A(n_2504),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2481),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2478),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2493),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2432),
.B(n_1835),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2525),
.B(n_1906),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2398),
.B(n_1916),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2479),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2434),
.B(n_1864),
.Y(n_2593)
);

OAI22xp5_ASAP7_75t_SL g2594 ( 
.A1(n_2383),
.A2(n_2314),
.B1(n_2220),
.B2(n_1666),
.Y(n_2594)
);

AND2x4_ASAP7_75t_L g2595 ( 
.A(n_2416),
.B(n_1948),
.Y(n_2595)
);

NOR2x1_ASAP7_75t_L g2596 ( 
.A(n_2374),
.B(n_1951),
.Y(n_2596)
);

BUFx12f_ASAP7_75t_L g2597 ( 
.A(n_2381),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_L g2598 ( 
.A(n_2391),
.B(n_2404),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2428),
.B(n_1980),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2493),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2480),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2485),
.Y(n_2602)
);

BUFx8_ASAP7_75t_L g2603 ( 
.A(n_2408),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2463),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2463),
.Y(n_2605)
);

BUFx3_ASAP7_75t_L g2606 ( 
.A(n_2505),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2488),
.Y(n_2607)
);

INVx2_ASAP7_75t_SL g2608 ( 
.A(n_2506),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2442),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2502),
.Y(n_2610)
);

OR2x2_ASAP7_75t_L g2611 ( 
.A(n_2375),
.B(n_1971),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2507),
.Y(n_2612)
);

OA21x2_ASAP7_75t_L g2613 ( 
.A1(n_2377),
.A2(n_1704),
.B(n_1703),
.Y(n_2613)
);

BUFx12f_ASAP7_75t_L g2614 ( 
.A(n_2486),
.Y(n_2614)
);

BUFx6f_ASAP7_75t_L g2615 ( 
.A(n_2444),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_SL g2616 ( 
.A(n_2420),
.B(n_1826),
.Y(n_2616)
);

BUFx6f_ASAP7_75t_L g2617 ( 
.A(n_2450),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2509),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2510),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2511),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_2452),
.Y(n_2621)
);

BUFx3_ASAP7_75t_L g2622 ( 
.A(n_2538),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2518),
.Y(n_2623)
);

BUFx6f_ASAP7_75t_L g2624 ( 
.A(n_2548),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2519),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2521),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2522),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2523),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_2477),
.Y(n_2629)
);

BUFx6f_ASAP7_75t_L g2630 ( 
.A(n_2500),
.Y(n_2630)
);

INVx6_ASAP7_75t_L g2631 ( 
.A(n_2491),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_2440),
.B(n_1830),
.Y(n_2632)
);

CKINVDCx6p67_ASAP7_75t_R g2633 ( 
.A(n_2379),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2527),
.Y(n_2634)
);

BUFx2_ASAP7_75t_L g2635 ( 
.A(n_2403),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2487),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_2528),
.Y(n_2637)
);

HB1xp67_ASAP7_75t_L g2638 ( 
.A(n_2395),
.Y(n_2638)
);

BUFx8_ASAP7_75t_L g2639 ( 
.A(n_2514),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2529),
.Y(n_2640)
);

AOI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_2396),
.A2(n_1840),
.B1(n_1863),
.B2(n_1859),
.Y(n_2641)
);

INVx3_ASAP7_75t_L g2642 ( 
.A(n_2531),
.Y(n_2642)
);

AOI22x1_ASAP7_75t_SL g2643 ( 
.A1(n_2421),
.A2(n_1709),
.B1(n_1720),
.B2(n_1696),
.Y(n_2643)
);

OA21x2_ASAP7_75t_L g2644 ( 
.A1(n_2378),
.A2(n_1715),
.B(n_1707),
.Y(n_2644)
);

OAI21x1_ASAP7_75t_L g2645 ( 
.A1(n_2414),
.A2(n_1755),
.B(n_1728),
.Y(n_2645)
);

AND2x6_ASAP7_75t_L g2646 ( 
.A(n_2419),
.B(n_1985),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2535),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2516),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2536),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2484),
.B(n_2059),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2539),
.Y(n_2651)
);

AOI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2393),
.A2(n_1870),
.B1(n_1902),
.B2(n_1881),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_2541),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_SL g2654 ( 
.A1(n_2431),
.A2(n_1747),
.B1(n_1760),
.B2(n_1722),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_2542),
.Y(n_2655)
);

BUFx6f_ASAP7_75t_L g2656 ( 
.A(n_2543),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2549),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2418),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2423),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2384),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2424),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2385),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2425),
.Y(n_2663)
);

BUFx6f_ASAP7_75t_L g2664 ( 
.A(n_2426),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2386),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2489),
.B(n_2110),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2537),
.B(n_2030),
.Y(n_2667)
);

NOR2xp33_ASAP7_75t_SL g2668 ( 
.A(n_2430),
.B(n_2445),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2388),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_2427),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2515),
.B(n_2122),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2429),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2389),
.Y(n_2673)
);

BUFx3_ASAP7_75t_L g2674 ( 
.A(n_2390),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2392),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2397),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2532),
.B(n_2130),
.Y(n_2677)
);

BUFx2_ASAP7_75t_L g2678 ( 
.A(n_2437),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2400),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2401),
.Y(n_2680)
);

AOI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2462),
.A2(n_1910),
.B1(n_1921),
.B2(n_1920),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_L g2682 ( 
.A(n_2433),
.Y(n_2682)
);

BUFx6f_ASAP7_75t_L g2683 ( 
.A(n_2435),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2402),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2446),
.B(n_2164),
.Y(n_2685)
);

BUFx6f_ASAP7_75t_L g2686 ( 
.A(n_2438),
.Y(n_2686)
);

INVx5_ASAP7_75t_L g2687 ( 
.A(n_2546),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2406),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2550),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2407),
.Y(n_2690)
);

INVx4_ASAP7_75t_L g2691 ( 
.A(n_2517),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2410),
.B(n_2061),
.Y(n_2692)
);

BUFx6f_ASAP7_75t_L g2693 ( 
.A(n_2439),
.Y(n_2693)
);

OA21x2_ASAP7_75t_L g2694 ( 
.A1(n_2411),
.A2(n_1763),
.B(n_1757),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2380),
.B(n_2190),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2447),
.B(n_2196),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2412),
.Y(n_2697)
);

INVx3_ASAP7_75t_L g2698 ( 
.A(n_2441),
.Y(n_2698)
);

BUFx6f_ASAP7_75t_L g2699 ( 
.A(n_2443),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2413),
.B(n_2102),
.Y(n_2700)
);

OAI22xp5_ASAP7_75t_L g2701 ( 
.A1(n_2459),
.A2(n_1967),
.B1(n_1972),
.B2(n_1924),
.Y(n_2701)
);

OA21x2_ASAP7_75t_L g2702 ( 
.A1(n_2415),
.A2(n_1818),
.B(n_1781),
.Y(n_2702)
);

BUFx6f_ASAP7_75t_L g2703 ( 
.A(n_2448),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2553),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2611),
.B(n_2490),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2674),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2552),
.Y(n_2707)
);

INVx3_ASAP7_75t_L g2708 ( 
.A(n_2660),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2624),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2659),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2661),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_2633),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2630),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2614),
.Y(n_2714)
);

BUFx3_ASAP7_75t_L g2715 ( 
.A(n_2606),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2559),
.Y(n_2716)
);

AO21x2_ASAP7_75t_L g2717 ( 
.A1(n_2573),
.A2(n_2394),
.B(n_2417),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2663),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_2585),
.Y(n_2719)
);

NOR2xp33_ASAP7_75t_R g2720 ( 
.A(n_2668),
.B(n_2482),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2648),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2664),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2672),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2571),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_2608),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_R g2726 ( 
.A(n_2689),
.B(n_2579),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_2582),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2572),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2566),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2682),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_2635),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2687),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2590),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2588),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_2562),
.Y(n_2735)
);

CKINVDCx20_ASAP7_75t_R g2736 ( 
.A(n_2631),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2639),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2602),
.Y(n_2738)
);

CKINVDCx20_ASAP7_75t_R g2739 ( 
.A(n_2638),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2636),
.Y(n_2740)
);

HB1xp67_ASAP7_75t_L g2741 ( 
.A(n_2695),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2646),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_2622),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2580),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2691),
.Y(n_2745)
);

HB1xp67_ASAP7_75t_L g2746 ( 
.A(n_2678),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2683),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2686),
.Y(n_2748)
);

NOR2xp67_ASAP7_75t_L g2749 ( 
.A(n_2598),
.B(n_2544),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2600),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_2565),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2603),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2632),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2693),
.Y(n_2754)
);

AOI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2551),
.A2(n_2576),
.B1(n_2577),
.B2(n_2681),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2671),
.B(n_2468),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2699),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2703),
.Y(n_2758)
);

BUFx6f_ASAP7_75t_L g2759 ( 
.A(n_2575),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2643),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2581),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_2667),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_2594),
.Y(n_2763)
);

CKINVDCx5p33_ASAP7_75t_R g2764 ( 
.A(n_2569),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2662),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2641),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2554),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2646),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2677),
.Y(n_2769)
);

OAI22xp5_ASAP7_75t_SL g2770 ( 
.A1(n_2654),
.A2(n_1813),
.B1(n_1815),
.B2(n_1793),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2650),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_R g2772 ( 
.A(n_2557),
.B(n_1820),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2665),
.Y(n_2773)
);

CKINVDCx20_ASAP7_75t_R g2774 ( 
.A(n_2616),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2555),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_R g2776 ( 
.A(n_2560),
.B(n_1824),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2669),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_2666),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_2652),
.Y(n_2779)
);

OAI22xp5_ASAP7_75t_SL g2780 ( 
.A1(n_2558),
.A2(n_1838),
.B1(n_1868),
.B2(n_1836),
.Y(n_2780)
);

CKINVDCx20_ASAP7_75t_R g2781 ( 
.A(n_2564),
.Y(n_2781)
);

INVxp67_ASAP7_75t_SL g2782 ( 
.A(n_2556),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_2574),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_2629),
.Y(n_2784)
);

CKINVDCx5p33_ASAP7_75t_R g2785 ( 
.A(n_2701),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2673),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_2561),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2675),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2609),
.Y(n_2789)
);

BUFx6f_ASAP7_75t_L g2790 ( 
.A(n_2583),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2615),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2578),
.B(n_2501),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_R g2793 ( 
.A(n_2584),
.B(n_1871),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_R g2794 ( 
.A(n_2589),
.B(n_1874),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2684),
.Y(n_2795)
);

CKINVDCx5p33_ASAP7_75t_R g2796 ( 
.A(n_2593),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_SL g2797 ( 
.A(n_2570),
.B(n_1926),
.Y(n_2797)
);

CKINVDCx5p33_ASAP7_75t_R g2798 ( 
.A(n_2591),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2595),
.B(n_2524),
.Y(n_2799)
);

CKINVDCx5p33_ASAP7_75t_R g2800 ( 
.A(n_2599),
.Y(n_2800)
);

OR2x2_ASAP7_75t_L g2801 ( 
.A(n_2563),
.B(n_2526),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2690),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2617),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2586),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2697),
.Y(n_2805)
);

BUFx10_ASAP7_75t_L g2806 ( 
.A(n_2685),
.Y(n_2806)
);

BUFx10_ASAP7_75t_L g2807 ( 
.A(n_2696),
.Y(n_2807)
);

CKINVDCx20_ASAP7_75t_R g2808 ( 
.A(n_2653),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_2621),
.Y(n_2809)
);

CKINVDCx5p33_ASAP7_75t_R g2810 ( 
.A(n_2604),
.Y(n_2810)
);

BUFx10_ASAP7_75t_L g2811 ( 
.A(n_2605),
.Y(n_2811)
);

CKINVDCx20_ASAP7_75t_R g2812 ( 
.A(n_2692),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_2640),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2676),
.Y(n_2814)
);

CKINVDCx5p33_ASAP7_75t_R g2815 ( 
.A(n_2656),
.Y(n_2815)
);

INVx3_ASAP7_75t_L g2816 ( 
.A(n_2679),
.Y(n_2816)
);

CKINVDCx20_ASAP7_75t_R g2817 ( 
.A(n_2700),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_2670),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2601),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2680),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2688),
.Y(n_2821)
);

CKINVDCx20_ASAP7_75t_R g2822 ( 
.A(n_2613),
.Y(n_2822)
);

CKINVDCx5p33_ASAP7_75t_R g2823 ( 
.A(n_2698),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2644),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_2618),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_2620),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2694),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2607),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2702),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2596),
.B(n_2474),
.Y(n_2830)
);

CKINVDCx5p33_ASAP7_75t_R g2831 ( 
.A(n_2623),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_2625),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2567),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2587),
.Y(n_2834)
);

BUFx10_ASAP7_75t_L g2835 ( 
.A(n_2592),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2568),
.Y(n_2836)
);

CKINVDCx5p33_ASAP7_75t_R g2837 ( 
.A(n_2626),
.Y(n_2837)
);

BUFx2_ASAP7_75t_L g2838 ( 
.A(n_2637),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_R g2839 ( 
.A(n_2642),
.B(n_1931),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2610),
.Y(n_2840)
);

BUFx3_ASAP7_75t_L g2841 ( 
.A(n_2655),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2649),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2657),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_2612),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2645),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2619),
.Y(n_2846)
);

CKINVDCx16_ASAP7_75t_R g2847 ( 
.A(n_2627),
.Y(n_2847)
);

CKINVDCx20_ASAP7_75t_R g2848 ( 
.A(n_2628),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2634),
.Y(n_2849)
);

CKINVDCx20_ASAP7_75t_R g2850 ( 
.A(n_2647),
.Y(n_2850)
);

BUFx10_ASAP7_75t_L g2851 ( 
.A(n_2651),
.Y(n_2851)
);

CKINVDCx5p33_ASAP7_75t_R g2852 ( 
.A(n_2553),
.Y(n_2852)
);

XNOR2x1_ASAP7_75t_L g2853 ( 
.A(n_2566),
.B(n_1976),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2667),
.B(n_2547),
.Y(n_2854)
);

CKINVDCx20_ASAP7_75t_R g2855 ( 
.A(n_2633),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_2553),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2630),
.Y(n_2857)
);

CKINVDCx20_ASAP7_75t_R g2858 ( 
.A(n_2633),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2658),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_R g2860 ( 
.A(n_2597),
.B(n_1961),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_2553),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_2553),
.Y(n_2862)
);

NAND2xp33_ASAP7_75t_R g2863 ( 
.A(n_2678),
.B(n_1982),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2658),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_R g2865 ( 
.A(n_2597),
.B(n_1965),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2658),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_2553),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2767),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2834),
.Y(n_2869)
);

BUFx6f_ASAP7_75t_L g2870 ( 
.A(n_2759),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2775),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2759),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2709),
.B(n_2449),
.Y(n_2873)
);

AO22x2_ASAP7_75t_L g2874 ( 
.A1(n_2853),
.A2(n_2007),
.B1(n_2257),
.B2(n_1843),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2811),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2840),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2762),
.B(n_2540),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2708),
.Y(n_2878)
);

INVx1_ASAP7_75t_SL g2879 ( 
.A(n_2769),
.Y(n_2879)
);

INVx3_ASAP7_75t_L g2880 ( 
.A(n_2811),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2756),
.B(n_2545),
.Y(n_2881)
);

BUFx6f_ASAP7_75t_L g2882 ( 
.A(n_2759),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_2719),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2816),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2846),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2789),
.B(n_2451),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2819),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2733),
.B(n_2453),
.Y(n_2888)
);

BUFx2_ASAP7_75t_L g2889 ( 
.A(n_2746),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2761),
.Y(n_2890)
);

CKINVDCx16_ASAP7_75t_R g2891 ( 
.A(n_2726),
.Y(n_2891)
);

INVx1_ASAP7_75t_SL g2892 ( 
.A(n_2839),
.Y(n_2892)
);

NAND2xp33_ASAP7_75t_SL g2893 ( 
.A(n_2753),
.B(n_2720),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2854),
.B(n_1657),
.Y(n_2894)
);

OR2x2_ASAP7_75t_L g2895 ( 
.A(n_2705),
.B(n_1683),
.Y(n_2895)
);

OR2x2_ASAP7_75t_L g2896 ( 
.A(n_2801),
.B(n_1706),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2765),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2828),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2741),
.B(n_2454),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2773),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2777),
.Y(n_2901)
);

BUFx6f_ASAP7_75t_L g2902 ( 
.A(n_2790),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2791),
.B(n_2455),
.Y(n_2903)
);

AO22x2_ASAP7_75t_L g2904 ( 
.A1(n_2770),
.A2(n_1740),
.B1(n_1821),
.B2(n_1731),
.Y(n_2904)
);

AND2x4_ASAP7_75t_L g2905 ( 
.A(n_2803),
.B(n_2456),
.Y(n_2905)
);

INVx4_ASAP7_75t_SL g2906 ( 
.A(n_2799),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2786),
.B(n_2176),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2830),
.B(n_2457),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2788),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2744),
.B(n_1953),
.Y(n_2910)
);

INVx3_ASAP7_75t_L g2911 ( 
.A(n_2790),
.Y(n_2911)
);

BUFx6f_ASAP7_75t_L g2912 ( 
.A(n_2804),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2814),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2795),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2804),
.Y(n_2915)
);

AND2x4_ASAP7_75t_L g2916 ( 
.A(n_2841),
.B(n_2458),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2820),
.Y(n_2917)
);

INVx1_ASAP7_75t_SL g2918 ( 
.A(n_2772),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2802),
.B(n_2460),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2805),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2821),
.Y(n_2921)
);

BUFx10_ASAP7_75t_L g2922 ( 
.A(n_2704),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2849),
.Y(n_2923)
);

OAI221xp5_ASAP7_75t_L g2924 ( 
.A1(n_2755),
.A2(n_2357),
.B1(n_1942),
.B2(n_2231),
.C(n_1899),
.Y(n_2924)
);

BUFx10_ASAP7_75t_L g2925 ( 
.A(n_2852),
.Y(n_2925)
);

HB1xp67_ASAP7_75t_L g2926 ( 
.A(n_2771),
.Y(n_2926)
);

NOR2xp33_ASAP7_75t_SL g2927 ( 
.A(n_2725),
.B(n_2714),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2778),
.B(n_1592),
.Y(n_2928)
);

BUFx3_ASAP7_75t_L g2929 ( 
.A(n_2809),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2787),
.B(n_1987),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2706),
.B(n_2464),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2716),
.Y(n_2932)
);

OAI22xp33_ASAP7_75t_L g2933 ( 
.A1(n_2785),
.A2(n_2085),
.B1(n_2099),
.B2(n_2094),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2824),
.B(n_2465),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2804),
.Y(n_2935)
);

INVx2_ASAP7_75t_SL g2936 ( 
.A(n_2807),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2749),
.B(n_2466),
.Y(n_2937)
);

CKINVDCx20_ASAP7_75t_R g2938 ( 
.A(n_2736),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_2807),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2724),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2818),
.B(n_2467),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2728),
.Y(n_2942)
);

INVx3_ASAP7_75t_L g2943 ( 
.A(n_2713),
.Y(n_2943)
);

BUFx3_ASAP7_75t_L g2944 ( 
.A(n_2813),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2734),
.Y(n_2945)
);

INVx5_ASAP7_75t_L g2946 ( 
.A(n_2806),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2827),
.B(n_2469),
.Y(n_2947)
);

INVx2_ASAP7_75t_SL g2948 ( 
.A(n_2806),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2750),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2829),
.Y(n_2950)
);

AND2x4_ASAP7_75t_L g2951 ( 
.A(n_2857),
.B(n_2470),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2833),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2844),
.B(n_1988),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2836),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2838),
.Y(n_2955)
);

AOI22xp33_ASAP7_75t_L g2956 ( 
.A1(n_2822),
.A2(n_1884),
.B1(n_1888),
.B2(n_1877),
.Y(n_2956)
);

AND2x6_ASAP7_75t_L g2957 ( 
.A(n_2710),
.B(n_2243),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2825),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2826),
.Y(n_2959)
);

OR2x2_ASAP7_75t_L g2960 ( 
.A(n_2847),
.B(n_2472),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2823),
.B(n_2473),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2793),
.B(n_2475),
.Y(n_2962)
);

INVx4_ASAP7_75t_L g2963 ( 
.A(n_2751),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2794),
.B(n_2476),
.Y(n_2964)
);

CKINVDCx5p33_ASAP7_75t_R g2965 ( 
.A(n_2856),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2845),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2845),
.Y(n_2967)
);

NOR2x1p5_ASAP7_75t_L g2968 ( 
.A(n_2737),
.B(n_2245),
.Y(n_2968)
);

BUFx8_ASAP7_75t_SL g2969 ( 
.A(n_2861),
.Y(n_2969)
);

HB1xp67_ASAP7_75t_L g2970 ( 
.A(n_2776),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2717),
.Y(n_2971)
);

INVx3_ASAP7_75t_L g2972 ( 
.A(n_2815),
.Y(n_2972)
);

BUFx2_ASAP7_75t_L g2973 ( 
.A(n_2742),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2717),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2784),
.B(n_1750),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2721),
.B(n_1758),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2835),
.Y(n_2977)
);

BUFx2_ASAP7_75t_L g2978 ( 
.A(n_2727),
.Y(n_2978)
);

AOI22xp33_ASAP7_75t_SL g2979 ( 
.A1(n_2797),
.A2(n_2006),
.B1(n_2033),
.B2(n_2000),
.Y(n_2979)
);

NAND3x1_ASAP7_75t_L g2980 ( 
.A(n_2764),
.B(n_1598),
.C(n_1596),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2711),
.B(n_2494),
.Y(n_2981)
);

NAND2xp33_ASAP7_75t_SL g2982 ( 
.A(n_2766),
.B(n_2038),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2831),
.Y(n_2983)
);

AND2x6_ASAP7_75t_L g2984 ( 
.A(n_2718),
.B(n_2722),
.Y(n_2984)
);

BUFx10_ASAP7_75t_L g2985 ( 
.A(n_2862),
.Y(n_2985)
);

INVx5_ASAP7_75t_L g2986 ( 
.A(n_2851),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2832),
.B(n_2837),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_2810),
.Y(n_2988)
);

BUFx3_ASAP7_75t_L g2989 ( 
.A(n_2808),
.Y(n_2989)
);

OR2x6_ASAP7_75t_L g2990 ( 
.A(n_2792),
.B(n_2295),
.Y(n_2990)
);

AND2x4_ASAP7_75t_L g2991 ( 
.A(n_2723),
.B(n_2495),
.Y(n_2991)
);

AND2x4_ASAP7_75t_L g2992 ( 
.A(n_2730),
.B(n_2496),
.Y(n_2992)
);

INVx3_ASAP7_75t_L g2993 ( 
.A(n_2747),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2842),
.Y(n_2994)
);

INVx4_ASAP7_75t_L g2995 ( 
.A(n_2743),
.Y(n_2995)
);

INVx3_ASAP7_75t_L g2996 ( 
.A(n_2748),
.Y(n_2996)
);

BUFx6f_ASAP7_75t_L g2997 ( 
.A(n_2754),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2843),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2735),
.B(n_2783),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2812),
.B(n_1599),
.Y(n_3000)
);

INVx5_ASAP7_75t_L g3001 ( 
.A(n_2732),
.Y(n_3001)
);

CKINVDCx5p33_ASAP7_75t_R g3002 ( 
.A(n_2867),
.Y(n_3002)
);

OR2x6_ASAP7_75t_SL g3003 ( 
.A(n_2763),
.B(n_2768),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2757),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2758),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2859),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2864),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2866),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2848),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2850),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2817),
.Y(n_3011)
);

BUFx3_ASAP7_75t_L g3012 ( 
.A(n_2855),
.Y(n_3012)
);

INVx4_ASAP7_75t_L g3013 ( 
.A(n_2712),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2798),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2800),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2779),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2745),
.B(n_1602),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2774),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2738),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2863),
.Y(n_3020)
);

INVx4_ASAP7_75t_SL g3021 ( 
.A(n_2780),
.Y(n_3021)
);

BUFx6f_ASAP7_75t_L g3022 ( 
.A(n_2731),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2740),
.B(n_1603),
.Y(n_3023)
);

INVx3_ASAP7_75t_L g3024 ( 
.A(n_2729),
.Y(n_3024)
);

AND3x4_ASAP7_75t_L g3025 ( 
.A(n_2781),
.B(n_1903),
.C(n_1896),
.Y(n_3025)
);

AND2x4_ASAP7_75t_L g3026 ( 
.A(n_2739),
.B(n_2497),
.Y(n_3026)
);

AND2x6_ASAP7_75t_L g3027 ( 
.A(n_2860),
.B(n_1601),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2865),
.B(n_1848),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2760),
.Y(n_3029)
);

BUFx6f_ASAP7_75t_L g3030 ( 
.A(n_2752),
.Y(n_3030)
);

INVx5_ASAP7_75t_L g3031 ( 
.A(n_2858),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2782),
.B(n_1605),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_SL g3033 ( 
.A(n_2707),
.B(n_2039),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_SL g3034 ( 
.A(n_2796),
.B(n_1612),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2782),
.B(n_1614),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2782),
.B(n_1616),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_2719),
.Y(n_3037)
);

HB1xp67_ASAP7_75t_L g3038 ( 
.A(n_2746),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_2709),
.B(n_2498),
.Y(n_3039)
);

HB1xp67_ASAP7_75t_L g3040 ( 
.A(n_2746),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2767),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2767),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_2796),
.B(n_1617),
.Y(n_3043)
);

INVx4_ASAP7_75t_SL g3044 ( 
.A(n_2799),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2767),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2767),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_2759),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2782),
.B(n_1618),
.Y(n_3048)
);

INVx4_ASAP7_75t_SL g3049 ( 
.A(n_2799),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2715),
.Y(n_3050)
);

INVx5_ASAP7_75t_L g3051 ( 
.A(n_2806),
.Y(n_3051)
);

BUFx3_ASAP7_75t_L g3052 ( 
.A(n_2715),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2834),
.Y(n_3053)
);

AND2x6_ASAP7_75t_L g3054 ( 
.A(n_2830),
.B(n_1606),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2782),
.B(n_1622),
.Y(n_3055)
);

INVx1_ASAP7_75t_SL g3056 ( 
.A(n_2769),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2834),
.Y(n_3057)
);

NAND2xp33_ASAP7_75t_L g3058 ( 
.A(n_2762),
.B(n_2032),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2782),
.B(n_1628),
.Y(n_3059)
);

CKINVDCx5p33_ASAP7_75t_R g3060 ( 
.A(n_2719),
.Y(n_3060)
);

INVx1_ASAP7_75t_SL g3061 ( 
.A(n_2769),
.Y(n_3061)
);

NAND2x1p5_ASAP7_75t_L g3062 ( 
.A(n_2709),
.B(n_2499),
.Y(n_3062)
);

AND2x4_ASAP7_75t_L g3063 ( 
.A(n_2709),
.B(n_1607),
.Y(n_3063)
);

HB1xp67_ASAP7_75t_L g3064 ( 
.A(n_2746),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2767),
.Y(n_3065)
);

BUFx2_ASAP7_75t_L g3066 ( 
.A(n_2746),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2834),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2767),
.Y(n_3068)
);

INVx1_ASAP7_75t_SL g3069 ( 
.A(n_2769),
.Y(n_3069)
);

CKINVDCx5p33_ASAP7_75t_R g3070 ( 
.A(n_2719),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2834),
.Y(n_3071)
);

OAI22xp5_ASAP7_75t_L g3072 ( 
.A1(n_2755),
.A2(n_1695),
.B1(n_1629),
.B2(n_1632),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2767),
.Y(n_3073)
);

AND2x6_ASAP7_75t_L g3074 ( 
.A(n_2830),
.B(n_1608),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2796),
.B(n_1634),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_2767),
.Y(n_3076)
);

AND2x4_ASAP7_75t_L g3077 ( 
.A(n_2709),
.B(n_1611),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2881),
.B(n_1947),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2910),
.B(n_2040),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2894),
.B(n_1635),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2869),
.Y(n_3081)
);

BUFx2_ASAP7_75t_L g3082 ( 
.A(n_2889),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_SL g3083 ( 
.A(n_2986),
.B(n_2048),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_2877),
.B(n_2070),
.Y(n_3084)
);

AOI22xp33_ASAP7_75t_L g3085 ( 
.A1(n_2924),
.A2(n_2093),
.B1(n_2113),
.B2(n_2083),
.Y(n_3085)
);

AND2x4_ASAP7_75t_L g3086 ( 
.A(n_2929),
.B(n_1613),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2937),
.B(n_1637),
.Y(n_3087)
);

O2A1O1Ixp33_ASAP7_75t_L g3088 ( 
.A1(n_2934),
.A2(n_1624),
.B(n_1633),
.C(n_1619),
.Y(n_3088)
);

CKINVDCx5p33_ASAP7_75t_R g3089 ( 
.A(n_2883),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2908),
.B(n_1639),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2950),
.Y(n_3091)
);

BUFx3_ASAP7_75t_L g3092 ( 
.A(n_2988),
.Y(n_3092)
);

NAND2x1p5_ASAP7_75t_L g3093 ( 
.A(n_2972),
.B(n_1636),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2868),
.Y(n_3094)
);

INVx8_ASAP7_75t_L g3095 ( 
.A(n_2946),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2871),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2876),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_3032),
.B(n_1646),
.Y(n_3098)
);

NOR2xp67_ASAP7_75t_L g3099 ( 
.A(n_2986),
.B(n_2057),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_3035),
.B(n_1648),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_3036),
.B(n_1652),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_3041),
.Y(n_3102)
);

INVx2_ASAP7_75t_SL g3103 ( 
.A(n_3066),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_3042),
.Y(n_3104)
);

AND2x4_ASAP7_75t_L g3105 ( 
.A(n_2944),
.B(n_1638),
.Y(n_3105)
);

OAI221xp5_ASAP7_75t_L g3106 ( 
.A1(n_3072),
.A2(n_1651),
.B1(n_1656),
.B2(n_1641),
.C(n_1640),
.Y(n_3106)
);

NAND2xp33_ASAP7_75t_SL g3107 ( 
.A(n_3037),
.B(n_3060),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_3048),
.B(n_1653),
.Y(n_3108)
);

INVxp33_ASAP7_75t_L g3109 ( 
.A(n_3038),
.Y(n_3109)
);

AOI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_2930),
.A2(n_2136),
.B1(n_2155),
.B2(n_2121),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_3055),
.B(n_1654),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_3059),
.B(n_1655),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2885),
.Y(n_3113)
);

INVx2_ASAP7_75t_SL g3114 ( 
.A(n_2873),
.Y(n_3114)
);

NOR2xp67_ASAP7_75t_L g3115 ( 
.A(n_3013),
.B(n_2062),
.Y(n_3115)
);

BUFx5_ASAP7_75t_L g3116 ( 
.A(n_2954),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2918),
.B(n_2252),
.Y(n_3117)
);

INVx2_ASAP7_75t_SL g3118 ( 
.A(n_3039),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_3045),
.Y(n_3119)
);

INVx8_ASAP7_75t_L g3120 ( 
.A(n_2946),
.Y(n_3120)
);

AND2x6_ASAP7_75t_SL g3121 ( 
.A(n_3029),
.B(n_1659),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_3020),
.A2(n_2275),
.B1(n_2276),
.B2(n_2268),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2890),
.Y(n_3123)
);

AND2x4_ASAP7_75t_L g3124 ( 
.A(n_3050),
.B(n_1662),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_SL g3125 ( 
.A(n_3030),
.Y(n_3125)
);

NAND2xp33_ASAP7_75t_L g3126 ( 
.A(n_3070),
.B(n_2069),
.Y(n_3126)
);

AND2x6_ASAP7_75t_L g3127 ( 
.A(n_2971),
.B(n_1663),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_L g3128 ( 
.A1(n_2897),
.A2(n_2283),
.B1(n_2306),
.B2(n_2277),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2967),
.A2(n_1670),
.B(n_1667),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_SL g3130 ( 
.A(n_2998),
.B(n_2313),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2870),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2900),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2987),
.B(n_1660),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2962),
.B(n_1661),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2964),
.B(n_1664),
.Y(n_3135)
);

INVx3_ASAP7_75t_L g3136 ( 
.A(n_2870),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2947),
.B(n_1665),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_2977),
.B(n_1669),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2901),
.B(n_1673),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_SL g3140 ( 
.A(n_2958),
.B(n_1675),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2909),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_2941),
.B(n_2016),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_3046),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2914),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2920),
.Y(n_3145)
);

INVx2_ASAP7_75t_SL g3146 ( 
.A(n_3040),
.Y(n_3146)
);

A2O1A1Ixp33_ASAP7_75t_L g3147 ( 
.A1(n_2974),
.A2(n_1672),
.B(n_1674),
.C(n_1671),
.Y(n_3147)
);

NOR2xp67_ASAP7_75t_L g3148 ( 
.A(n_3051),
.B(n_2081),
.Y(n_3148)
);

BUFx6f_ASAP7_75t_SL g3149 ( 
.A(n_3030),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_SL g3150 ( 
.A1(n_2979),
.A2(n_2097),
.B1(n_2112),
.B2(n_2084),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_2959),
.B(n_1676),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_3053),
.B(n_1678),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_3057),
.B(n_1681),
.Y(n_3153)
);

OAI22xp33_ASAP7_75t_L g3154 ( 
.A1(n_2896),
.A2(n_2120),
.B1(n_2135),
.B2(n_2116),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_2983),
.B(n_1682),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_3065),
.Y(n_3156)
);

NOR2xp33_ASAP7_75t_L g3157 ( 
.A(n_2892),
.B(n_2953),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_SL g3158 ( 
.A(n_2994),
.B(n_1685),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3068),
.Y(n_3159)
);

NOR2xp67_ASAP7_75t_L g3160 ( 
.A(n_3051),
.B(n_2154),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3067),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_3071),
.B(n_1688),
.Y(n_3162)
);

INVx8_ASAP7_75t_L g3163 ( 
.A(n_2984),
.Y(n_3163)
);

NAND2xp33_ASAP7_75t_L g3164 ( 
.A(n_3054),
.B(n_2165),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_3000),
.B(n_1691),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2961),
.B(n_2123),
.Y(n_3166)
);

NOR2xp33_ASAP7_75t_L g3167 ( 
.A(n_2970),
.B(n_1692),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2956),
.B(n_1698),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_3073),
.Y(n_3169)
);

AOI22xp5_ASAP7_75t_L g3170 ( 
.A1(n_2923),
.A2(n_1701),
.B1(n_1708),
.B2(n_1705),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2931),
.B(n_1710),
.Y(n_3171)
);

NOR2xp33_ASAP7_75t_L g3172 ( 
.A(n_3016),
.B(n_1713),
.Y(n_3172)
);

O2A1O1Ixp5_ASAP7_75t_L g3173 ( 
.A1(n_2913),
.A2(n_2042),
.B(n_2047),
.C(n_2003),
.Y(n_3173)
);

AOI22xp33_ASAP7_75t_L g3174 ( 
.A1(n_2933),
.A2(n_2114),
.B1(n_2118),
.B2(n_2111),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2888),
.B(n_1714),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3076),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2887),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2899),
.B(n_1716),
.Y(n_3178)
);

BUFx5_ASAP7_75t_L g3179 ( 
.A(n_2984),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_SL g3180 ( 
.A(n_2893),
.B(n_1717),
.Y(n_3180)
);

AND2x4_ASAP7_75t_L g3181 ( 
.A(n_3052),
.B(n_1686),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_2875),
.B(n_1712),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_3023),
.B(n_1724),
.Y(n_3183)
);

OR2x2_ASAP7_75t_L g3184 ( 
.A(n_2895),
.B(n_2194),
.Y(n_3184)
);

OR2x2_ASAP7_75t_L g3185 ( 
.A(n_2960),
.B(n_2200),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2898),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_SL g3187 ( 
.A(n_3017),
.B(n_1729),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_L g3188 ( 
.A(n_2879),
.B(n_1733),
.Y(n_3188)
);

BUFx6f_ASAP7_75t_L g3189 ( 
.A(n_2872),
.Y(n_3189)
);

AOI22xp33_ASAP7_75t_L g3190 ( 
.A1(n_3074),
.A2(n_2289),
.B1(n_2301),
.B2(n_2278),
.Y(n_3190)
);

AOI22xp33_ASAP7_75t_L g3191 ( 
.A1(n_2904),
.A2(n_2344),
.B1(n_2316),
.B2(n_1725),
.Y(n_3191)
);

AOI22xp5_ASAP7_75t_L g3192 ( 
.A1(n_3058),
.A2(n_1752),
.B1(n_1754),
.B2(n_1749),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2932),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2945),
.Y(n_3194)
);

BUFx3_ASAP7_75t_L g3195 ( 
.A(n_2938),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2917),
.B(n_1759),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_2975),
.B(n_2123),
.Y(n_3197)
);

NAND2x1_ASAP7_75t_L g3198 ( 
.A(n_2940),
.B(n_1719),
.Y(n_3198)
);

AND2x6_ASAP7_75t_L g3199 ( 
.A(n_3022),
.B(n_1726),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2955),
.A2(n_1765),
.B1(n_1767),
.B2(n_1762),
.Y(n_3200)
);

NAND2xp33_ASAP7_75t_L g3201 ( 
.A(n_2999),
.B(n_2202),
.Y(n_3201)
);

CKINVDCx5p33_ASAP7_75t_R g3202 ( 
.A(n_2969),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2921),
.B(n_1771),
.Y(n_3203)
);

BUFx8_ASAP7_75t_L g3204 ( 
.A(n_2978),
.Y(n_3204)
);

NAND3xp33_ASAP7_75t_L g3205 ( 
.A(n_2982),
.B(n_1773),
.C(n_1772),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2942),
.B(n_1775),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2949),
.B(n_1777),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2976),
.B(n_2175),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_2891),
.B(n_1780),
.Y(n_3209)
);

AOI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_3034),
.A2(n_1786),
.B1(n_1787),
.B2(n_1785),
.Y(n_3210)
);

OAI22xp33_ASAP7_75t_L g3211 ( 
.A1(n_3033),
.A2(n_2207),
.B1(n_2234),
.B2(n_2206),
.Y(n_3211)
);

NOR2x1p5_ASAP7_75t_L g3212 ( 
.A(n_2880),
.B(n_2238),
.Y(n_3212)
);

NAND3xp33_ASAP7_75t_L g3213 ( 
.A(n_3043),
.B(n_1790),
.C(n_1789),
.Y(n_3213)
);

CKINVDCx5p33_ASAP7_75t_R g3214 ( 
.A(n_2965),
.Y(n_3214)
);

AO221x1_ASAP7_75t_L g3215 ( 
.A1(n_2874),
.A2(n_1738),
.B1(n_1739),
.B2(n_1730),
.C(n_1727),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2878),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_L g3217 ( 
.A(n_3056),
.B(n_1795),
.Y(n_3217)
);

INVxp67_ASAP7_75t_L g3218 ( 
.A(n_3064),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_2919),
.A2(n_1742),
.B(n_1741),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2886),
.Y(n_3220)
);

NAND3xp33_ASAP7_75t_L g3221 ( 
.A(n_3075),
.B(n_1807),
.C(n_1797),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_2995),
.B(n_1808),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2872),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_2927),
.B(n_1809),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2903),
.Y(n_3225)
);

INVx3_ASAP7_75t_L g3226 ( 
.A(n_2882),
.Y(n_3226)
);

AOI22xp33_ASAP7_75t_L g3227 ( 
.A1(n_2884),
.A2(n_1770),
.B1(n_1774),
.B2(n_1769),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_3061),
.B(n_1819),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_3069),
.B(n_1823),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2952),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2905),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2951),
.Y(n_3232)
);

A2O1A1Ixp33_ASAP7_75t_L g3233 ( 
.A1(n_2907),
.A2(n_1788),
.B(n_1792),
.C(n_1784),
.Y(n_3233)
);

OR2x6_ASAP7_75t_L g3234 ( 
.A(n_2963),
.B(n_1794),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_SL g3235 ( 
.A(n_3019),
.B(n_1831),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_2882),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2981),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2916),
.B(n_1837),
.Y(n_3238)
);

NOR2xp33_ASAP7_75t_L g3239 ( 
.A(n_2926),
.B(n_1841),
.Y(n_3239)
);

AOI22xp33_ASAP7_75t_L g3240 ( 
.A1(n_3021),
.A2(n_1800),
.B1(n_1801),
.B2(n_1798),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2991),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3028),
.B(n_2208),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_2902),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2992),
.Y(n_3244)
);

OR2x2_ASAP7_75t_L g3245 ( 
.A(n_3011),
.B(n_3009),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_3015),
.B(n_1844),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2993),
.B(n_1851),
.Y(n_3247)
);

INVx2_ASAP7_75t_SL g3248 ( 
.A(n_3026),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_2928),
.B(n_1856),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2996),
.B(n_1858),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3004),
.Y(n_3251)
);

BUFx2_ASAP7_75t_L g3252 ( 
.A(n_3010),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3006),
.Y(n_3253)
);

NOR3xp33_ASAP7_75t_L g3254 ( 
.A(n_3018),
.B(n_1865),
.C(n_1861),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3007),
.Y(n_3255)
);

AND2x6_ASAP7_75t_SL g3256 ( 
.A(n_3014),
.B(n_1803),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_3025),
.A2(n_1814),
.B1(n_1827),
.B2(n_1812),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3008),
.B(n_1866),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2943),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_2911),
.B(n_1869),
.Y(n_3260)
);

BUFx6f_ASAP7_75t_L g3261 ( 
.A(n_2902),
.Y(n_3261)
);

INVx2_ASAP7_75t_SL g3262 ( 
.A(n_2912),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2915),
.B(n_1875),
.Y(n_3263)
);

NOR2xp67_ASAP7_75t_L g3264 ( 
.A(n_3031),
.B(n_2250),
.Y(n_3264)
);

INVx3_ASAP7_75t_L g3265 ( 
.A(n_2935),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2997),
.B(n_1879),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_3005),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3005),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3047),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3047),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3063),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_3077),
.B(n_1880),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_2936),
.A2(n_1839),
.B(n_1829),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2957),
.B(n_1882),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3062),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2957),
.B(n_1883),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_2906),
.B(n_2208),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_SL g3278 ( 
.A(n_3001),
.B(n_1887),
.Y(n_3278)
);

INVx5_ASAP7_75t_L g3279 ( 
.A(n_3027),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3044),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3049),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2939),
.B(n_1889),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_3024),
.B(n_1891),
.Y(n_3283)
);

INVx8_ASAP7_75t_L g3284 ( 
.A(n_3031),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_SL g3285 ( 
.A(n_3001),
.B(n_1892),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_2973),
.A2(n_1901),
.B1(n_1904),
.B2(n_1894),
.Y(n_3286)
);

OR2x6_ASAP7_75t_L g3287 ( 
.A(n_2989),
.B(n_1842),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2990),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2948),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3027),
.B(n_1905),
.Y(n_3290)
);

INVx2_ASAP7_75t_SL g3291 ( 
.A(n_3012),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2980),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2968),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_SL g3294 ( 
.A(n_3002),
.B(n_1908),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_SL g3295 ( 
.A(n_2922),
.B(n_1911),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2925),
.B(n_1912),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2985),
.B(n_1913),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3003),
.B(n_1914),
.Y(n_3298)
);

INVx2_ASAP7_75t_SL g3299 ( 
.A(n_2881),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_2881),
.B(n_2351),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2894),
.B(n_1923),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_2894),
.A2(n_1852),
.B1(n_1854),
.B2(n_1847),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_2986),
.B(n_1925),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_2894),
.B(n_1928),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_SL g3305 ( 
.A(n_2986),
.B(n_1930),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2894),
.B(n_1932),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2869),
.Y(n_3307)
);

NAND3xp33_ASAP7_75t_L g3308 ( 
.A(n_2894),
.B(n_1937),
.C(n_1936),
.Y(n_3308)
);

AOI22xp5_ASAP7_75t_L g3309 ( 
.A1(n_2894),
.A2(n_1940),
.B1(n_1941),
.B2(n_1938),
.Y(n_3309)
);

AOI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_2894),
.A2(n_1946),
.B1(n_1949),
.B2(n_1945),
.Y(n_3310)
);

NOR2xp67_ASAP7_75t_SL g3311 ( 
.A(n_2986),
.B(n_1857),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_2910),
.B(n_1952),
.Y(n_3312)
);

BUFx3_ASAP7_75t_L g3313 ( 
.A(n_2988),
.Y(n_3313)
);

INVxp67_ASAP7_75t_SL g3314 ( 
.A(n_2950),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2869),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_SL g3316 ( 
.A(n_2986),
.B(n_1957),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2894),
.B(n_1962),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2894),
.B(n_1963),
.Y(n_3318)
);

INVx2_ASAP7_75t_SL g3319 ( 
.A(n_2881),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_2966),
.A2(n_1862),
.B(n_1860),
.Y(n_3320)
);

A2O1A1Ixp33_ASAP7_75t_L g3321 ( 
.A1(n_2894),
.A2(n_1876),
.B(n_1878),
.C(n_1867),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2894),
.B(n_1968),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_2910),
.B(n_1969),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2986),
.B(n_1973),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_2950),
.Y(n_3325)
);

AOI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_2894),
.A2(n_1977),
.B1(n_1979),
.B2(n_1975),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2950),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_2869),
.Y(n_3328)
);

NAND2xp33_ASAP7_75t_L g3329 ( 
.A(n_2883),
.B(n_2262),
.Y(n_3329)
);

INVxp67_ASAP7_75t_L g3330 ( 
.A(n_2881),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2894),
.B(n_1991),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2894),
.B(n_1995),
.Y(n_3332)
);

INVxp67_ASAP7_75t_L g3333 ( 
.A(n_2881),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_SL g3334 ( 
.A(n_2986),
.B(n_1996),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_2910),
.B(n_1997),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3312),
.B(n_1998),
.Y(n_3336)
);

INVx3_ASAP7_75t_L g3337 ( 
.A(n_3092),
.Y(n_3337)
);

OAI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3314),
.A2(n_2002),
.B1(n_2005),
.B2(n_2001),
.Y(n_3338)
);

BUFx6f_ASAP7_75t_L g3339 ( 
.A(n_3131),
.Y(n_3339)
);

BUFx8_ASAP7_75t_L g3340 ( 
.A(n_3125),
.Y(n_3340)
);

BUFx6f_ASAP7_75t_L g3341 ( 
.A(n_3131),
.Y(n_3341)
);

OAI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_3323),
.A2(n_3335),
.B(n_3325),
.Y(n_3342)
);

BUFx2_ASAP7_75t_L g3343 ( 
.A(n_3082),
.Y(n_3343)
);

O2A1O1Ixp33_ASAP7_75t_L g3344 ( 
.A1(n_3079),
.A2(n_1886),
.B(n_1890),
.C(n_1885),
.Y(n_3344)
);

BUFx6f_ASAP7_75t_L g3345 ( 
.A(n_3189),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_3157),
.B(n_2008),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3080),
.B(n_2009),
.Y(n_3347)
);

INVx4_ASAP7_75t_L g3348 ( 
.A(n_3313),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3301),
.B(n_2010),
.Y(n_3349)
);

OA21x2_ASAP7_75t_L g3350 ( 
.A1(n_3147),
.A2(n_1898),
.B(n_1895),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_SL g3351 ( 
.A(n_3299),
.B(n_2011),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3304),
.B(n_2012),
.Y(n_3352)
);

BUFx2_ASAP7_75t_SL g3353 ( 
.A(n_3149),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3081),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3306),
.B(n_2013),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3097),
.Y(n_3356)
);

BUFx12f_ASAP7_75t_L g3357 ( 
.A(n_3204),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_3091),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_3319),
.B(n_2020),
.Y(n_3359)
);

OAI22xp5_ASAP7_75t_L g3360 ( 
.A1(n_3317),
.A2(n_2023),
.B1(n_2024),
.B2(n_2022),
.Y(n_3360)
);

O2A1O1Ixp33_ASAP7_75t_L g3361 ( 
.A1(n_3318),
.A2(n_1915),
.B(n_1922),
.C(n_1909),
.Y(n_3361)
);

AOI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3098),
.A2(n_1929),
.B(n_1927),
.Y(n_3362)
);

AO21x1_ASAP7_75t_L g3363 ( 
.A1(n_3322),
.A2(n_1935),
.B(n_1933),
.Y(n_3363)
);

OAI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3327),
.A2(n_1943),
.B(n_1939),
.Y(n_3364)
);

AOI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_3100),
.A2(n_1954),
.B(n_1950),
.Y(n_3365)
);

CKINVDCx5p33_ASAP7_75t_R g3366 ( 
.A(n_3089),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3101),
.A2(n_1958),
.B(n_1955),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3331),
.B(n_3332),
.Y(n_3368)
);

BUFx6f_ASAP7_75t_L g3369 ( 
.A(n_3189),
.Y(n_3369)
);

AOI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_3084),
.A2(n_2028),
.B1(n_2029),
.B2(n_2025),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3094),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_3142),
.B(n_3166),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3108),
.A2(n_1970),
.B(n_1966),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3133),
.B(n_2034),
.Y(n_3374)
);

O2A1O1Ixp5_ASAP7_75t_L g3375 ( 
.A1(n_3111),
.A2(n_1986),
.B(n_1989),
.C(n_1983),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3078),
.B(n_3300),
.Y(n_3376)
);

NOR2x1_ASAP7_75t_L g3377 ( 
.A(n_3213),
.B(n_1990),
.Y(n_3377)
);

OR2x6_ASAP7_75t_L g3378 ( 
.A(n_3284),
.B(n_1992),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_3330),
.B(n_3333),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3112),
.A2(n_1994),
.B(n_1993),
.Y(n_3380)
);

OAI22xp5_ASAP7_75t_L g3381 ( 
.A1(n_3113),
.A2(n_2044),
.B1(n_2046),
.B2(n_2043),
.Y(n_3381)
);

BUFx8_ASAP7_75t_L g3382 ( 
.A(n_3103),
.Y(n_3382)
);

NOR2xp67_ASAP7_75t_L g3383 ( 
.A(n_3214),
.B(n_2323),
.Y(n_3383)
);

OAI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3123),
.A2(n_2051),
.B1(n_2053),
.B2(n_2050),
.Y(n_3384)
);

INVx3_ASAP7_75t_L g3385 ( 
.A(n_3223),
.Y(n_3385)
);

NAND2xp33_ASAP7_75t_L g3386 ( 
.A(n_3179),
.B(n_3116),
.Y(n_3386)
);

A2O1A1Ixp33_ASAP7_75t_L g3387 ( 
.A1(n_3249),
.A2(n_2019),
.B(n_2021),
.C(n_2018),
.Y(n_3387)
);

AOI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_3165),
.A2(n_2060),
.B1(n_2063),
.B2(n_2056),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3197),
.B(n_2329),
.Y(n_3389)
);

AOI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_3127),
.A2(n_2037),
.B1(n_2041),
.B2(n_2031),
.Y(n_3390)
);

O2A1O1Ixp33_ASAP7_75t_L g3391 ( 
.A1(n_3106),
.A2(n_2054),
.B(n_2055),
.C(n_2052),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3146),
.B(n_2065),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3137),
.B(n_2066),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3087),
.A2(n_2068),
.B(n_2058),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_3208),
.B(n_2330),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3132),
.B(n_2067),
.Y(n_3396)
);

A2O1A1Ixp33_ASAP7_75t_L g3397 ( 
.A1(n_3172),
.A2(n_2073),
.B(n_2076),
.C(n_2074),
.Y(n_3397)
);

AND3x4_ASAP7_75t_L g3398 ( 
.A(n_3264),
.B(n_3254),
.C(n_3195),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_L g3399 ( 
.A(n_3110),
.B(n_2071),
.Y(n_3399)
);

NOR2xp67_ASAP7_75t_L g3400 ( 
.A(n_3279),
.B(n_2331),
.Y(n_3400)
);

AOI21x1_ASAP7_75t_L g3401 ( 
.A1(n_3193),
.A2(n_2119),
.B(n_2115),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3141),
.B(n_2075),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3144),
.B(n_2077),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_3109),
.B(n_2079),
.Y(n_3404)
);

INVx1_ASAP7_75t_SL g3405 ( 
.A(n_3245),
.Y(n_3405)
);

A2O1A1Ixp33_ASAP7_75t_L g3406 ( 
.A1(n_3308),
.A2(n_2128),
.B(n_2131),
.C(n_2125),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3145),
.B(n_2080),
.Y(n_3407)
);

INVx2_ASAP7_75t_SL g3408 ( 
.A(n_3124),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3161),
.B(n_2087),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3187),
.A2(n_2145),
.B(n_2144),
.Y(n_3410)
);

AOI21x1_ASAP7_75t_L g3411 ( 
.A1(n_3194),
.A2(n_2149),
.B(n_2147),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3307),
.B(n_3315),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3328),
.B(n_2088),
.Y(n_3413)
);

NAND2xp33_ASAP7_75t_L g3414 ( 
.A(n_3179),
.B(n_2342),
.Y(n_3414)
);

AOI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_3171),
.A2(n_2151),
.B(n_2150),
.Y(n_3415)
);

BUFx6f_ASAP7_75t_L g3416 ( 
.A(n_3223),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3096),
.Y(n_3417)
);

INVx6_ASAP7_75t_L g3418 ( 
.A(n_3095),
.Y(n_3418)
);

INVx3_ASAP7_75t_L g3419 ( 
.A(n_3261),
.Y(n_3419)
);

AOI33xp33_ASAP7_75t_L g3420 ( 
.A1(n_3257),
.A2(n_2184),
.A3(n_2178),
.B1(n_2187),
.B2(n_2182),
.B3(n_2170),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3283),
.A2(n_2091),
.B1(n_2092),
.B2(n_2090),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_3134),
.A2(n_2192),
.B(n_2189),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3102),
.Y(n_3423)
);

AOI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_3135),
.A2(n_3119),
.B(n_3104),
.Y(n_3424)
);

INVx4_ASAP7_75t_L g3425 ( 
.A(n_3095),
.Y(n_3425)
);

HB1xp67_ASAP7_75t_L g3426 ( 
.A(n_3218),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3143),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_3122),
.B(n_2095),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3090),
.B(n_2096),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_3127),
.A2(n_2199),
.B1(n_2201),
.B2(n_2197),
.Y(n_3430)
);

INVx3_ASAP7_75t_L g3431 ( 
.A(n_3261),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3242),
.B(n_3175),
.Y(n_3432)
);

NOR2xp33_ASAP7_75t_SL g3433 ( 
.A(n_3202),
.B(n_2098),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_SL g3434 ( 
.A(n_3284),
.B(n_3120),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_L g3435 ( 
.A(n_3188),
.B(n_2100),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3178),
.B(n_2104),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3127),
.B(n_2105),
.Y(n_3437)
);

NOR2xp67_ASAP7_75t_L g3438 ( 
.A(n_3221),
.B(n_2106),
.Y(n_3438)
);

OAI21xp33_ASAP7_75t_L g3439 ( 
.A1(n_3085),
.A2(n_3310),
.B(n_3309),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3156),
.Y(n_3440)
);

AOI21xp33_ASAP7_75t_L g3441 ( 
.A1(n_3168),
.A2(n_2117),
.B(n_2109),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3251),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3217),
.B(n_2124),
.Y(n_3443)
);

OAI21xp33_ASAP7_75t_L g3444 ( 
.A1(n_3326),
.A2(n_2127),
.B(n_2126),
.Y(n_3444)
);

INVx4_ASAP7_75t_L g3445 ( 
.A(n_3120),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3159),
.B(n_2129),
.Y(n_3446)
);

A2O1A1Ixp33_ASAP7_75t_L g3447 ( 
.A1(n_3167),
.A2(n_2218),
.B(n_2219),
.C(n_2213),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_3169),
.A2(n_2240),
.B(n_2222),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3107),
.B(n_3116),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3176),
.Y(n_3450)
);

BUFx6f_ASAP7_75t_L g3451 ( 
.A(n_3262),
.Y(n_3451)
);

AO21x1_ASAP7_75t_L g3452 ( 
.A1(n_3129),
.A2(n_2247),
.B(n_2241),
.Y(n_3452)
);

O2A1O1Ixp5_ASAP7_75t_L g3453 ( 
.A1(n_3183),
.A2(n_2263),
.B(n_2265),
.C(n_2261),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_3116),
.B(n_2132),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3177),
.Y(n_3455)
);

INVx2_ASAP7_75t_SL g3456 ( 
.A(n_3181),
.Y(n_3456)
);

O2A1O1Ixp33_ASAP7_75t_L g3457 ( 
.A1(n_3321),
.A2(n_2269),
.B(n_2273),
.C(n_2267),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3255),
.Y(n_3458)
);

NOR2x1_ASAP7_75t_L g3459 ( 
.A(n_3205),
.B(n_2279),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3186),
.B(n_2133),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_3280),
.B(n_2282),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3230),
.Y(n_3462)
);

AND2x2_ASAP7_75t_SL g3463 ( 
.A(n_3128),
.B(n_2285),
.Y(n_3463)
);

OAI321xp33_ASAP7_75t_L g3464 ( 
.A1(n_3150),
.A2(n_2307),
.A3(n_2294),
.B1(n_2315),
.B2(n_2304),
.C(n_2288),
.Y(n_3464)
);

OAI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3139),
.A2(n_2318),
.B(n_2317),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3253),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3216),
.B(n_2138),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3184),
.B(n_2139),
.Y(n_3468)
);

A2O1A1Ixp33_ASAP7_75t_L g3469 ( 
.A1(n_3239),
.A2(n_2320),
.B(n_2321),
.C(n_2319),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3259),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3130),
.B(n_2140),
.Y(n_3471)
);

AO21x1_ASAP7_75t_L g3472 ( 
.A1(n_3320),
.A2(n_2343),
.B(n_2341),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3117),
.B(n_2142),
.Y(n_3473)
);

NOR2xp33_ASAP7_75t_L g3474 ( 
.A(n_3252),
.B(n_2148),
.Y(n_3474)
);

INVx1_ASAP7_75t_SL g3475 ( 
.A(n_3086),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_3206),
.A2(n_2350),
.B(n_2348),
.Y(n_3476)
);

AOI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3201),
.A2(n_2153),
.B1(n_2156),
.B2(n_2152),
.Y(n_3477)
);

AOI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_3207),
.A2(n_2360),
.B(n_2356),
.Y(n_3478)
);

OR2x6_ASAP7_75t_L g3479 ( 
.A(n_3163),
.B(n_340),
.Y(n_3479)
);

NAND2x1p5_ASAP7_75t_L g3480 ( 
.A(n_3136),
.B(n_340),
.Y(n_3480)
);

OAI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_3152),
.A2(n_2158),
.B(n_2157),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_3247),
.A2(n_2160),
.B(n_2159),
.Y(n_3482)
);

AO21x1_ASAP7_75t_L g3483 ( 
.A1(n_3180),
.A2(n_342),
.B(n_341),
.Y(n_3483)
);

AOI22xp5_ASAP7_75t_L g3484 ( 
.A1(n_3140),
.A2(n_2163),
.B1(n_2167),
.B2(n_2161),
.Y(n_3484)
);

AOI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_3250),
.A2(n_2169),
.B(n_2168),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3198),
.Y(n_3486)
);

OAI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3153),
.A2(n_2172),
.B(n_2171),
.Y(n_3487)
);

OAI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_3162),
.A2(n_2174),
.B(n_2173),
.Y(n_3488)
);

AND2x4_ASAP7_75t_L g3489 ( 
.A(n_3281),
.B(n_2177),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_3266),
.A2(n_2181),
.B(n_2179),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3173),
.Y(n_3491)
);

AO21x1_ASAP7_75t_L g3492 ( 
.A1(n_3088),
.A2(n_342),
.B(n_341),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3267),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3268),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3196),
.B(n_2183),
.Y(n_3495)
);

HB1xp67_ASAP7_75t_L g3496 ( 
.A(n_3248),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_3138),
.A2(n_2188),
.B(n_2186),
.Y(n_3497)
);

AOI21x1_ASAP7_75t_L g3498 ( 
.A1(n_3203),
.A2(n_344),
.B(n_343),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3260),
.A2(n_2205),
.B(n_2204),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3269),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3232),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3185),
.B(n_2209),
.Y(n_3502)
);

INVx1_ASAP7_75t_SL g3503 ( 
.A(n_3105),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3220),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3263),
.A2(n_2211),
.B(n_2210),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3270),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3258),
.B(n_2212),
.Y(n_3507)
);

NOR2xp67_ASAP7_75t_L g3508 ( 
.A(n_3291),
.B(n_2214),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3246),
.A2(n_2217),
.B(n_2215),
.Y(n_3509)
);

AOI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_3151),
.A2(n_2223),
.B(n_2221),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3225),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3155),
.A2(n_2226),
.B(n_2225),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_3158),
.A2(n_2230),
.B(n_2229),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_3093),
.B(n_2232),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3231),
.Y(n_3515)
);

BUFx12f_ASAP7_75t_L g3516 ( 
.A(n_3199),
.Y(n_3516)
);

AOI21x1_ASAP7_75t_L g3517 ( 
.A1(n_3235),
.A2(n_346),
.B(n_345),
.Y(n_3517)
);

O2A1O1Ixp33_ASAP7_75t_SL g3518 ( 
.A1(n_3233),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_3518)
);

BUFx6f_ASAP7_75t_L g3519 ( 
.A(n_3226),
.Y(n_3519)
);

AOI21xp33_ASAP7_75t_L g3520 ( 
.A1(n_3238),
.A2(n_2235),
.B(n_2233),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3240),
.B(n_2236),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3154),
.B(n_2237),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_3083),
.B(n_2239),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3182),
.B(n_2244),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3118),
.A2(n_2248),
.B(n_2246),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3114),
.A2(n_2251),
.B(n_2249),
.Y(n_3526)
);

A2O1A1Ixp33_ASAP7_75t_L g3527 ( 
.A1(n_3192),
.A2(n_2255),
.B(n_2256),
.C(n_2254),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3282),
.A2(n_2259),
.B(n_2258),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3227),
.B(n_2260),
.Y(n_3529)
);

AND2x6_ASAP7_75t_SL g3530 ( 
.A(n_3298),
.B(n_3287),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3302),
.B(n_2264),
.Y(n_3531)
);

AOI21x1_ASAP7_75t_L g3532 ( 
.A1(n_3219),
.A2(n_348),
.B(n_347),
.Y(n_3532)
);

NAND3xp33_ASAP7_75t_L g3533 ( 
.A(n_3126),
.B(n_2270),
.C(n_2266),
.Y(n_3533)
);

OAI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3228),
.A2(n_3229),
.B(n_3272),
.Y(n_3534)
);

CKINVDCx20_ASAP7_75t_R g3535 ( 
.A(n_3294),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3237),
.A2(n_2272),
.B(n_2271),
.Y(n_3536)
);

OAI21xp5_ASAP7_75t_L g3537 ( 
.A1(n_3274),
.A2(n_3276),
.B(n_3273),
.Y(n_3537)
);

AOI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_3241),
.A2(n_3244),
.B(n_3275),
.Y(n_3538)
);

OAI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3210),
.A2(n_2281),
.B(n_2280),
.Y(n_3539)
);

AOI21xp5_ASAP7_75t_L g3540 ( 
.A1(n_3222),
.A2(n_2286),
.B(n_2284),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3236),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_3099),
.B(n_2287),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3115),
.B(n_2290),
.Y(n_3543)
);

AOI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3163),
.A2(n_2292),
.B(n_2291),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3243),
.Y(n_3545)
);

INVx2_ASAP7_75t_SL g3546 ( 
.A(n_3271),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3265),
.Y(n_3547)
);

BUFx6f_ASAP7_75t_L g3548 ( 
.A(n_3339),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_SL g3549 ( 
.A(n_3342),
.B(n_3292),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3386),
.A2(n_3290),
.B(n_3164),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3368),
.B(n_3329),
.Y(n_3551)
);

INVxp33_ASAP7_75t_SL g3552 ( 
.A(n_3366),
.Y(n_3552)
);

AND2x4_ASAP7_75t_L g3553 ( 
.A(n_3337),
.B(n_3293),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3432),
.B(n_3211),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_3405),
.B(n_3289),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3537),
.A2(n_3297),
.B(n_3296),
.Y(n_3556)
);

BUFx12f_ASAP7_75t_L g3557 ( 
.A(n_3340),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3356),
.Y(n_3558)
);

BUFx3_ASAP7_75t_L g3559 ( 
.A(n_3418),
.Y(n_3559)
);

O2A1O1Ixp5_ASAP7_75t_SL g3560 ( 
.A1(n_3491),
.A2(n_3303),
.B(n_3316),
.C(n_3305),
.Y(n_3560)
);

NOR2xp33_ASAP7_75t_L g3561 ( 
.A(n_3346),
.B(n_3209),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3435),
.B(n_3224),
.Y(n_3562)
);

INVxp67_ASAP7_75t_L g3563 ( 
.A(n_3343),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_3424),
.A2(n_3334),
.B(n_3324),
.Y(n_3564)
);

NOR2x1_ASAP7_75t_L g3565 ( 
.A(n_3353),
.B(n_3212),
.Y(n_3565)
);

OAI22xp5_ASAP7_75t_L g3566 ( 
.A1(n_3412),
.A2(n_3160),
.B1(n_3148),
.B2(n_3286),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_SL g3567 ( 
.A(n_3372),
.B(n_3277),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_3449),
.A2(n_3285),
.B(n_3278),
.Y(n_3568)
);

OAI22xp5_ASAP7_75t_SL g3569 ( 
.A1(n_3399),
.A2(n_3535),
.B1(n_3428),
.B2(n_3463),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3376),
.B(n_3288),
.Y(n_3570)
);

HB1xp67_ASAP7_75t_L g3571 ( 
.A(n_3426),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_SL g3572 ( 
.A(n_3474),
.B(n_3170),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_3454),
.A2(n_3295),
.B(n_3234),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3442),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3458),
.Y(n_3575)
);

O2A1O1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_3336),
.A2(n_3200),
.B(n_3234),
.C(n_3191),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3374),
.B(n_3215),
.Y(n_3577)
);

AOI22xp33_ASAP7_75t_L g3578 ( 
.A1(n_3471),
.A2(n_3174),
.B1(n_3199),
.B2(n_3190),
.Y(n_3578)
);

NOR2x1_ASAP7_75t_L g3579 ( 
.A(n_3425),
.B(n_3199),
.Y(n_3579)
);

HB1xp67_ASAP7_75t_L g3580 ( 
.A(n_3341),
.Y(n_3580)
);

OAI22xp5_ASAP7_75t_L g3581 ( 
.A1(n_3347),
.A2(n_2296),
.B1(n_2297),
.B2(n_2293),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_3443),
.B(n_2298),
.Y(n_3582)
);

NAND2xp33_ASAP7_75t_SL g3583 ( 
.A(n_3398),
.B(n_3311),
.Y(n_3583)
);

O2A1O1Ixp33_ASAP7_75t_L g3584 ( 
.A1(n_3465),
.A2(n_3344),
.B(n_3522),
.C(n_3387),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3462),
.Y(n_3585)
);

INVx5_ASAP7_75t_L g3586 ( 
.A(n_3418),
.Y(n_3586)
);

OAI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3349),
.A2(n_2303),
.B1(n_2305),
.B2(n_2300),
.Y(n_3587)
);

AND2x4_ASAP7_75t_L g3588 ( 
.A(n_3408),
.B(n_2308),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3534),
.A2(n_3355),
.B(n_3352),
.Y(n_3589)
);

AO32x1_ASAP7_75t_L g3590 ( 
.A1(n_3360),
.A2(n_3121),
.A3(n_3256),
.B1(n_3),
.B2(n_1),
.Y(n_3590)
);

BUFx6f_ASAP7_75t_L g3591 ( 
.A(n_3341),
.Y(n_3591)
);

INVxp67_ASAP7_75t_L g3592 ( 
.A(n_3496),
.Y(n_3592)
);

O2A1O1Ixp33_ASAP7_75t_SL g3593 ( 
.A1(n_3527),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3414),
.A2(n_3393),
.B(n_3495),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3436),
.B(n_2324),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_3382),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3429),
.A2(n_2326),
.B(n_2325),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3507),
.B(n_2332),
.Y(n_3598)
);

A2O1A1Ixp33_ASAP7_75t_L g3599 ( 
.A1(n_3473),
.A2(n_3441),
.B(n_3523),
.C(n_3361),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_3538),
.A2(n_2335),
.B(n_2333),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_SL g3601 ( 
.A(n_3546),
.B(n_2337),
.Y(n_3601)
);

AOI22xp5_ASAP7_75t_L g3602 ( 
.A1(n_3383),
.A2(n_2339),
.B1(n_2340),
.B2(n_2338),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_3345),
.Y(n_3603)
);

HB1xp67_ASAP7_75t_L g3604 ( 
.A(n_3369),
.Y(n_3604)
);

AND2x4_ASAP7_75t_L g3605 ( 
.A(n_3456),
.B(n_2345),
.Y(n_3605)
);

NOR2x1_ASAP7_75t_L g3606 ( 
.A(n_3445),
.B(n_2346),
.Y(n_3606)
);

OAI22xp5_ASAP7_75t_SL g3607 ( 
.A1(n_3479),
.A2(n_2349),
.B1(n_2352),
.B2(n_2347),
.Y(n_3607)
);

A2O1A1Ixp33_ASAP7_75t_L g3608 ( 
.A1(n_3539),
.A2(n_2354),
.B(n_2355),
.C(n_2353),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_3379),
.B(n_2358),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3420),
.B(n_4),
.Y(n_3610)
);

OAI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3358),
.A2(n_351),
.B1(n_352),
.B2(n_349),
.Y(n_3611)
);

BUFx6f_ASAP7_75t_L g3612 ( 
.A(n_3416),
.Y(n_3612)
);

NOR2xp33_ASAP7_75t_R g3613 ( 
.A(n_3434),
.B(n_353),
.Y(n_3613)
);

BUFx3_ASAP7_75t_L g3614 ( 
.A(n_3416),
.Y(n_3614)
);

NAND3xp33_ASAP7_75t_L g3615 ( 
.A(n_3388),
.B(n_4),
.C(n_5),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_R g3616 ( 
.A(n_3385),
.B(n_354),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_L g3617 ( 
.A(n_3404),
.B(n_354),
.Y(n_3617)
);

OAI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3466),
.A2(n_358),
.B1(n_359),
.B2(n_355),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_3475),
.B(n_359),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3468),
.B(n_5),
.Y(n_3620)
);

NOR3xp33_ASAP7_75t_L g3621 ( 
.A(n_3464),
.B(n_3520),
.C(n_3543),
.Y(n_3621)
);

BUFx6f_ASAP7_75t_L g3622 ( 
.A(n_3451),
.Y(n_3622)
);

O2A1O1Ixp33_ASAP7_75t_L g3623 ( 
.A1(n_3397),
.A2(n_361),
.B(n_362),
.C(n_360),
.Y(n_3623)
);

O2A1O1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3447),
.A2(n_361),
.B(n_362),
.C(n_360),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_L g3625 ( 
.A(n_3503),
.B(n_363),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_SL g3626 ( 
.A(n_3514),
.B(n_365),
.Y(n_3626)
);

OAI22xp5_ASAP7_75t_L g3627 ( 
.A1(n_3493),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_3627)
);

AO21x2_ASAP7_75t_L g3628 ( 
.A1(n_3401),
.A2(n_7),
.B(n_8),
.Y(n_3628)
);

AOI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_3351),
.A2(n_368),
.B(n_366),
.Y(n_3629)
);

OAI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_3494),
.A2(n_370),
.B1(n_372),
.B2(n_369),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3389),
.B(n_9),
.Y(n_3631)
);

BUFx8_ASAP7_75t_SL g3632 ( 
.A(n_3357),
.Y(n_3632)
);

INVx3_ASAP7_75t_L g3633 ( 
.A(n_3519),
.Y(n_3633)
);

NOR2xp33_ASAP7_75t_R g3634 ( 
.A(n_3419),
.B(n_369),
.Y(n_3634)
);

O2A1O1Ixp33_ASAP7_75t_L g3635 ( 
.A1(n_3469),
.A2(n_374),
.B(n_375),
.C(n_373),
.Y(n_3635)
);

BUFx12f_ASAP7_75t_L g3636 ( 
.A(n_3516),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3371),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_SL g3638 ( 
.A1(n_3364),
.A2(n_374),
.B(n_373),
.Y(n_3638)
);

OAI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_3417),
.A2(n_378),
.B1(n_379),
.B2(n_376),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3423),
.Y(n_3640)
);

HB1xp67_ASAP7_75t_L g3641 ( 
.A(n_3431),
.Y(n_3641)
);

NOR2xp33_ASAP7_75t_L g3642 ( 
.A(n_3502),
.B(n_381),
.Y(n_3642)
);

NOR2xp33_ASAP7_75t_L g3643 ( 
.A(n_3444),
.B(n_383),
.Y(n_3643)
);

NAND2x1p5_ASAP7_75t_L g3644 ( 
.A(n_3519),
.B(n_383),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3395),
.B(n_9),
.Y(n_3645)
);

INVx5_ASAP7_75t_L g3646 ( 
.A(n_3378),
.Y(n_3646)
);

NAND2x1p5_ASAP7_75t_L g3647 ( 
.A(n_3541),
.B(n_384),
.Y(n_3647)
);

AO32x2_ASAP7_75t_L g3648 ( 
.A1(n_3381),
.A2(n_12),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3427),
.Y(n_3649)
);

BUFx3_ASAP7_75t_L g3650 ( 
.A(n_3545),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_SL g3651 ( 
.A(n_3504),
.B(n_384),
.Y(n_3651)
);

O2A1O1Ixp33_ASAP7_75t_L g3652 ( 
.A1(n_3406),
.A2(n_386),
.B(n_387),
.C(n_385),
.Y(n_3652)
);

AND2x6_ASAP7_75t_L g3653 ( 
.A(n_3486),
.B(n_10),
.Y(n_3653)
);

BUFx6f_ASAP7_75t_L g3654 ( 
.A(n_3461),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_R g3655 ( 
.A(n_3433),
.B(n_385),
.Y(n_3655)
);

AOI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_3359),
.A2(n_389),
.B(n_388),
.Y(n_3656)
);

OAI22x1_ASAP7_75t_L g3657 ( 
.A1(n_3480),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_3657)
);

BUFx3_ASAP7_75t_L g3658 ( 
.A(n_3547),
.Y(n_3658)
);

OAI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3440),
.A2(n_390),
.B1(n_391),
.B2(n_389),
.Y(n_3659)
);

NOR2xp33_ASAP7_75t_R g3660 ( 
.A(n_3530),
.B(n_390),
.Y(n_3660)
);

AOI21x1_ASAP7_75t_L g3661 ( 
.A1(n_3411),
.A2(n_393),
.B(n_391),
.Y(n_3661)
);

O2A1O1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3391),
.A2(n_394),
.B(n_395),
.C(n_393),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3450),
.Y(n_3663)
);

A2O1A1Ixp33_ASAP7_75t_SL g3664 ( 
.A1(n_3481),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_3664)
);

AOI22xp33_ASAP7_75t_L g3665 ( 
.A1(n_3363),
.A2(n_3511),
.B1(n_3515),
.B2(n_3487),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3455),
.Y(n_3666)
);

NAND3xp33_ASAP7_75t_SL g3667 ( 
.A(n_3370),
.B(n_14),
.C(n_15),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3396),
.B(n_15),
.Y(n_3668)
);

INVx1_ASAP7_75t_SL g3669 ( 
.A(n_3524),
.Y(n_3669)
);

O2A1O1Ixp33_ASAP7_75t_L g3670 ( 
.A1(n_3488),
.A2(n_397),
.B(n_398),
.C(n_396),
.Y(n_3670)
);

AOI221xp5_ASAP7_75t_L g3671 ( 
.A1(n_3422),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.C(n_20),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3446),
.A2(n_400),
.B(n_399),
.Y(n_3672)
);

A2O1A1Ixp33_ASAP7_75t_L g3673 ( 
.A1(n_3375),
.A2(n_20),
.B(n_17),
.C(n_19),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3402),
.B(n_17),
.Y(n_3674)
);

BUFx6f_ASAP7_75t_L g3675 ( 
.A(n_3501),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3403),
.B(n_3407),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3409),
.B(n_19),
.Y(n_3677)
);

BUFx6f_ASAP7_75t_L g3678 ( 
.A(n_3489),
.Y(n_3678)
);

AND2x6_ASAP7_75t_L g3679 ( 
.A(n_3500),
.B(n_20),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3506),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3460),
.A2(n_401),
.B(n_400),
.Y(n_3681)
);

A2O1A1Ixp33_ASAP7_75t_L g3682 ( 
.A1(n_3453),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3682)
);

AOI22xp33_ASAP7_75t_L g3683 ( 
.A1(n_3531),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3470),
.Y(n_3684)
);

INVx3_ASAP7_75t_L g3685 ( 
.A(n_3479),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3413),
.B(n_22),
.Y(n_3686)
);

A2O1A1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3482),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_3687)
);

AOI21x1_ASAP7_75t_L g3688 ( 
.A1(n_3532),
.A2(n_403),
.B(n_402),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3467),
.Y(n_3689)
);

BUFx3_ASAP7_75t_L g3690 ( 
.A(n_3437),
.Y(n_3690)
);

BUFx6f_ASAP7_75t_L g3691 ( 
.A(n_3517),
.Y(n_3691)
);

AO32x1_ASAP7_75t_L g3692 ( 
.A1(n_3338),
.A2(n_27),
.A3(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_3692)
);

AOI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_3536),
.A2(n_405),
.B(n_404),
.Y(n_3693)
);

NOR3xp33_ASAP7_75t_SL g3694 ( 
.A(n_3533),
.B(n_27),
.C(n_28),
.Y(n_3694)
);

NOR3xp33_ASAP7_75t_SL g3695 ( 
.A(n_3542),
.B(n_29),
.C(n_30),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3350),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3521),
.B(n_404),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3421),
.B(n_405),
.Y(n_3698)
);

O2A1O1Ixp5_ASAP7_75t_L g3699 ( 
.A1(n_3492),
.A2(n_407),
.B(n_408),
.C(n_406),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_3508),
.B(n_3400),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3394),
.B(n_29),
.Y(n_3701)
);

BUFx12f_ASAP7_75t_L g3702 ( 
.A(n_3392),
.Y(n_3702)
);

INVx1_ASAP7_75t_SL g3703 ( 
.A(n_3459),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_SL g3704 ( 
.A(n_3438),
.B(n_407),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3498),
.Y(n_3705)
);

AOI22xp5_ASAP7_75t_L g3706 ( 
.A1(n_3377),
.A2(n_410),
.B1(n_411),
.B2(n_409),
.Y(n_3706)
);

A2O1A1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_3485),
.A2(n_3365),
.B(n_3367),
.C(n_3362),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_SL g3708 ( 
.A(n_3477),
.B(n_411),
.Y(n_3708)
);

NOR2xp33_ASAP7_75t_R g3709 ( 
.A(n_3529),
.B(n_412),
.Y(n_3709)
);

NAND3xp33_ASAP7_75t_SL g3710 ( 
.A(n_3484),
.B(n_30),
.C(n_31),
.Y(n_3710)
);

INVx3_ASAP7_75t_L g3711 ( 
.A(n_3483),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3373),
.B(n_31),
.Y(n_3712)
);

O2A1O1Ixp33_ASAP7_75t_SL g3713 ( 
.A1(n_3540),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3390),
.B(n_413),
.Y(n_3714)
);

NOR2xp33_ASAP7_75t_L g3715 ( 
.A(n_3490),
.B(n_414),
.Y(n_3715)
);

A2O1A1Ixp33_ASAP7_75t_L g3716 ( 
.A1(n_3380),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_3716)
);

OAI21xp33_ASAP7_75t_L g3717 ( 
.A1(n_3430),
.A2(n_32),
.B(n_33),
.Y(n_3717)
);

O2A1O1Ixp33_ASAP7_75t_L g3718 ( 
.A1(n_3518),
.A2(n_418),
.B(n_419),
.C(n_417),
.Y(n_3718)
);

NOR2xp67_ASAP7_75t_L g3719 ( 
.A(n_3525),
.B(n_3526),
.Y(n_3719)
);

A2O1A1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_3499),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_3720)
);

INVx4_ASAP7_75t_L g3721 ( 
.A(n_3452),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3528),
.B(n_424),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3384),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_R g3724 ( 
.A(n_3544),
.B(n_424),
.Y(n_3724)
);

OAI22xp5_ASAP7_75t_L g3725 ( 
.A1(n_3505),
.A2(n_426),
.B1(n_427),
.B2(n_425),
.Y(n_3725)
);

AOI21x1_ASAP7_75t_L g3726 ( 
.A1(n_3415),
.A2(n_429),
.B(n_428),
.Y(n_3726)
);

AOI21xp5_ASAP7_75t_L g3727 ( 
.A1(n_3448),
.A2(n_431),
.B(n_430),
.Y(n_3727)
);

INVx5_ASAP7_75t_L g3728 ( 
.A(n_3457),
.Y(n_3728)
);

OAI22x1_ASAP7_75t_L g3729 ( 
.A1(n_3472),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_3729)
);

OAI22xp5_ASAP7_75t_L g3730 ( 
.A1(n_3510),
.A2(n_434),
.B1(n_435),
.B2(n_433),
.Y(n_3730)
);

A2O1A1Ixp33_ASAP7_75t_L g3731 ( 
.A1(n_3410),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3512),
.A2(n_436),
.B1(n_437),
.B2(n_434),
.Y(n_3732)
);

BUFx6f_ASAP7_75t_L g3733 ( 
.A(n_3476),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3478),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3513),
.B(n_437),
.Y(n_3735)
);

INVx2_ASAP7_75t_SL g3736 ( 
.A(n_3509),
.Y(n_3736)
);

AOI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_3497),
.A2(n_439),
.B(n_438),
.Y(n_3737)
);

A2O1A1Ixp33_ASAP7_75t_L g3738 ( 
.A1(n_3439),
.A2(n_41),
.B(n_38),
.C(n_40),
.Y(n_3738)
);

NOR2xp33_ASAP7_75t_L g3739 ( 
.A(n_3346),
.B(n_438),
.Y(n_3739)
);

BUFx6f_ASAP7_75t_L g3740 ( 
.A(n_3339),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3354),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3368),
.B(n_40),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3354),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3354),
.Y(n_3744)
);

AOI22xp33_ASAP7_75t_L g3745 ( 
.A1(n_3439),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3354),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3354),
.Y(n_3747)
);

AOI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_3435),
.A2(n_442),
.B1(n_444),
.B2(n_441),
.Y(n_3748)
);

NOR2xp33_ASAP7_75t_L g3749 ( 
.A(n_3346),
.B(n_441),
.Y(n_3749)
);

NAND2x1p5_ASAP7_75t_L g3750 ( 
.A(n_3348),
.B(n_445),
.Y(n_3750)
);

AOI21xp5_ASAP7_75t_L g3751 ( 
.A1(n_3386),
.A2(n_446),
.B(n_445),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3354),
.Y(n_3752)
);

O2A1O1Ixp33_ASAP7_75t_L g3753 ( 
.A1(n_3346),
.A2(n_447),
.B(n_448),
.C(n_446),
.Y(n_3753)
);

OR2x6_ASAP7_75t_L g3754 ( 
.A(n_3353),
.B(n_447),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3354),
.Y(n_3755)
);

NOR2xp33_ASAP7_75t_L g3756 ( 
.A(n_3346),
.B(n_449),
.Y(n_3756)
);

O2A1O1Ixp33_ASAP7_75t_L g3757 ( 
.A1(n_3346),
.A2(n_452),
.B(n_453),
.C(n_451),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3354),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3744),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3746),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3755),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3569),
.B(n_452),
.Y(n_3762)
);

O2A1O1Ixp5_ASAP7_75t_L g3763 ( 
.A1(n_3599),
.A2(n_3739),
.B(n_3756),
.C(n_3749),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3758),
.Y(n_3764)
);

OAI21xp5_ASAP7_75t_SL g3765 ( 
.A1(n_3562),
.A2(n_44),
.B(n_45),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3676),
.B(n_46),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_SL g3767 ( 
.A(n_3551),
.B(n_454),
.Y(n_3767)
);

NAND3xp33_ASAP7_75t_SL g3768 ( 
.A(n_3655),
.B(n_46),
.C(n_47),
.Y(n_3768)
);

INVx4_ASAP7_75t_L g3769 ( 
.A(n_3586),
.Y(n_3769)
);

INVxp67_ASAP7_75t_L g3770 ( 
.A(n_3571),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3556),
.A2(n_456),
.B(n_455),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3649),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3594),
.A2(n_456),
.B(n_455),
.Y(n_3773)
);

NAND3x1_ASAP7_75t_L g3774 ( 
.A(n_3617),
.B(n_46),
.C(n_47),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3589),
.A2(n_458),
.B(n_457),
.Y(n_3775)
);

AOI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3550),
.A2(n_459),
.B(n_458),
.Y(n_3776)
);

OAI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_3561),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3584),
.A2(n_460),
.B(n_459),
.Y(n_3778)
);

INVx4_ASAP7_75t_L g3779 ( 
.A(n_3586),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3558),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3689),
.B(n_48),
.Y(n_3781)
);

NOR2xp67_ASAP7_75t_L g3782 ( 
.A(n_3592),
.B(n_49),
.Y(n_3782)
);

OAI21x1_ASAP7_75t_L g3783 ( 
.A1(n_3696),
.A2(n_50),
.B(n_51),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3742),
.B(n_50),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3703),
.B(n_461),
.Y(n_3785)
);

OAI21x1_ASAP7_75t_L g3786 ( 
.A1(n_3564),
.A2(n_52),
.B(n_53),
.Y(n_3786)
);

A2O1A1Ixp33_ASAP7_75t_L g3787 ( 
.A1(n_3576),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_L g3788 ( 
.A1(n_3707),
.A2(n_463),
.B(n_462),
.Y(n_3788)
);

BUFx6f_ASAP7_75t_L g3789 ( 
.A(n_3622),
.Y(n_3789)
);

CKINVDCx5p33_ASAP7_75t_R g3790 ( 
.A(n_3552),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3736),
.A2(n_465),
.B(n_464),
.Y(n_3791)
);

AO21x1_ASAP7_75t_L g3792 ( 
.A1(n_3670),
.A2(n_466),
.B(n_465),
.Y(n_3792)
);

CKINVDCx11_ASAP7_75t_R g3793 ( 
.A(n_3557),
.Y(n_3793)
);

AND3x4_ASAP7_75t_L g3794 ( 
.A(n_3565),
.B(n_55),
.C(n_57),
.Y(n_3794)
);

AO31x2_ASAP7_75t_L g3795 ( 
.A1(n_3705),
.A2(n_58),
.A3(n_55),
.B(n_57),
.Y(n_3795)
);

OAI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_3595),
.A2(n_59),
.B(n_60),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3554),
.B(n_60),
.Y(n_3797)
);

AOI221xp5_ASAP7_75t_L g3798 ( 
.A1(n_3698),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.C(n_65),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3669),
.B(n_63),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3574),
.Y(n_3800)
);

INVxp67_ASAP7_75t_SL g3801 ( 
.A(n_3563),
.Y(n_3801)
);

OAI21x1_ASAP7_75t_L g3802 ( 
.A1(n_3560),
.A2(n_64),
.B(n_65),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3642),
.B(n_64),
.Y(n_3803)
);

CKINVDCx20_ASAP7_75t_R g3804 ( 
.A(n_3632),
.Y(n_3804)
);

AO31x2_ASAP7_75t_L g3805 ( 
.A1(n_3721),
.A2(n_67),
.A3(n_65),
.B(n_66),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3723),
.B(n_66),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3688),
.A2(n_67),
.B(n_68),
.Y(n_3807)
);

INVxp67_ASAP7_75t_L g3808 ( 
.A(n_3580),
.Y(n_3808)
);

OAI21x1_ASAP7_75t_L g3809 ( 
.A1(n_3568),
.A2(n_67),
.B(n_68),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3549),
.B(n_68),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3609),
.B(n_69),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3575),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3741),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3572),
.B(n_3697),
.Y(n_3814)
);

OAI21x1_ASAP7_75t_L g3815 ( 
.A1(n_3661),
.A2(n_69),
.B(n_70),
.Y(n_3815)
);

O2A1O1Ixp5_ASAP7_75t_SL g3816 ( 
.A1(n_3711),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3598),
.B(n_71),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3668),
.B(n_71),
.Y(n_3818)
);

AOI22xp5_ASAP7_75t_L g3819 ( 
.A1(n_3621),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_3819)
);

AO32x2_ASAP7_75t_L g3820 ( 
.A1(n_3611),
.A2(n_74),
.A3(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3743),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3674),
.B(n_75),
.Y(n_3822)
);

OAI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3578),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3677),
.B(n_76),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3686),
.B(n_77),
.Y(n_3825)
);

BUFx2_ASAP7_75t_L g3826 ( 
.A(n_3603),
.Y(n_3826)
);

AO31x2_ASAP7_75t_L g3827 ( 
.A1(n_3673),
.A2(n_81),
.A3(n_79),
.B(n_80),
.Y(n_3827)
);

AND2x4_ASAP7_75t_L g3828 ( 
.A(n_3559),
.B(n_470),
.Y(n_3828)
);

OAI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3577),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_3829)
);

AO21x1_ASAP7_75t_L g3830 ( 
.A1(n_3643),
.A2(n_473),
.B(n_471),
.Y(n_3830)
);

AO31x2_ASAP7_75t_L g3831 ( 
.A1(n_3729),
.A2(n_84),
.A3(n_82),
.B(n_83),
.Y(n_3831)
);

BUFx2_ASAP7_75t_L g3832 ( 
.A(n_3604),
.Y(n_3832)
);

OA21x2_ASAP7_75t_L g3833 ( 
.A1(n_3751),
.A2(n_82),
.B(n_84),
.Y(n_3833)
);

AO21x2_ASAP7_75t_L g3834 ( 
.A1(n_3719),
.A2(n_86),
.B(n_87),
.Y(n_3834)
);

O2A1O1Ixp5_ASAP7_75t_L g3835 ( 
.A1(n_3708),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_3835)
);

AOI22xp33_ASAP7_75t_L g3836 ( 
.A1(n_3667),
.A2(n_89),
.B1(n_86),
.B2(n_87),
.Y(n_3836)
);

AOI21x1_ASAP7_75t_L g3837 ( 
.A1(n_3573),
.A2(n_89),
.B(n_90),
.Y(n_3837)
);

OAI21x1_ASAP7_75t_L g3838 ( 
.A1(n_3726),
.A2(n_89),
.B(n_90),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3690),
.B(n_475),
.Y(n_3839)
);

OAI21x1_ASAP7_75t_L g3840 ( 
.A1(n_3734),
.A2(n_90),
.B(n_91),
.Y(n_3840)
);

AO31x2_ASAP7_75t_L g3841 ( 
.A1(n_3682),
.A2(n_93),
.A3(n_91),
.B(n_92),
.Y(n_3841)
);

NAND3x1_ASAP7_75t_L g3842 ( 
.A(n_3748),
.B(n_91),
.C(n_92),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3665),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3747),
.Y(n_3844)
);

AO21x2_ASAP7_75t_L g3845 ( 
.A1(n_3722),
.A2(n_95),
.B(n_96),
.Y(n_3845)
);

AOI21xp5_ASAP7_75t_L g3846 ( 
.A1(n_3566),
.A2(n_3582),
.B(n_3733),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3752),
.Y(n_3847)
);

OAI22xp5_ASAP7_75t_L g3848 ( 
.A1(n_3570),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_3848)
);

INVx1_ASAP7_75t_SL g3849 ( 
.A(n_3555),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3694),
.B(n_95),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3733),
.A2(n_478),
.B(n_477),
.Y(n_3851)
);

AOI21x1_ASAP7_75t_L g3852 ( 
.A1(n_3700),
.A2(n_98),
.B(n_99),
.Y(n_3852)
);

A2O1A1Ixp33_ASAP7_75t_L g3853 ( 
.A1(n_3715),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_3853)
);

OAI22x1_ASAP7_75t_L g3854 ( 
.A1(n_3615),
.A2(n_103),
.B1(n_100),
.B2(n_101),
.Y(n_3854)
);

AO32x2_ASAP7_75t_L g3855 ( 
.A1(n_3618),
.A2(n_104),
.A3(n_100),
.B1(n_103),
.B2(n_105),
.Y(n_3855)
);

OR2x2_ASAP7_75t_L g3856 ( 
.A(n_3620),
.B(n_477),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3638),
.A2(n_480),
.B(n_479),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3745),
.B(n_103),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3680),
.Y(n_3859)
);

AOI21xp5_ASAP7_75t_SL g3860 ( 
.A1(n_3738),
.A2(n_481),
.B(n_480),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3585),
.Y(n_3861)
);

OAI22x1_ASAP7_75t_L g3862 ( 
.A1(n_3706),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_3862)
);

OAI21x1_ASAP7_75t_L g3863 ( 
.A1(n_3737),
.A2(n_105),
.B(n_107),
.Y(n_3863)
);

INVx5_ASAP7_75t_L g3864 ( 
.A(n_3548),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3610),
.B(n_108),
.Y(n_3865)
);

AO31x2_ASAP7_75t_L g3866 ( 
.A1(n_3687),
.A2(n_110),
.A3(n_108),
.B(n_109),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3631),
.B(n_108),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3728),
.A2(n_482),
.B(n_481),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3637),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3645),
.B(n_110),
.Y(n_3870)
);

NOR2xp33_ASAP7_75t_L g3871 ( 
.A(n_3567),
.B(n_3626),
.Y(n_3871)
);

OAI21x1_ASAP7_75t_L g3872 ( 
.A1(n_3693),
.A2(n_111),
.B(n_112),
.Y(n_3872)
);

OAI21x1_ASAP7_75t_SL g3873 ( 
.A1(n_3718),
.A2(n_111),
.B(n_112),
.Y(n_3873)
);

NOR4xp25_ASAP7_75t_L g3874 ( 
.A(n_3753),
.B(n_113),
.C(n_111),
.D(n_112),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3728),
.A2(n_484),
.B(n_483),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3633),
.B(n_484),
.Y(n_3876)
);

OAI22xp5_ASAP7_75t_L g3877 ( 
.A1(n_3608),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_3877)
);

AO21x2_ASAP7_75t_L g3878 ( 
.A1(n_3664),
.A2(n_113),
.B(n_114),
.Y(n_3878)
);

BUFx3_ASAP7_75t_L g3879 ( 
.A(n_3614),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3640),
.Y(n_3880)
);

AO31x2_ASAP7_75t_L g3881 ( 
.A1(n_3720),
.A2(n_116),
.A3(n_114),
.B(n_115),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3684),
.Y(n_3882)
);

OAI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3695),
.A2(n_3650),
.B1(n_3658),
.B2(n_3675),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3663),
.Y(n_3884)
);

INVx4_ASAP7_75t_L g3885 ( 
.A(n_3591),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3666),
.Y(n_3886)
);

AO31x2_ASAP7_75t_L g3887 ( 
.A1(n_3731),
.A2(n_119),
.A3(n_117),
.B(n_118),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3701),
.Y(n_3888)
);

CKINVDCx5p33_ASAP7_75t_R g3889 ( 
.A(n_3636),
.Y(n_3889)
);

AO31x2_ASAP7_75t_L g3890 ( 
.A1(n_3730),
.A2(n_120),
.A3(n_118),
.B(n_119),
.Y(n_3890)
);

AOI21x1_ASAP7_75t_L g3891 ( 
.A1(n_3600),
.A2(n_119),
.B(n_120),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3612),
.Y(n_3892)
);

OAI22xp5_ASAP7_75t_L g3893 ( 
.A1(n_3675),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3691),
.A2(n_486),
.B(n_485),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3691),
.A2(n_487),
.B(n_486),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3717),
.B(n_121),
.Y(n_3896)
);

OAI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3641),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_3897)
);

BUFx5_ASAP7_75t_L g3898 ( 
.A(n_3653),
.Y(n_3898)
);

INVxp67_ASAP7_75t_L g3899 ( 
.A(n_3612),
.Y(n_3899)
);

NOR2x1_ASAP7_75t_SL g3900 ( 
.A(n_3628),
.B(n_489),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3714),
.B(n_124),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3593),
.A2(n_491),
.B(n_490),
.Y(n_3902)
);

CKINVDCx5p33_ASAP7_75t_R g3903 ( 
.A(n_3596),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3683),
.B(n_125),
.Y(n_3904)
);

OAI21x1_ASAP7_75t_L g3905 ( 
.A1(n_3699),
.A2(n_3681),
.B(n_3672),
.Y(n_3905)
);

BUFx6f_ASAP7_75t_L g3906 ( 
.A(n_3740),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3597),
.B(n_126),
.Y(n_3907)
);

NOR2x1_ASAP7_75t_SL g3908 ( 
.A(n_3710),
.B(n_492),
.Y(n_3908)
);

CKINVDCx5p33_ASAP7_75t_R g3909 ( 
.A(n_3660),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3712),
.Y(n_3910)
);

NOR4xp25_ASAP7_75t_L g3911 ( 
.A(n_3757),
.B(n_129),
.C(n_127),
.D(n_128),
.Y(n_3911)
);

BUFx2_ASAP7_75t_L g3912 ( 
.A(n_3740),
.Y(n_3912)
);

OAI21x1_ASAP7_75t_SL g3913 ( 
.A1(n_3623),
.A2(n_127),
.B(n_128),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3651),
.Y(n_3914)
);

AOI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_3727),
.A2(n_495),
.B(n_494),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3713),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3735),
.Y(n_3917)
);

OAI22xp5_ASAP7_75t_L g3918 ( 
.A1(n_3601),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3679),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3581),
.B(n_129),
.Y(n_3920)
);

OAI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3685),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3587),
.B(n_131),
.Y(n_3922)
);

OAI22xp5_ASAP7_75t_L g3923 ( 
.A1(n_3646),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3624),
.A2(n_497),
.B(n_496),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3619),
.B(n_3704),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3553),
.B(n_133),
.Y(n_3926)
);

AOI21xp33_ASAP7_75t_L g3927 ( 
.A1(n_3662),
.A2(n_133),
.B(n_134),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_SL g3928 ( 
.A(n_3763),
.B(n_3724),
.Y(n_3928)
);

OAI22xp5_ASAP7_75t_L g3929 ( 
.A1(n_3814),
.A2(n_3702),
.B1(n_3646),
.B2(n_3754),
.Y(n_3929)
);

CKINVDCx20_ASAP7_75t_R g3930 ( 
.A(n_3804),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3761),
.Y(n_3931)
);

AOI22x1_ASAP7_75t_L g3932 ( 
.A1(n_3796),
.A2(n_3854),
.B1(n_3778),
.B2(n_3862),
.Y(n_3932)
);

CKINVDCx11_ASAP7_75t_R g3933 ( 
.A(n_3793),
.Y(n_3933)
);

OR2x2_ASAP7_75t_L g3934 ( 
.A(n_3917),
.B(n_3647),
.Y(n_3934)
);

AOI22x1_ASAP7_75t_L g3935 ( 
.A1(n_3788),
.A2(n_3657),
.B1(n_3629),
.B2(n_3656),
.Y(n_3935)
);

CKINVDCx5p33_ASAP7_75t_R g3936 ( 
.A(n_3790),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3780),
.Y(n_3937)
);

AO31x2_ASAP7_75t_L g3938 ( 
.A1(n_3792),
.A2(n_3732),
.A3(n_3716),
.B(n_3725),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3849),
.B(n_3583),
.Y(n_3939)
);

OAI21x1_ASAP7_75t_L g3940 ( 
.A1(n_3786),
.A2(n_3652),
.B(n_3635),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3812),
.Y(n_3941)
);

NOR2xp33_ASAP7_75t_R g3942 ( 
.A(n_3903),
.B(n_3678),
.Y(n_3942)
);

HB1xp67_ASAP7_75t_L g3943 ( 
.A(n_3770),
.Y(n_3943)
);

NAND2x1p5_ASAP7_75t_L g3944 ( 
.A(n_3769),
.B(n_3779),
.Y(n_3944)
);

AOI21x1_ASAP7_75t_L g3945 ( 
.A1(n_3846),
.A2(n_3630),
.B(n_3627),
.Y(n_3945)
);

AOI21x1_ASAP7_75t_L g3946 ( 
.A1(n_3891),
.A2(n_3659),
.B(n_3639),
.Y(n_3946)
);

OAI21xp5_ASAP7_75t_L g3947 ( 
.A1(n_3924),
.A2(n_3671),
.B(n_3602),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3888),
.B(n_3644),
.Y(n_3948)
);

OR2x2_ASAP7_75t_L g3949 ( 
.A(n_3910),
.B(n_3625),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3813),
.Y(n_3950)
);

OAI21x1_ASAP7_75t_L g3951 ( 
.A1(n_3905),
.A2(n_3579),
.B(n_3606),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3821),
.Y(n_3952)
);

BUFx3_ASAP7_75t_L g3953 ( 
.A(n_3789),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3844),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3847),
.Y(n_3955)
);

NOR2x1_ASAP7_75t_R g3956 ( 
.A(n_3889),
.B(n_3678),
.Y(n_3956)
);

OAI21x1_ASAP7_75t_L g3957 ( 
.A1(n_3809),
.A2(n_3750),
.B(n_3692),
.Y(n_3957)
);

OAI21x1_ASAP7_75t_L g3958 ( 
.A1(n_3838),
.A2(n_3648),
.B(n_3679),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3797),
.B(n_3709),
.Y(n_3959)
);

INVx6_ASAP7_75t_L g3960 ( 
.A(n_3864),
.Y(n_3960)
);

OAI21x1_ASAP7_75t_L g3961 ( 
.A1(n_3776),
.A2(n_3648),
.B(n_3590),
.Y(n_3961)
);

OAI21x1_ASAP7_75t_L g3962 ( 
.A1(n_3840),
.A2(n_3590),
.B(n_3613),
.Y(n_3962)
);

OAI21x1_ASAP7_75t_L g3963 ( 
.A1(n_3815),
.A2(n_3634),
.B(n_3616),
.Y(n_3963)
);

OAI21x1_ASAP7_75t_L g3964 ( 
.A1(n_3807),
.A2(n_3754),
.B(n_3607),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3859),
.Y(n_3965)
);

OAI21x1_ASAP7_75t_L g3966 ( 
.A1(n_3863),
.A2(n_3654),
.B(n_137),
.Y(n_3966)
);

AOI221xp5_ASAP7_75t_L g3967 ( 
.A1(n_3874),
.A2(n_3605),
.B1(n_3588),
.B2(n_3654),
.C(n_140),
.Y(n_3967)
);

OA21x2_ASAP7_75t_L g3968 ( 
.A1(n_3802),
.A2(n_138),
.B(n_139),
.Y(n_3968)
);

AO21x2_ASAP7_75t_L g3969 ( 
.A1(n_3771),
.A2(n_139),
.B(n_140),
.Y(n_3969)
);

AND2x4_ASAP7_75t_L g3970 ( 
.A(n_3826),
.B(n_498),
.Y(n_3970)
);

OAI22xp5_ASAP7_75t_L g3971 ( 
.A1(n_3762),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_3971)
);

OAI21x1_ASAP7_75t_L g3972 ( 
.A1(n_3872),
.A2(n_141),
.B(n_142),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_3800),
.Y(n_3973)
);

OAI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3787),
.A2(n_141),
.B(n_142),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3772),
.Y(n_3975)
);

OR2x2_ASAP7_75t_L g3976 ( 
.A(n_3901),
.B(n_3759),
.Y(n_3976)
);

BUFx3_ASAP7_75t_L g3977 ( 
.A(n_3789),
.Y(n_3977)
);

BUFx3_ASAP7_75t_L g3978 ( 
.A(n_3912),
.Y(n_3978)
);

AOI221xp5_ASAP7_75t_L g3979 ( 
.A1(n_3911),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.C(n_146),
.Y(n_3979)
);

INVx3_ASAP7_75t_SL g3980 ( 
.A(n_3864),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3882),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3861),
.Y(n_3982)
);

AOI322xp5_ASAP7_75t_L g3983 ( 
.A1(n_3798),
.A2(n_148),
.A3(n_147),
.B1(n_145),
.B2(n_143),
.C1(n_144),
.C2(n_146),
.Y(n_3983)
);

AND2x4_ASAP7_75t_L g3984 ( 
.A(n_3832),
.B(n_3879),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3869),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3760),
.Y(n_3986)
);

OAI222xp33_ASAP7_75t_L g3987 ( 
.A1(n_3819),
.A2(n_147),
.B1(n_149),
.B2(n_145),
.C1(n_146),
.C2(n_148),
.Y(n_3987)
);

OR2x6_ASAP7_75t_L g3988 ( 
.A(n_3860),
.B(n_499),
.Y(n_3988)
);

OAI21x1_ASAP7_75t_L g3989 ( 
.A1(n_3773),
.A2(n_147),
.B(n_148),
.Y(n_3989)
);

OAI21x1_ASAP7_75t_L g3990 ( 
.A1(n_3837),
.A2(n_149),
.B(n_150),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_3892),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3764),
.Y(n_3992)
);

OR2x6_ASAP7_75t_L g3993 ( 
.A(n_3883),
.B(n_500),
.Y(n_3993)
);

OA21x2_ASAP7_75t_L g3994 ( 
.A1(n_3775),
.A2(n_152),
.B(n_153),
.Y(n_3994)
);

HB1xp67_ASAP7_75t_L g3995 ( 
.A(n_3801),
.Y(n_3995)
);

OAI21x1_ASAP7_75t_L g3996 ( 
.A1(n_3783),
.A2(n_153),
.B(n_154),
.Y(n_3996)
);

AOI221xp5_ASAP7_75t_SL g3997 ( 
.A1(n_3853),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.C(n_157),
.Y(n_3997)
);

AOI22xp33_ASAP7_75t_L g3998 ( 
.A1(n_3768),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_3998)
);

OAI22xp5_ASAP7_75t_L g3999 ( 
.A1(n_3871),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3880),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3766),
.B(n_502),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3767),
.B(n_502),
.Y(n_4002)
);

OAI21x1_ASAP7_75t_SL g4003 ( 
.A1(n_3830),
.A2(n_158),
.B(n_159),
.Y(n_4003)
);

AOI221xp5_ASAP7_75t_L g4004 ( 
.A1(n_3803),
.A2(n_3927),
.B1(n_3811),
.B2(n_3765),
.C(n_3823),
.Y(n_4004)
);

OAI22xp5_ASAP7_75t_L g4005 ( 
.A1(n_3774),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3884),
.Y(n_4006)
);

AO21x1_ASAP7_75t_L g4007 ( 
.A1(n_3902),
.A2(n_161),
.B(n_162),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3886),
.Y(n_4008)
);

OA21x2_ASAP7_75t_L g4009 ( 
.A1(n_3916),
.A2(n_162),
.B(n_163),
.Y(n_4009)
);

OAI21x1_ASAP7_75t_L g4010 ( 
.A1(n_3915),
.A2(n_163),
.B(n_164),
.Y(n_4010)
);

HB1xp67_ASAP7_75t_L g4011 ( 
.A(n_3914),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3865),
.B(n_503),
.Y(n_4012)
);

A2O1A1Ixp33_ASAP7_75t_L g4013 ( 
.A1(n_3857),
.A2(n_505),
.B(n_506),
.C(n_504),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3784),
.B(n_504),
.Y(n_4014)
);

AO31x2_ASAP7_75t_L g4015 ( 
.A1(n_3900),
.A2(n_166),
.A3(n_164),
.B(n_165),
.Y(n_4015)
);

NAND2x1p5_ASAP7_75t_L g4016 ( 
.A(n_3885),
.B(n_507),
.Y(n_4016)
);

AND2x4_ASAP7_75t_L g4017 ( 
.A(n_3808),
.B(n_507),
.Y(n_4017)
);

OAI21x1_ASAP7_75t_L g4018 ( 
.A1(n_3791),
.A2(n_165),
.B(n_166),
.Y(n_4018)
);

OAI21x1_ASAP7_75t_L g4019 ( 
.A1(n_3851),
.A2(n_167),
.B(n_168),
.Y(n_4019)
);

CKINVDCx20_ASAP7_75t_R g4020 ( 
.A(n_3909),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3805),
.Y(n_4021)
);

OA21x2_ASAP7_75t_L g4022 ( 
.A1(n_3810),
.A2(n_3875),
.B(n_3868),
.Y(n_4022)
);

AOI21x1_ASAP7_75t_L g4023 ( 
.A1(n_3852),
.A2(n_3843),
.B(n_3806),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_L g4024 ( 
.A1(n_3877),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_4024)
);

INVx3_ASAP7_75t_L g4025 ( 
.A(n_3906),
.Y(n_4025)
);

NOR2xp33_ASAP7_75t_L g4026 ( 
.A(n_3925),
.B(n_508),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3833),
.Y(n_4027)
);

OAI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_3835),
.A2(n_169),
.B(n_170),
.Y(n_4028)
);

AOI22xp33_ASAP7_75t_L g4029 ( 
.A1(n_3836),
.A2(n_173),
.B1(n_170),
.B2(n_172),
.Y(n_4029)
);

OAI21x1_ASAP7_75t_L g4030 ( 
.A1(n_3816),
.A2(n_3895),
.B(n_3894),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3805),
.Y(n_4031)
);

OAI21x1_ASAP7_75t_L g4032 ( 
.A1(n_3873),
.A2(n_173),
.B(n_174),
.Y(n_4032)
);

NAND2x1p5_ASAP7_75t_L g4033 ( 
.A(n_3919),
.B(n_509),
.Y(n_4033)
);

OAI21x1_ASAP7_75t_L g4034 ( 
.A1(n_3913),
.A2(n_175),
.B(n_176),
.Y(n_4034)
);

NOR2x1_ASAP7_75t_SL g4035 ( 
.A(n_3834),
.B(n_509),
.Y(n_4035)
);

AND2x6_ASAP7_75t_L g4036 ( 
.A(n_3907),
.B(n_510),
.Y(n_4036)
);

A2O1A1Ixp33_ASAP7_75t_L g4037 ( 
.A1(n_3920),
.A2(n_512),
.B(n_513),
.C(n_510),
.Y(n_4037)
);

AND2x4_ASAP7_75t_L g4038 ( 
.A(n_3899),
.B(n_512),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3795),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3908),
.B(n_3781),
.Y(n_4040)
);

INVx4_ASAP7_75t_L g4041 ( 
.A(n_3876),
.Y(n_4041)
);

OR2x6_ASAP7_75t_L g4042 ( 
.A(n_4041),
.B(n_3828),
.Y(n_4042)
);

CKINVDCx5p33_ASAP7_75t_R g4043 ( 
.A(n_3933),
.Y(n_4043)
);

AO31x2_ASAP7_75t_L g4044 ( 
.A1(n_4021),
.A2(n_3829),
.A3(n_3777),
.B(n_3848),
.Y(n_4044)
);

OAI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_3928),
.A2(n_3842),
.B(n_3922),
.Y(n_4045)
);

OA21x2_ASAP7_75t_L g4046 ( 
.A1(n_3990),
.A2(n_3839),
.B(n_3822),
.Y(n_4046)
);

A2O1A1Ixp33_ASAP7_75t_L g4047 ( 
.A1(n_3947),
.A2(n_3818),
.B(n_3825),
.C(n_3824),
.Y(n_4047)
);

CKINVDCx5p33_ASAP7_75t_R g4048 ( 
.A(n_3936),
.Y(n_4048)
);

AND2x4_ASAP7_75t_L g4049 ( 
.A(n_3984),
.B(n_3866),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3995),
.B(n_3850),
.Y(n_4050)
);

A2O1A1Ixp33_ASAP7_75t_L g4051 ( 
.A1(n_3974),
.A2(n_3858),
.B(n_3817),
.C(n_3904),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_SL g4052 ( 
.A1(n_3932),
.A2(n_3898),
.B1(n_3878),
.B2(n_3918),
.Y(n_4052)
);

OAI21x1_ASAP7_75t_L g4053 ( 
.A1(n_3951),
.A2(n_3896),
.B(n_3893),
.Y(n_4053)
);

AO31x2_ASAP7_75t_L g4054 ( 
.A1(n_4031),
.A2(n_3897),
.A3(n_3921),
.B(n_3923),
.Y(n_4054)
);

OAI21x1_ASAP7_75t_L g4055 ( 
.A1(n_3940),
.A2(n_3870),
.B(n_3867),
.Y(n_4055)
);

HB1xp67_ASAP7_75t_L g4056 ( 
.A(n_4011),
.Y(n_4056)
);

AOI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3935),
.A2(n_3845),
.B(n_3898),
.Y(n_4057)
);

OA21x2_ASAP7_75t_L g4058 ( 
.A1(n_3957),
.A2(n_3785),
.B(n_3799),
.Y(n_4058)
);

BUFx2_ASAP7_75t_L g4059 ( 
.A(n_3943),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3937),
.Y(n_4060)
);

OAI21x1_ASAP7_75t_L g4061 ( 
.A1(n_4027),
.A2(n_3926),
.B(n_3856),
.Y(n_4061)
);

OAI21x1_ASAP7_75t_L g4062 ( 
.A1(n_3945),
.A2(n_3898),
.B(n_3782),
.Y(n_4062)
);

BUFx6f_ASAP7_75t_L g4063 ( 
.A(n_3953),
.Y(n_4063)
);

AO31x2_ASAP7_75t_L g4064 ( 
.A1(n_4039),
.A2(n_3820),
.A3(n_3855),
.B(n_3827),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3941),
.Y(n_4065)
);

A2O1A1Ixp33_ASAP7_75t_L g4066 ( 
.A1(n_3967),
.A2(n_3794),
.B(n_3898),
.C(n_3881),
.Y(n_4066)
);

BUFx6f_ASAP7_75t_L g4067 ( 
.A(n_3977),
.Y(n_4067)
);

AO31x2_ASAP7_75t_L g4068 ( 
.A1(n_4007),
.A2(n_3841),
.A3(n_3831),
.B(n_3890),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_SL g4069 ( 
.A(n_4040),
.B(n_3831),
.Y(n_4069)
);

BUFx2_ASAP7_75t_L g4070 ( 
.A(n_3978),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3976),
.B(n_3887),
.Y(n_4071)
);

INVx3_ASAP7_75t_L g4072 ( 
.A(n_3960),
.Y(n_4072)
);

OAI21x1_ASAP7_75t_L g4073 ( 
.A1(n_3966),
.A2(n_3841),
.B(n_3887),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3973),
.Y(n_4074)
);

OAI21x1_ASAP7_75t_L g4075 ( 
.A1(n_3972),
.A2(n_3890),
.B(n_177),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3950),
.Y(n_4076)
);

AOI21x1_ASAP7_75t_L g4077 ( 
.A1(n_4023),
.A2(n_177),
.B(n_178),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3952),
.Y(n_4078)
);

A2O1A1Ixp33_ASAP7_75t_L g4079 ( 
.A1(n_4004),
.A2(n_515),
.B(n_516),
.C(n_514),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3986),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3992),
.Y(n_4081)
);

OAI22xp33_ASAP7_75t_L g4082 ( 
.A1(n_3988),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_4000),
.B(n_514),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_4008),
.B(n_515),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3954),
.Y(n_4085)
);

BUFx4f_ASAP7_75t_SL g4086 ( 
.A(n_3930),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3955),
.Y(n_4087)
);

OA21x2_ASAP7_75t_L g4088 ( 
.A1(n_3961),
.A2(n_181),
.B(n_182),
.Y(n_4088)
);

OAI21x1_ASAP7_75t_SL g4089 ( 
.A1(n_4003),
.A2(n_183),
.B(n_184),
.Y(n_4089)
);

AO21x2_ASAP7_75t_L g4090 ( 
.A1(n_4035),
.A2(n_4030),
.B(n_3969),
.Y(n_4090)
);

OA21x2_ASAP7_75t_L g4091 ( 
.A1(n_3958),
.A2(n_183),
.B(n_185),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_3988),
.A2(n_185),
.B(n_186),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3949),
.B(n_517),
.Y(n_4093)
);

AOI21xp5_ASAP7_75t_L g4094 ( 
.A1(n_4028),
.A2(n_185),
.B(n_187),
.Y(n_4094)
);

OA21x2_ASAP7_75t_L g4095 ( 
.A1(n_3996),
.A2(n_187),
.B(n_188),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3931),
.B(n_517),
.Y(n_4096)
);

HB1xp67_ASAP7_75t_L g4097 ( 
.A(n_3982),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3965),
.Y(n_4098)
);

OR2x2_ASAP7_75t_L g4099 ( 
.A(n_3985),
.B(n_518),
.Y(n_4099)
);

AOI22xp33_ASAP7_75t_L g4100 ( 
.A1(n_4036),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_4100)
);

OA21x2_ASAP7_75t_L g4101 ( 
.A1(n_3962),
.A2(n_190),
.B(n_191),
.Y(n_4101)
);

AOI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_4022),
.A2(n_3994),
.B(n_4013),
.Y(n_4102)
);

NAND2x1p5_ASAP7_75t_L g4103 ( 
.A(n_3939),
.B(n_519),
.Y(n_4103)
);

OAI21xp33_ASAP7_75t_L g4104 ( 
.A1(n_3983),
.A2(n_192),
.B(n_193),
.Y(n_4104)
);

NAND3xp33_ASAP7_75t_L g4105 ( 
.A(n_3979),
.B(n_193),
.C(n_194),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_4006),
.B(n_520),
.Y(n_4106)
);

AND2x4_ASAP7_75t_L g4107 ( 
.A(n_3975),
.B(n_521),
.Y(n_4107)
);

OR2x2_ASAP7_75t_L g4108 ( 
.A(n_3948),
.B(n_3934),
.Y(n_4108)
);

HB1xp67_ASAP7_75t_L g4109 ( 
.A(n_3981),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_3989),
.A2(n_195),
.B(n_196),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_4009),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_4015),
.Y(n_4112)
);

BUFx2_ASAP7_75t_L g4113 ( 
.A(n_3942),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4026),
.B(n_4036),
.Y(n_4114)
);

AO21x1_ASAP7_75t_L g4115 ( 
.A1(n_4005),
.A2(n_195),
.B(n_196),
.Y(n_4115)
);

BUFx3_ASAP7_75t_L g4116 ( 
.A(n_4025),
.Y(n_4116)
);

OAI21xp5_ASAP7_75t_L g4117 ( 
.A1(n_4037),
.A2(n_196),
.B(n_197),
.Y(n_4117)
);

AO21x2_ASAP7_75t_L g4118 ( 
.A1(n_3946),
.A2(n_197),
.B(n_198),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4015),
.Y(n_4119)
);

AO31x2_ASAP7_75t_L g4120 ( 
.A1(n_3999),
.A2(n_202),
.A3(n_200),
.B(n_201),
.Y(n_4120)
);

BUFx2_ASAP7_75t_L g4121 ( 
.A(n_3980),
.Y(n_4121)
);

OAI21x1_ASAP7_75t_L g4122 ( 
.A1(n_4010),
.A2(n_4019),
.B(n_4018),
.Y(n_4122)
);

INVx2_ASAP7_75t_L g4123 ( 
.A(n_3968),
.Y(n_4123)
);

CKINVDCx20_ASAP7_75t_R g4124 ( 
.A(n_4020),
.Y(n_4124)
);

OA21x2_ASAP7_75t_L g4125 ( 
.A1(n_4032),
.A2(n_200),
.B(n_201),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4002),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4012),
.Y(n_4127)
);

BUFx4_ASAP7_75t_R g4128 ( 
.A(n_3956),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_4034),
.Y(n_4129)
);

AOI21xp33_ASAP7_75t_SL g4130 ( 
.A1(n_3929),
.A2(n_202),
.B(n_203),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4001),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3959),
.B(n_523),
.Y(n_4132)
);

OAI21x1_ASAP7_75t_SL g4133 ( 
.A1(n_4024),
.A2(n_3971),
.B(n_4014),
.Y(n_4133)
);

OAI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_3963),
.A2(n_204),
.B(n_205),
.Y(n_4134)
);

HB1xp67_ASAP7_75t_L g4135 ( 
.A(n_3964),
.Y(n_4135)
);

OR2x6_ASAP7_75t_L g4136 ( 
.A(n_3993),
.B(n_524),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_3991),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3987),
.A2(n_204),
.B(n_205),
.Y(n_4138)
);

OA21x2_ASAP7_75t_L g4139 ( 
.A1(n_3997),
.A2(n_206),
.B(n_207),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4036),
.Y(n_4140)
);

AO22x1_ASAP7_75t_L g4141 ( 
.A1(n_3970),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_4141)
);

BUFx8_ASAP7_75t_SL g4142 ( 
.A(n_3993),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3938),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4085),
.Y(n_4144)
);

HB1xp67_ASAP7_75t_L g4145 ( 
.A(n_4056),
.Y(n_4145)
);

BUFx3_ASAP7_75t_L g4146 ( 
.A(n_4086),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4060),
.Y(n_4147)
);

INVx3_ASAP7_75t_L g4148 ( 
.A(n_4116),
.Y(n_4148)
);

AO21x1_ASAP7_75t_SL g4149 ( 
.A1(n_4135),
.A2(n_3998),
.B(n_4029),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4070),
.B(n_4108),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_4087),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4050),
.B(n_4140),
.Y(n_4152)
);

INVx4_ASAP7_75t_L g4153 ( 
.A(n_4128),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4109),
.B(n_4017),
.Y(n_4154)
);

AND2x4_ASAP7_75t_L g4155 ( 
.A(n_4049),
.B(n_4038),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_4065),
.Y(n_4156)
);

AO21x2_ASAP7_75t_L g4157 ( 
.A1(n_4119),
.A2(n_3944),
.B(n_4033),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4076),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_4121),
.B(n_4016),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_4078),
.Y(n_4160)
);

INVx2_ASAP7_75t_L g4161 ( 
.A(n_4098),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4080),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4081),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4112),
.Y(n_4164)
);

HB1xp67_ASAP7_75t_L g4165 ( 
.A(n_4071),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_4074),
.Y(n_4166)
);

CKINVDCx11_ASAP7_75t_R g4167 ( 
.A(n_4124),
.Y(n_4167)
);

INVxp67_ASAP7_75t_L g4168 ( 
.A(n_4127),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4111),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4143),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4123),
.Y(n_4171)
);

NOR2xp67_ASAP7_75t_L g4172 ( 
.A(n_4126),
.B(n_208),
.Y(n_4172)
);

OR2x2_ASAP7_75t_L g4173 ( 
.A(n_4069),
.B(n_525),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4129),
.Y(n_4174)
);

BUFx12f_ASAP7_75t_L g4175 ( 
.A(n_4043),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4073),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_4104),
.A2(n_527),
.B1(n_528),
.B2(n_526),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_4061),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4064),
.Y(n_4179)
);

INVxp67_ASAP7_75t_SL g4180 ( 
.A(n_4055),
.Y(n_4180)
);

NOR2xp33_ASAP7_75t_L g4181 ( 
.A(n_4114),
.B(n_526),
.Y(n_4181)
);

INVx3_ASAP7_75t_L g4182 ( 
.A(n_4063),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4106),
.Y(n_4183)
);

INVx3_ASAP7_75t_L g4184 ( 
.A(n_4067),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_4137),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4091),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4088),
.Y(n_4187)
);

HB1xp67_ASAP7_75t_L g4188 ( 
.A(n_4090),
.Y(n_4188)
);

AO21x2_ASAP7_75t_L g4189 ( 
.A1(n_4077),
.A2(n_209),
.B(n_210),
.Y(n_4189)
);

NOR2xp33_ASAP7_75t_L g4190 ( 
.A(n_4142),
.B(n_529),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_4099),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4083),
.Y(n_4192)
);

INVx4_ASAP7_75t_L g4193 ( 
.A(n_4042),
.Y(n_4193)
);

BUFx3_ASAP7_75t_L g4194 ( 
.A(n_4072),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4084),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4068),
.Y(n_4196)
);

OA21x2_ASAP7_75t_L g4197 ( 
.A1(n_4134),
.A2(n_530),
.B(n_529),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4068),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_4122),
.Y(n_4199)
);

AO21x2_ASAP7_75t_L g4200 ( 
.A1(n_4102),
.A2(n_209),
.B(n_210),
.Y(n_4200)
);

HB1xp67_ASAP7_75t_L g4201 ( 
.A(n_4058),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_4131),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4101),
.Y(n_4203)
);

OR2x2_ASAP7_75t_L g4204 ( 
.A(n_4093),
.B(n_530),
.Y(n_4204)
);

HB1xp67_ASAP7_75t_L g4205 ( 
.A(n_4053),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_4096),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_4107),
.Y(n_4207)
);

HB1xp67_ASAP7_75t_L g4208 ( 
.A(n_4046),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4075),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4118),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4095),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4125),
.Y(n_4212)
);

INVx3_ASAP7_75t_SL g4213 ( 
.A(n_4048),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_4062),
.Y(n_4214)
);

INVx2_ASAP7_75t_SL g4215 ( 
.A(n_4132),
.Y(n_4215)
);

INVx3_ASAP7_75t_L g4216 ( 
.A(n_4136),
.Y(n_4216)
);

BUFx5_ASAP7_75t_L g4217 ( 
.A(n_4057),
.Y(n_4217)
);

AO21x2_ASAP7_75t_L g4218 ( 
.A1(n_4130),
.A2(n_211),
.B(n_212),
.Y(n_4218)
);

OR2x2_ASAP7_75t_L g4219 ( 
.A(n_4047),
.B(n_531),
.Y(n_4219)
);

AND2x4_ASAP7_75t_L g4220 ( 
.A(n_4045),
.B(n_532),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4120),
.Y(n_4221)
);

INVx2_ASAP7_75t_L g4222 ( 
.A(n_4089),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4120),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4110),
.Y(n_4224)
);

HB1xp67_ASAP7_75t_L g4225 ( 
.A(n_4139),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4115),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4103),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4044),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4054),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4133),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4052),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_4141),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4066),
.B(n_533),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4094),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4092),
.B(n_4100),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4105),
.Y(n_4236)
);

HB1xp67_ASAP7_75t_L g4237 ( 
.A(n_4117),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_4082),
.Y(n_4238)
);

INVx3_ASAP7_75t_L g4239 ( 
.A(n_4051),
.Y(n_4239)
);

OR2x2_ASAP7_75t_L g4240 ( 
.A(n_4079),
.B(n_4138),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4097),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4097),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4097),
.Y(n_4243)
);

BUFx2_ASAP7_75t_SL g4244 ( 
.A(n_4113),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4097),
.Y(n_4245)
);

HB1xp67_ASAP7_75t_L g4246 ( 
.A(n_4056),
.Y(n_4246)
);

BUFx2_ASAP7_75t_L g4247 ( 
.A(n_4059),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4085),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4097),
.Y(n_4249)
);

NAND3xp33_ASAP7_75t_L g4250 ( 
.A(n_4239),
.B(n_536),
.C(n_534),
.Y(n_4250)
);

AND2x6_ASAP7_75t_L g4251 ( 
.A(n_4230),
.B(n_537),
.Y(n_4251)
);

BUFx6f_ASAP7_75t_L g4252 ( 
.A(n_4175),
.Y(n_4252)
);

AOI22xp5_ASAP7_75t_L g4253 ( 
.A1(n_4231),
.A2(n_539),
.B1(n_540),
.B2(n_538),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4169),
.Y(n_4254)
);

OAI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_4240),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_4255)
);

OAI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_4234),
.A2(n_542),
.B(n_541),
.Y(n_4256)
);

OAI211xp5_ASAP7_75t_L g4257 ( 
.A1(n_4226),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_4257)
);

AOI221xp5_ASAP7_75t_L g4258 ( 
.A1(n_4233),
.A2(n_218),
.B1(n_215),
.B2(n_217),
.C(n_219),
.Y(n_4258)
);

AOI22xp5_ASAP7_75t_L g4259 ( 
.A1(n_4236),
.A2(n_542),
.B1(n_543),
.B2(n_541),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4225),
.A2(n_217),
.B(n_218),
.Y(n_4260)
);

AOI22xp33_ASAP7_75t_L g4261 ( 
.A1(n_4235),
.A2(n_547),
.B1(n_548),
.B2(n_546),
.Y(n_4261)
);

OAI211xp5_ASAP7_75t_L g4262 ( 
.A1(n_4219),
.A2(n_220),
.B(n_218),
.C(n_219),
.Y(n_4262)
);

AOI22xp33_ASAP7_75t_L g4263 ( 
.A1(n_4149),
.A2(n_549),
.B1(n_550),
.B2(n_548),
.Y(n_4263)
);

OAI22xp5_ASAP7_75t_L g4264 ( 
.A1(n_4177),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4150),
.B(n_221),
.Y(n_4265)
);

OAI22xp5_ASAP7_75t_L g4266 ( 
.A1(n_4238),
.A2(n_225),
.B1(n_222),
.B2(n_224),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4171),
.Y(n_4267)
);

INVx4_ASAP7_75t_SL g4268 ( 
.A(n_4213),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_4145),
.B(n_4246),
.Y(n_4269)
);

OAI21x1_ASAP7_75t_L g4270 ( 
.A1(n_4214),
.A2(n_222),
.B(n_224),
.Y(n_4270)
);

NAND2x1_ASAP7_75t_L g4271 ( 
.A(n_4178),
.B(n_224),
.Y(n_4271)
);

OAI22xp5_ASAP7_75t_SL g4272 ( 
.A1(n_4153),
.A2(n_229),
.B1(n_226),
.B2(n_227),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4147),
.Y(n_4273)
);

OR2x6_ASAP7_75t_L g4274 ( 
.A(n_4244),
.B(n_551),
.Y(n_4274)
);

AOI22xp33_ASAP7_75t_SL g4275 ( 
.A1(n_4220),
.A2(n_553),
.B1(n_554),
.B2(n_552),
.Y(n_4275)
);

AOI22xp33_ASAP7_75t_L g4276 ( 
.A1(n_4197),
.A2(n_555),
.B1(n_556),
.B2(n_554),
.Y(n_4276)
);

OAI21x1_ASAP7_75t_L g4277 ( 
.A1(n_4199),
.A2(n_230),
.B(n_231),
.Y(n_4277)
);

OAI22xp5_ASAP7_75t_L g4278 ( 
.A1(n_4232),
.A2(n_4227),
.B1(n_4173),
.B2(n_4222),
.Y(n_4278)
);

OAI21x1_ASAP7_75t_L g4279 ( 
.A1(n_4196),
.A2(n_4198),
.B(n_4176),
.Y(n_4279)
);

AOI22xp33_ASAP7_75t_L g4280 ( 
.A1(n_4224),
.A2(n_557),
.B1(n_559),
.B2(n_555),
.Y(n_4280)
);

OAI211xp5_ASAP7_75t_L g4281 ( 
.A1(n_4221),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4152),
.B(n_232),
.Y(n_4282)
);

AO31x2_ASAP7_75t_L g4283 ( 
.A1(n_4187),
.A2(n_234),
.A3(n_232),
.B(n_233),
.Y(n_4283)
);

OAI22xp5_ASAP7_75t_L g4284 ( 
.A1(n_4168),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_4284)
);

OAI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_4216),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_4285)
);

AOI22xp33_ASAP7_75t_L g4286 ( 
.A1(n_4200),
.A2(n_564),
.B1(n_566),
.B2(n_563),
.Y(n_4286)
);

O2A1O1Ixp33_ASAP7_75t_L g4287 ( 
.A1(n_4223),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_4287)
);

BUFx2_ASAP7_75t_SL g4288 ( 
.A(n_4146),
.Y(n_4288)
);

AND2x2_ASAP7_75t_L g4289 ( 
.A(n_4191),
.B(n_236),
.Y(n_4289)
);

NAND3xp33_ASAP7_75t_L g4290 ( 
.A(n_4205),
.B(n_566),
.C(n_564),
.Y(n_4290)
);

OAI22xp5_ASAP7_75t_L g4291 ( 
.A1(n_4183),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_4291)
);

AO21x2_ASAP7_75t_L g4292 ( 
.A1(n_4188),
.A2(n_238),
.B(n_239),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4158),
.Y(n_4293)
);

AOI221xp5_ASAP7_75t_L g4294 ( 
.A1(n_4181),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.C(n_243),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4241),
.B(n_568),
.Y(n_4295)
);

AND2x4_ASAP7_75t_L g4296 ( 
.A(n_4242),
.B(n_4243),
.Y(n_4296)
);

OAI22xp5_ASAP7_75t_L g4297 ( 
.A1(n_4192),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_4297)
);

AOI221xp5_ASAP7_75t_L g4298 ( 
.A1(n_4195),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.C(n_244),
.Y(n_4298)
);

AND2x4_ASAP7_75t_L g4299 ( 
.A(n_4245),
.B(n_569),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4156),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4160),
.Y(n_4301)
);

INVx4_ASAP7_75t_L g4302 ( 
.A(n_4182),
.Y(n_4302)
);

OAI22xp33_ASAP7_75t_L g4303 ( 
.A1(n_4193),
.A2(n_4172),
.B1(n_4215),
.B2(n_4210),
.Y(n_4303)
);

AOI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_4180),
.A2(n_244),
.B(n_245),
.Y(n_4304)
);

BUFx4f_ASAP7_75t_SL g4305 ( 
.A(n_4194),
.Y(n_4305)
);

NAND3xp33_ASAP7_75t_L g4306 ( 
.A(n_4228),
.B(n_573),
.C(n_572),
.Y(n_4306)
);

AOI21x1_ASAP7_75t_L g4307 ( 
.A1(n_4201),
.A2(n_246),
.B(n_247),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4161),
.Y(n_4308)
);

INVx4_ASAP7_75t_L g4309 ( 
.A(n_4184),
.Y(n_4309)
);

AOI22xp5_ASAP7_75t_L g4310 ( 
.A1(n_4218),
.A2(n_575),
.B1(n_576),
.B2(n_574),
.Y(n_4310)
);

AOI22xp33_ASAP7_75t_L g4311 ( 
.A1(n_4190),
.A2(n_4206),
.B1(n_4159),
.B2(n_4207),
.Y(n_4311)
);

INVx3_ASAP7_75t_L g4312 ( 
.A(n_4148),
.Y(n_4312)
);

AND2x4_ASAP7_75t_L g4313 ( 
.A(n_4249),
.B(n_574),
.Y(n_4313)
);

AOI22xp33_ASAP7_75t_L g4314 ( 
.A1(n_4189),
.A2(n_577),
.B1(n_578),
.B2(n_575),
.Y(n_4314)
);

AND2x4_ASAP7_75t_L g4315 ( 
.A(n_4185),
.B(n_4162),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4170),
.Y(n_4316)
);

AOI22xp33_ASAP7_75t_L g4317 ( 
.A1(n_4209),
.A2(n_582),
.B1(n_584),
.B2(n_580),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4144),
.Y(n_4318)
);

OAI22xp33_ASAP7_75t_L g4319 ( 
.A1(n_4154),
.A2(n_585),
.B1(n_586),
.B2(n_584),
.Y(n_4319)
);

OAI22xp5_ASAP7_75t_L g4320 ( 
.A1(n_4155),
.A2(n_251),
.B1(n_248),
.B2(n_250),
.Y(n_4320)
);

OAI22xp33_ASAP7_75t_L g4321 ( 
.A1(n_4186),
.A2(n_587),
.B1(n_588),
.B2(n_585),
.Y(n_4321)
);

OAI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_4229),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4151),
.B(n_250),
.Y(n_4323)
);

OR2x2_ASAP7_75t_L g4324 ( 
.A(n_4174),
.B(n_252),
.Y(n_4324)
);

AND2x4_ASAP7_75t_L g4325 ( 
.A(n_4163),
.B(n_587),
.Y(n_4325)
);

HB1xp67_ASAP7_75t_L g4326 ( 
.A(n_4208),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_SL g4327 ( 
.A1(n_4157),
.A2(n_590),
.B(n_589),
.Y(n_4327)
);

OAI22xp5_ASAP7_75t_SL g4328 ( 
.A1(n_4204),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_4328)
);

BUFx2_ASAP7_75t_L g4329 ( 
.A(n_4248),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4166),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4212),
.B(n_591),
.Y(n_4331)
);

AO21x2_ASAP7_75t_L g4332 ( 
.A1(n_4203),
.A2(n_4179),
.B(n_4211),
.Y(n_4332)
);

OA21x2_ASAP7_75t_L g4333 ( 
.A1(n_4164),
.A2(n_256),
.B(n_257),
.Y(n_4333)
);

AOI22xp33_ASAP7_75t_L g4334 ( 
.A1(n_4217),
.A2(n_595),
.B1(n_596),
.B2(n_593),
.Y(n_4334)
);

HB1xp67_ASAP7_75t_L g4335 ( 
.A(n_4217),
.Y(n_4335)
);

AOI21xp5_ASAP7_75t_L g4336 ( 
.A1(n_4217),
.A2(n_258),
.B(n_259),
.Y(n_4336)
);

BUFx3_ASAP7_75t_L g4337 ( 
.A(n_4175),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4202),
.Y(n_4338)
);

CKINVDCx5p33_ASAP7_75t_R g4339 ( 
.A(n_4167),
.Y(n_4339)
);

OAI22xp5_ASAP7_75t_L g4340 ( 
.A1(n_4239),
.A2(n_261),
.B1(n_258),
.B2(n_260),
.Y(n_4340)
);

INVxp33_ASAP7_75t_L g4341 ( 
.A(n_4167),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4150),
.B(n_260),
.Y(n_4342)
);

OAI22xp5_ASAP7_75t_SL g4343 ( 
.A1(n_4153),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_4343)
);

OR2x2_ASAP7_75t_L g4344 ( 
.A(n_4165),
.B(n_261),
.Y(n_4344)
);

OAI33xp33_ASAP7_75t_L g4345 ( 
.A1(n_4226),
.A2(n_265),
.A3(n_267),
.B1(n_263),
.B2(n_264),
.B3(n_266),
.Y(n_4345)
);

CKINVDCx20_ASAP7_75t_R g4346 ( 
.A(n_4167),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_4150),
.B(n_264),
.Y(n_4347)
);

AOI22xp33_ASAP7_75t_L g4348 ( 
.A1(n_4239),
.A2(n_598),
.B1(n_599),
.B2(n_597),
.Y(n_4348)
);

AOI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_4239),
.A2(n_598),
.B1(n_600),
.B2(n_597),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4150),
.B(n_265),
.Y(n_4350)
);

HB1xp67_ASAP7_75t_L g4351 ( 
.A(n_4165),
.Y(n_4351)
);

BUFx2_ASAP7_75t_L g4352 ( 
.A(n_4247),
.Y(n_4352)
);

AOI22xp33_ASAP7_75t_SL g4353 ( 
.A1(n_4237),
.A2(n_601),
.B1(n_602),
.B2(n_600),
.Y(n_4353)
);

NAND2x1p5_ASAP7_75t_L g4354 ( 
.A(n_4247),
.B(n_603),
.Y(n_4354)
);

AOI22xp33_ASAP7_75t_L g4355 ( 
.A1(n_4239),
.A2(n_604),
.B1(n_605),
.B2(n_603),
.Y(n_4355)
);

OR2x2_ASAP7_75t_L g4356 ( 
.A(n_4165),
.B(n_266),
.Y(n_4356)
);

OAI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_4239),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4169),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4150),
.B(n_271),
.Y(n_4359)
);

HB1xp67_ASAP7_75t_L g4360 ( 
.A(n_4351),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4312),
.B(n_273),
.Y(n_4361)
);

OR2x2_ASAP7_75t_L g4362 ( 
.A(n_4329),
.B(n_273),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4254),
.Y(n_4363)
);

AND2x4_ASAP7_75t_L g4364 ( 
.A(n_4296),
.B(n_4302),
.Y(n_4364)
);

BUFx2_ASAP7_75t_SL g4365 ( 
.A(n_4346),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4315),
.B(n_606),
.Y(n_4366)
);

HB1xp67_ASAP7_75t_L g4367 ( 
.A(n_4332),
.Y(n_4367)
);

NAND3xp33_ASAP7_75t_L g4368 ( 
.A(n_4336),
.B(n_275),
.C(n_276),
.Y(n_4368)
);

BUFx3_ASAP7_75t_L g4369 ( 
.A(n_4305),
.Y(n_4369)
);

AOI22xp5_ASAP7_75t_L g4370 ( 
.A1(n_4262),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4358),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4316),
.Y(n_4372)
);

AND2x4_ASAP7_75t_L g4373 ( 
.A(n_4309),
.B(n_607),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4278),
.B(n_607),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_4311),
.B(n_278),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4273),
.Y(n_4376)
);

NAND2xp33_ASAP7_75t_L g4377 ( 
.A(n_4339),
.B(n_4252),
.Y(n_4377)
);

HB1xp67_ASAP7_75t_L g4378 ( 
.A(n_4318),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4293),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4300),
.B(n_279),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4267),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4330),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4301),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4338),
.B(n_608),
.Y(n_4384)
);

AND2x2_ASAP7_75t_L g4385 ( 
.A(n_4308),
.B(n_280),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4279),
.Y(n_4386)
);

HB1xp67_ASAP7_75t_L g4387 ( 
.A(n_4324),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4265),
.B(n_281),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4333),
.Y(n_4389)
);

OAI221xp5_ASAP7_75t_SL g4390 ( 
.A1(n_4294),
.A2(n_4258),
.B1(n_4263),
.B2(n_4253),
.C(n_4259),
.Y(n_4390)
);

HB1xp67_ASAP7_75t_L g4391 ( 
.A(n_4344),
.Y(n_4391)
);

HB1xp67_ASAP7_75t_L g4392 ( 
.A(n_4356),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4335),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_4303),
.B(n_4331),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_4342),
.B(n_281),
.Y(n_4395)
);

INVx1_ASAP7_75t_SL g4396 ( 
.A(n_4288),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4323),
.Y(n_4397)
);

OR2x2_ASAP7_75t_L g4398 ( 
.A(n_4295),
.B(n_282),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4347),
.B(n_282),
.Y(n_4399)
);

NOR2x1p5_ASAP7_75t_L g4400 ( 
.A(n_4337),
.B(n_282),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4299),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4350),
.B(n_283),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4292),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4307),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_4313),
.Y(n_4405)
);

INVx2_ASAP7_75t_SL g4406 ( 
.A(n_4268),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4325),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4283),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4359),
.B(n_284),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_4289),
.Y(n_4410)
);

HB1xp67_ASAP7_75t_L g4411 ( 
.A(n_4271),
.Y(n_4411)
);

AND2x2_ASAP7_75t_L g4412 ( 
.A(n_4341),
.B(n_285),
.Y(n_4412)
);

OR2x2_ASAP7_75t_L g4413 ( 
.A(n_4282),
.B(n_285),
.Y(n_4413)
);

BUFx6f_ASAP7_75t_L g4414 ( 
.A(n_4252),
.Y(n_4414)
);

AND2x4_ASAP7_75t_L g4415 ( 
.A(n_4274),
.B(n_611),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4270),
.Y(n_4416)
);

HB1xp67_ASAP7_75t_L g4417 ( 
.A(n_4277),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4251),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4251),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_4354),
.B(n_287),
.Y(n_4420)
);

INVx3_ASAP7_75t_L g4421 ( 
.A(n_4327),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4306),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4290),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4260),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4287),
.Y(n_4425)
);

OR2x2_ASAP7_75t_L g4426 ( 
.A(n_4304),
.B(n_287),
.Y(n_4426)
);

INVxp67_ASAP7_75t_SL g4427 ( 
.A(n_4250),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4276),
.B(n_288),
.Y(n_4428)
);

BUFx6f_ASAP7_75t_L g4429 ( 
.A(n_4272),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_4256),
.B(n_612),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_4310),
.B(n_613),
.Y(n_4431)
);

HB1xp67_ASAP7_75t_L g4432 ( 
.A(n_4284),
.Y(n_4432)
);

AND2x2_ASAP7_75t_L g4433 ( 
.A(n_4275),
.B(n_288),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4328),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4281),
.Y(n_4435)
);

BUFx3_ASAP7_75t_L g4436 ( 
.A(n_4343),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4322),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4319),
.B(n_613),
.Y(n_4438)
);

NAND2x1_ASAP7_75t_L g4439 ( 
.A(n_4286),
.B(n_289),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4255),
.Y(n_4440)
);

INVx2_ASAP7_75t_SL g4441 ( 
.A(n_4320),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_4297),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4291),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4334),
.B(n_615),
.Y(n_4444)
);

OR2x2_ASAP7_75t_L g4445 ( 
.A(n_4266),
.B(n_291),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4257),
.Y(n_4446)
);

OR2x2_ASAP7_75t_L g4447 ( 
.A(n_4285),
.B(n_291),
.Y(n_4447)
);

AOI22xp33_ASAP7_75t_L g4448 ( 
.A1(n_4345),
.A2(n_617),
.B1(n_618),
.B2(n_616),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4261),
.B(n_292),
.Y(n_4449)
);

AND2x2_ASAP7_75t_L g4450 ( 
.A(n_4314),
.B(n_292),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4340),
.Y(n_4451)
);

BUFx2_ASAP7_75t_L g4452 ( 
.A(n_4321),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_4357),
.Y(n_4453)
);

INVxp67_ASAP7_75t_SL g4454 ( 
.A(n_4280),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4264),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4353),
.Y(n_4456)
);

BUFx2_ASAP7_75t_L g4457 ( 
.A(n_4298),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4317),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4348),
.B(n_293),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4349),
.Y(n_4460)
);

NOR2x1p5_ASAP7_75t_L g4461 ( 
.A(n_4355),
.B(n_294),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4269),
.B(n_619),
.Y(n_4462)
);

HB1xp67_ASAP7_75t_L g4463 ( 
.A(n_4326),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4254),
.Y(n_4464)
);

AND2x4_ASAP7_75t_L g4465 ( 
.A(n_4352),
.B(n_620),
.Y(n_4465)
);

AND2x2_ASAP7_75t_L g4466 ( 
.A(n_4352),
.B(n_295),
.Y(n_4466)
);

OR2x2_ASAP7_75t_L g4467 ( 
.A(n_4351),
.B(n_295),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4352),
.B(n_296),
.Y(n_4468)
);

OAI221xp5_ASAP7_75t_SL g4469 ( 
.A1(n_4294),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.C(n_300),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4254),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4254),
.Y(n_4471)
);

BUFx3_ASAP7_75t_L g4472 ( 
.A(n_4369),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4418),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_4419),
.Y(n_4474)
);

AND2x4_ASAP7_75t_SL g4475 ( 
.A(n_4414),
.B(n_298),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4387),
.B(n_300),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4391),
.B(n_300),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4371),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4386),
.Y(n_4479)
);

NAND3xp33_ASAP7_75t_L g4480 ( 
.A(n_4368),
.B(n_301),
.C(n_302),
.Y(n_4480)
);

OR2x2_ASAP7_75t_L g4481 ( 
.A(n_4360),
.B(n_301),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4372),
.Y(n_4482)
);

OR2x2_ASAP7_75t_L g4483 ( 
.A(n_4392),
.B(n_4389),
.Y(n_4483)
);

NAND3xp33_ASAP7_75t_L g4484 ( 
.A(n_4457),
.B(n_4425),
.C(n_4423),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_L g4485 ( 
.A(n_4406),
.B(n_623),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4376),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4393),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_4422),
.B(n_623),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4379),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4464),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4416),
.B(n_624),
.Y(n_4491)
);

OA21x2_ASAP7_75t_L g4492 ( 
.A1(n_4394),
.A2(n_303),
.B(n_304),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4417),
.B(n_626),
.Y(n_4493)
);

AND2x4_ASAP7_75t_L g4494 ( 
.A(n_4407),
.B(n_304),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_4397),
.B(n_4410),
.Y(n_4495)
);

AND2x4_ASAP7_75t_L g4496 ( 
.A(n_4401),
.B(n_4405),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4463),
.B(n_305),
.Y(n_4497)
);

INVx3_ASAP7_75t_L g4498 ( 
.A(n_4465),
.Y(n_4498)
);

OR2x2_ASAP7_75t_L g4499 ( 
.A(n_4408),
.B(n_307),
.Y(n_4499)
);

AND2x2_ASAP7_75t_L g4500 ( 
.A(n_4378),
.B(n_308),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4470),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4424),
.B(n_4403),
.Y(n_4502)
);

AND2x4_ASAP7_75t_L g4503 ( 
.A(n_4361),
.B(n_309),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4471),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4381),
.Y(n_4505)
);

AND2x2_ASAP7_75t_L g4506 ( 
.A(n_4383),
.B(n_309),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4382),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4404),
.B(n_627),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4380),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4385),
.Y(n_4510)
);

OR2x2_ASAP7_75t_L g4511 ( 
.A(n_4462),
.B(n_310),
.Y(n_4511)
);

NAND2x1p5_ASAP7_75t_L g4512 ( 
.A(n_4373),
.B(n_4362),
.Y(n_4512)
);

AND2x4_ASAP7_75t_SL g4513 ( 
.A(n_4415),
.B(n_311),
.Y(n_4513)
);

OAI22xp5_ASAP7_75t_L g4514 ( 
.A1(n_4448),
.A2(n_4390),
.B1(n_4454),
.B2(n_4430),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4384),
.Y(n_4515)
);

INVx3_ASAP7_75t_R g4516 ( 
.A(n_4467),
.Y(n_4516)
);

NOR2xp33_ASAP7_75t_L g4517 ( 
.A(n_4377),
.B(n_627),
.Y(n_4517)
);

INVx1_ASAP7_75t_SL g4518 ( 
.A(n_4365),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4366),
.B(n_628),
.Y(n_4519)
);

OR2x2_ASAP7_75t_L g4520 ( 
.A(n_4440),
.B(n_312),
.Y(n_4520)
);

AND2x2_ASAP7_75t_L g4521 ( 
.A(n_4466),
.B(n_313),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4432),
.B(n_628),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_4374),
.B(n_629),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4367),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4468),
.B(n_313),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_4437),
.B(n_629),
.Y(n_4526)
);

OR2x2_ASAP7_75t_L g4527 ( 
.A(n_4451),
.B(n_314),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4453),
.B(n_315),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4442),
.B(n_315),
.Y(n_4529)
);

OR2x2_ASAP7_75t_L g4530 ( 
.A(n_4443),
.B(n_316),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4398),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4455),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4441),
.B(n_317),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4375),
.B(n_630),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4412),
.B(n_318),
.Y(n_4535)
);

OAI22xp33_ASAP7_75t_L g4536 ( 
.A1(n_4429),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4413),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4420),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4435),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4426),
.Y(n_4540)
);

OR2x6_ASAP7_75t_SL g4541 ( 
.A(n_4456),
.B(n_320),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4460),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4400),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4388),
.B(n_320),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4395),
.B(n_321),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4399),
.B(n_322),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4402),
.B(n_322),
.Y(n_4547)
);

INVx3_ASAP7_75t_L g4548 ( 
.A(n_4429),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4409),
.B(n_323),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4434),
.B(n_323),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4458),
.B(n_4436),
.Y(n_4551)
);

INVxp67_ASAP7_75t_R g4552 ( 
.A(n_4433),
.Y(n_4552)
);

INVxp67_ASAP7_75t_L g4553 ( 
.A(n_4446),
.Y(n_4553)
);

INVx3_ASAP7_75t_L g4554 ( 
.A(n_4431),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4445),
.Y(n_4555)
);

OR2x2_ASAP7_75t_L g4556 ( 
.A(n_4447),
.B(n_324),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4438),
.Y(n_4557)
);

NAND3xp33_ASAP7_75t_L g4558 ( 
.A(n_4469),
.B(n_324),
.C(n_325),
.Y(n_4558)
);

AND2x2_ASAP7_75t_L g4559 ( 
.A(n_4449),
.B(n_325),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4428),
.Y(n_4560)
);

INVx2_ASAP7_75t_L g4561 ( 
.A(n_4439),
.Y(n_4561)
);

OAI21xp5_ASAP7_75t_SL g4562 ( 
.A1(n_4370),
.A2(n_326),
.B(n_327),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4459),
.B(n_327),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4461),
.B(n_329),
.Y(n_4564)
);

OR2x2_ASAP7_75t_L g4565 ( 
.A(n_4444),
.B(n_329),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4450),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4363),
.Y(n_4567)
);

NAND2x1p5_ASAP7_75t_L g4568 ( 
.A(n_4396),
.B(n_330),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4364),
.B(n_330),
.Y(n_4569)
);

OR2x2_ASAP7_75t_L g4570 ( 
.A(n_4360),
.B(n_331),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_4427),
.B(n_631),
.Y(n_4571)
);

OR2x2_ASAP7_75t_L g4572 ( 
.A(n_4360),
.B(n_331),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4427),
.B(n_632),
.Y(n_4573)
);

INVxp67_ASAP7_75t_SL g4574 ( 
.A(n_4411),
.Y(n_4574)
);

INVx2_ASAP7_75t_SL g4575 ( 
.A(n_4406),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4418),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4363),
.Y(n_4577)
);

OAI22xp5_ASAP7_75t_L g4578 ( 
.A1(n_4452),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4364),
.B(n_333),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4363),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4363),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4363),
.Y(n_4582)
);

OAI221xp5_ASAP7_75t_L g4583 ( 
.A1(n_4457),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.C(n_337),
.Y(n_4583)
);

HB1xp67_ASAP7_75t_L g4584 ( 
.A(n_4360),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4427),
.B(n_633),
.Y(n_4585)
);

AND2x4_ASAP7_75t_L g4586 ( 
.A(n_4406),
.B(n_336),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4364),
.B(n_337),
.Y(n_4587)
);

OR2x2_ASAP7_75t_L g4588 ( 
.A(n_4360),
.B(n_338),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4427),
.B(n_634),
.Y(n_4589)
);

AND2x4_ASAP7_75t_L g4590 ( 
.A(n_4406),
.B(n_338),
.Y(n_4590)
);

INVxp67_ASAP7_75t_L g4591 ( 
.A(n_4411),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4363),
.Y(n_4592)
);

INVx2_ASAP7_75t_L g4593 ( 
.A(n_4418),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4363),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4427),
.B(n_634),
.Y(n_4595)
);

BUFx2_ASAP7_75t_L g4596 ( 
.A(n_4411),
.Y(n_4596)
);

BUFx2_ASAP7_75t_L g4597 ( 
.A(n_4411),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4427),
.B(n_636),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4427),
.B(n_637),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4364),
.B(n_339),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4363),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4364),
.B(n_637),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4363),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4364),
.B(n_638),
.Y(n_4604)
);

BUFx6f_ASAP7_75t_L g4605 ( 
.A(n_4414),
.Y(n_4605)
);

BUFx2_ASAP7_75t_SL g4606 ( 
.A(n_4406),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4363),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4363),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4363),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4363),
.Y(n_4610)
);

HB1xp67_ASAP7_75t_L g4611 ( 
.A(n_4360),
.Y(n_4611)
);

OAI221xp5_ASAP7_75t_L g4612 ( 
.A1(n_4457),
.A2(n_641),
.B1(n_639),
.B2(n_640),
.C(n_642),
.Y(n_4612)
);

INVx1_ASAP7_75t_SL g4613 ( 
.A(n_4396),
.Y(n_4613)
);

NAND2x1_ASAP7_75t_SL g4614 ( 
.A(n_4421),
.B(n_639),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4364),
.B(n_641),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4363),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4418),
.Y(n_4617)
);

OR2x2_ASAP7_75t_L g4618 ( 
.A(n_4360),
.B(n_642),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4363),
.Y(n_4619)
);

OR2x2_ASAP7_75t_L g4620 ( 
.A(n_4360),
.B(n_643),
.Y(n_4620)
);

INVx3_ASAP7_75t_L g4621 ( 
.A(n_4605),
.Y(n_4621)
);

OAI31xp33_ASAP7_75t_L g4622 ( 
.A1(n_4514),
.A2(n_1583),
.A3(n_1584),
.B(n_1582),
.Y(n_4622)
);

NAND3xp33_ASAP7_75t_L g4623 ( 
.A(n_4484),
.B(n_644),
.C(n_646),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4557),
.B(n_644),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4606),
.B(n_647),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4478),
.Y(n_4626)
);

AND2x2_ASAP7_75t_L g4627 ( 
.A(n_4575),
.B(n_647),
.Y(n_4627)
);

NAND2x1_ASAP7_75t_L g4628 ( 
.A(n_4596),
.B(n_4597),
.Y(n_4628)
);

INVx1_ASAP7_75t_SL g4629 ( 
.A(n_4614),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4482),
.Y(n_4630)
);

OAI33xp33_ASAP7_75t_L g4631 ( 
.A1(n_4578),
.A2(n_651),
.A3(n_653),
.B1(n_649),
.B2(n_650),
.B3(n_652),
.Y(n_4631)
);

OAI221xp5_ASAP7_75t_L g4632 ( 
.A1(n_4562),
.A2(n_653),
.B1(n_650),
.B2(n_651),
.C(n_654),
.Y(n_4632)
);

INVxp67_ASAP7_75t_SL g4633 ( 
.A(n_4548),
.Y(n_4633)
);

NOR3xp33_ASAP7_75t_SL g4634 ( 
.A(n_4558),
.B(n_4583),
.C(n_4536),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4486),
.Y(n_4635)
);

OAI33xp33_ASAP7_75t_L g4636 ( 
.A1(n_4553),
.A2(n_657),
.A3(n_659),
.B1(n_655),
.B2(n_656),
.B3(n_658),
.Y(n_4636)
);

NOR2x1_ASAP7_75t_L g4637 ( 
.A(n_4492),
.B(n_655),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4489),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4490),
.Y(n_4639)
);

OAI21xp5_ASAP7_75t_SL g4640 ( 
.A1(n_4480),
.A2(n_661),
.B(n_660),
.Y(n_4640)
);

INVxp67_ASAP7_75t_L g4641 ( 
.A(n_4541),
.Y(n_4641)
);

NAND3xp33_ASAP7_75t_L g4642 ( 
.A(n_4612),
.B(n_662),
.C(n_663),
.Y(n_4642)
);

BUFx3_ASAP7_75t_L g4643 ( 
.A(n_4472),
.Y(n_4643)
);

BUFx2_ASAP7_75t_L g4644 ( 
.A(n_4574),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4501),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_SL g4646 ( 
.A(n_4613),
.B(n_666),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4504),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4567),
.Y(n_4648)
);

OR2x2_ASAP7_75t_L g4649 ( 
.A(n_4542),
.B(n_667),
.Y(n_4649)
);

OR2x2_ASAP7_75t_L g4650 ( 
.A(n_4483),
.B(n_667),
.Y(n_4650)
);

NAND3xp33_ASAP7_75t_L g4651 ( 
.A(n_4502),
.B(n_668),
.C(n_669),
.Y(n_4651)
);

AOI21x1_ASAP7_75t_L g4652 ( 
.A1(n_4493),
.A2(n_1586),
.B(n_1576),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4577),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4539),
.B(n_4540),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4518),
.Y(n_4655)
);

HB1xp67_ASAP7_75t_L g4656 ( 
.A(n_4516),
.Y(n_4656)
);

NAND3xp33_ASAP7_75t_L g4657 ( 
.A(n_4591),
.B(n_670),
.C(n_672),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4580),
.Y(n_4658)
);

OR2x2_ASAP7_75t_L g4659 ( 
.A(n_4531),
.B(n_674),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4555),
.B(n_675),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4496),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_4473),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4581),
.Y(n_4663)
);

HB1xp67_ASAP7_75t_L g4664 ( 
.A(n_4584),
.Y(n_4664)
);

OAI31xp33_ASAP7_75t_L g4665 ( 
.A1(n_4568),
.A2(n_1569),
.A3(n_1570),
.B(n_1568),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4474),
.Y(n_4666)
);

OAI31xp33_ASAP7_75t_SL g4667 ( 
.A1(n_4561),
.A2(n_678),
.A3(n_679),
.B(n_677),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4582),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4495),
.B(n_676),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4537),
.B(n_681),
.Y(n_4670)
);

AOI22xp5_ASAP7_75t_L g4671 ( 
.A1(n_4532),
.A2(n_4593),
.B1(n_4617),
.B2(n_4576),
.Y(n_4671)
);

INVx4_ASAP7_75t_L g4672 ( 
.A(n_4586),
.Y(n_4672)
);

OAI33xp33_ASAP7_75t_L g4673 ( 
.A1(n_4571),
.A2(n_687),
.A3(n_689),
.B1(n_684),
.B2(n_685),
.B3(n_688),
.Y(n_4673)
);

NAND3xp33_ASAP7_75t_L g4674 ( 
.A(n_4573),
.B(n_684),
.C(n_685),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4592),
.Y(n_4675)
);

INVx2_ASAP7_75t_L g4676 ( 
.A(n_4538),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4594),
.Y(n_4677)
);

AOI221xp5_ASAP7_75t_L g4678 ( 
.A1(n_4585),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.C(n_696),
.Y(n_4678)
);

OAI21xp5_ASAP7_75t_L g4679 ( 
.A1(n_4589),
.A2(n_694),
.B(n_695),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4551),
.B(n_697),
.Y(n_4680)
);

AO21x2_ASAP7_75t_L g4681 ( 
.A1(n_4524),
.A2(n_698),
.B(n_699),
.Y(n_4681)
);

NAND3xp33_ASAP7_75t_L g4682 ( 
.A(n_4595),
.B(n_698),
.C(n_700),
.Y(n_4682)
);

AND2x4_ASAP7_75t_L g4683 ( 
.A(n_4611),
.B(n_1585),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4554),
.B(n_702),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4601),
.Y(n_4685)
);

AOI21xp33_ASAP7_75t_SL g4686 ( 
.A1(n_4543),
.A2(n_1575),
.B(n_1574),
.Y(n_4686)
);

BUFx6f_ASAP7_75t_L g4687 ( 
.A(n_4590),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4603),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4607),
.Y(n_4689)
);

INVx3_ASAP7_75t_L g4690 ( 
.A(n_4498),
.Y(n_4690)
);

NOR3xp33_ASAP7_75t_L g4691 ( 
.A(n_4598),
.B(n_4599),
.C(n_4523),
.Y(n_4691)
);

OAI22xp33_ASAP7_75t_L g4692 ( 
.A1(n_4552),
.A2(n_708),
.B1(n_706),
.B2(n_707),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4608),
.Y(n_4693)
);

OAI211xp5_ASAP7_75t_SL g4694 ( 
.A1(n_4488),
.A2(n_710),
.B(n_708),
.C(n_709),
.Y(n_4694)
);

NOR2xp33_ASAP7_75t_R g4695 ( 
.A(n_4517),
.B(n_709),
.Y(n_4695)
);

AOI221xp5_ASAP7_75t_L g4696 ( 
.A1(n_4508),
.A2(n_714),
.B1(n_711),
.B2(n_713),
.C(n_715),
.Y(n_4696)
);

OAI33xp33_ASAP7_75t_L g4697 ( 
.A1(n_4522),
.A2(n_717),
.A3(n_720),
.B1(n_715),
.B2(n_716),
.B3(n_719),
.Y(n_4697)
);

OAI31xp33_ASAP7_75t_SL g4698 ( 
.A1(n_4564),
.A2(n_720),
.A3(n_721),
.B(n_717),
.Y(n_4698)
);

INVxp67_ASAP7_75t_L g4699 ( 
.A(n_4499),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4515),
.B(n_716),
.Y(n_4700)
);

AOI22xp33_ASAP7_75t_L g4701 ( 
.A1(n_4566),
.A2(n_723),
.B1(n_721),
.B2(n_722),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4609),
.Y(n_4702)
);

HB1xp67_ASAP7_75t_L g4703 ( 
.A(n_4505),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4509),
.B(n_722),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_4479),
.Y(n_4705)
);

OR2x2_ASAP7_75t_L g4706 ( 
.A(n_4487),
.B(n_4510),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4610),
.Y(n_4707)
);

INVx3_ASAP7_75t_L g4708 ( 
.A(n_4512),
.Y(n_4708)
);

AOI221xp5_ASAP7_75t_L g4709 ( 
.A1(n_4491),
.A2(n_726),
.B1(n_723),
.B2(n_725),
.C(n_727),
.Y(n_4709)
);

BUFx2_ASAP7_75t_L g4710 ( 
.A(n_4500),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4616),
.Y(n_4711)
);

AOI322xp5_ASAP7_75t_L g4712 ( 
.A1(n_4550),
.A2(n_733),
.A3(n_732),
.B1(n_730),
.B2(n_728),
.C1(n_729),
.C2(n_731),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4619),
.Y(n_4713)
);

INVx1_ASAP7_75t_SL g4714 ( 
.A(n_4475),
.Y(n_4714)
);

NAND3xp33_ASAP7_75t_L g4715 ( 
.A(n_4565),
.B(n_729),
.C(n_730),
.Y(n_4715)
);

AOI22xp33_ASAP7_75t_L g4716 ( 
.A1(n_4560),
.A2(n_733),
.B1(n_731),
.B2(n_732),
.Y(n_4716)
);

NOR3xp33_ASAP7_75t_SL g4717 ( 
.A(n_4485),
.B(n_734),
.C(n_735),
.Y(n_4717)
);

INVx2_ASAP7_75t_L g4718 ( 
.A(n_4507),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4506),
.B(n_734),
.Y(n_4719)
);

OR2x2_ASAP7_75t_L g4720 ( 
.A(n_4520),
.B(n_735),
.Y(n_4720)
);

INVx1_ASAP7_75t_SL g4721 ( 
.A(n_4513),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_4569),
.Y(n_4722)
);

AND2x2_ASAP7_75t_SL g4723 ( 
.A(n_4477),
.B(n_736),
.Y(n_4723)
);

NAND4xp25_ASAP7_75t_L g4724 ( 
.A(n_4526),
.B(n_739),
.C(n_740),
.D(n_738),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4579),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4481),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4527),
.B(n_737),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4570),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4656),
.B(n_4637),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4664),
.Y(n_4730)
);

NAND3x1_ASAP7_75t_SL g4731 ( 
.A(n_4665),
.B(n_4497),
.C(n_4476),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4633),
.B(n_4533),
.Y(n_4732)
);

AND2x4_ASAP7_75t_SL g4733 ( 
.A(n_4687),
.B(n_4587),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4655),
.B(n_4529),
.Y(n_4734)
);

HB1xp67_ASAP7_75t_SL g4735 ( 
.A(n_4643),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4710),
.B(n_4528),
.Y(n_4736)
);

HB1xp67_ASAP7_75t_L g4737 ( 
.A(n_4644),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4641),
.B(n_4530),
.Y(n_4738)
);

AND2x4_ASAP7_75t_L g4739 ( 
.A(n_4672),
.B(n_4600),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4687),
.Y(n_4740)
);

AND2x2_ASAP7_75t_L g4741 ( 
.A(n_4690),
.B(n_4602),
.Y(n_4741)
);

OR2x2_ASAP7_75t_L g4742 ( 
.A(n_4726),
.B(n_4556),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4708),
.B(n_4604),
.Y(n_4743)
);

AND2x4_ASAP7_75t_L g4744 ( 
.A(n_4621),
.B(n_4615),
.Y(n_4744)
);

BUFx2_ASAP7_75t_L g4745 ( 
.A(n_4628),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4629),
.B(n_4535),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4718),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4722),
.B(n_4559),
.Y(n_4748)
);

NAND4xp25_ASAP7_75t_L g4749 ( 
.A(n_4622),
.B(n_4534),
.C(n_4519),
.D(n_4563),
.Y(n_4749)
);

INVx3_ASAP7_75t_L g4750 ( 
.A(n_4683),
.Y(n_4750)
);

OR2x2_ASAP7_75t_L g4751 ( 
.A(n_4728),
.B(n_4572),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4626),
.Y(n_4752)
);

INVx1_ASAP7_75t_SL g4753 ( 
.A(n_4714),
.Y(n_4753)
);

NAND2x1_ASAP7_75t_L g4754 ( 
.A(n_4683),
.B(n_4588),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4699),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4630),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4725),
.B(n_4494),
.Y(n_4757)
);

OR2x2_ASAP7_75t_L g4758 ( 
.A(n_4706),
.B(n_4618),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4661),
.B(n_4521),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4676),
.B(n_4620),
.Y(n_4760)
);

HB1xp67_ASAP7_75t_L g4761 ( 
.A(n_4650),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4698),
.B(n_4503),
.Y(n_4762)
);

OR2x2_ASAP7_75t_L g4763 ( 
.A(n_4654),
.B(n_4511),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4635),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4638),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4691),
.B(n_4525),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4625),
.Y(n_4767)
);

OAI221xp5_ASAP7_75t_L g4768 ( 
.A1(n_4634),
.A2(n_4546),
.B1(n_4547),
.B2(n_4545),
.C(n_4544),
.Y(n_4768)
);

NOR2x1_ASAP7_75t_L g4769 ( 
.A(n_4681),
.B(n_4549),
.Y(n_4769)
);

INVx2_ASAP7_75t_L g4770 ( 
.A(n_4660),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4680),
.B(n_741),
.Y(n_4771)
);

INVx2_ASAP7_75t_L g4772 ( 
.A(n_4662),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4666),
.Y(n_4773)
);

NOR3xp33_ASAP7_75t_L g4774 ( 
.A(n_4632),
.B(n_742),
.C(n_743),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4639),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4645),
.Y(n_4776)
);

NOR2xp33_ASAP7_75t_L g4777 ( 
.A(n_4721),
.B(n_747),
.Y(n_4777)
);

AND2x4_ASAP7_75t_L g4778 ( 
.A(n_4627),
.B(n_4684),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4647),
.Y(n_4779)
);

INVx2_ASAP7_75t_SL g4780 ( 
.A(n_4723),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4648),
.Y(n_4781)
);

OR2x6_ASAP7_75t_L g4782 ( 
.A(n_4640),
.B(n_749),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4704),
.B(n_4670),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4669),
.B(n_750),
.Y(n_4784)
);

NOR3xp33_ASAP7_75t_L g4785 ( 
.A(n_4642),
.B(n_751),
.C(n_752),
.Y(n_4785)
);

OR2x2_ASAP7_75t_L g4786 ( 
.A(n_4703),
.B(n_1583),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4653),
.Y(n_4787)
);

INVx2_ASAP7_75t_L g4788 ( 
.A(n_4705),
.Y(n_4788)
);

AND2x2_ASAP7_75t_L g4789 ( 
.A(n_4700),
.B(n_755),
.Y(n_4789)
);

NAND3xp33_ASAP7_75t_SL g4790 ( 
.A(n_4678),
.B(n_756),
.C(n_758),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4658),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4671),
.B(n_759),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4663),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4668),
.Y(n_4794)
);

INVx2_ASAP7_75t_L g4795 ( 
.A(n_4659),
.Y(n_4795)
);

BUFx2_ASAP7_75t_L g4796 ( 
.A(n_4695),
.Y(n_4796)
);

INVx2_ASAP7_75t_SL g4797 ( 
.A(n_4720),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4667),
.B(n_761),
.Y(n_4798)
);

OR2x2_ASAP7_75t_L g4799 ( 
.A(n_4649),
.B(n_1570),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_L g4800 ( 
.A(n_4624),
.B(n_761),
.Y(n_4800)
);

AND2x4_ASAP7_75t_L g4801 ( 
.A(n_4715),
.B(n_4623),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_4727),
.B(n_762),
.Y(n_4802)
);

A2O1A1Ixp33_ASAP7_75t_L g4803 ( 
.A1(n_4712),
.A2(n_766),
.B(n_767),
.C(n_764),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4780),
.B(n_4753),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4755),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4746),
.B(n_4675),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4796),
.B(n_4677),
.Y(n_4807)
);

AND2x2_ASAP7_75t_L g4808 ( 
.A(n_4732),
.B(n_4685),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4769),
.B(n_4686),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_L g4810 ( 
.A(n_4736),
.B(n_4692),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4783),
.B(n_4674),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4767),
.B(n_4682),
.Y(n_4812)
);

AND2x2_ASAP7_75t_L g4813 ( 
.A(n_4739),
.B(n_4688),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4743),
.B(n_4689),
.Y(n_4814)
);

INVx2_ASAP7_75t_L g4815 ( 
.A(n_4733),
.Y(n_4815)
);

AND2x2_ASAP7_75t_L g4816 ( 
.A(n_4741),
.B(n_4693),
.Y(n_4816)
);

NAND2xp33_ASAP7_75t_L g4817 ( 
.A(n_4785),
.B(n_4717),
.Y(n_4817)
);

OR2x2_ASAP7_75t_L g4818 ( 
.A(n_4738),
.B(n_4702),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4730),
.Y(n_4819)
);

AND2x2_ASAP7_75t_L g4820 ( 
.A(n_4740),
.B(n_4707),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4742),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4750),
.B(n_4646),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4734),
.B(n_4679),
.Y(n_4823)
);

AND2x4_ASAP7_75t_L g4824 ( 
.A(n_4744),
.B(n_4711),
.Y(n_4824)
);

INVxp67_ASAP7_75t_SL g4825 ( 
.A(n_4735),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4786),
.Y(n_4826)
);

OR2x2_ASAP7_75t_L g4827 ( 
.A(n_4729),
.B(n_4713),
.Y(n_4827)
);

OAI21xp5_ASAP7_75t_L g4828 ( 
.A1(n_4803),
.A2(n_4651),
.B(n_4657),
.Y(n_4828)
);

INVx2_ASAP7_75t_L g4829 ( 
.A(n_4745),
.Y(n_4829)
);

NAND2xp67_ASAP7_75t_L g4830 ( 
.A(n_4770),
.B(n_4719),
.Y(n_4830)
);

OR2x2_ASAP7_75t_L g4831 ( 
.A(n_4766),
.B(n_4724),
.Y(n_4831)
);

AND3x2_ASAP7_75t_L g4832 ( 
.A(n_4774),
.B(n_4696),
.C(n_4709),
.Y(n_4832)
);

HB1xp67_ASAP7_75t_L g4833 ( 
.A(n_4754),
.Y(n_4833)
);

INVxp67_ASAP7_75t_L g4834 ( 
.A(n_4762),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4751),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4759),
.B(n_4652),
.Y(n_4836)
);

HB1xp67_ASAP7_75t_L g4837 ( 
.A(n_4761),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4797),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4748),
.Y(n_4839)
);

INVx2_ASAP7_75t_L g4840 ( 
.A(n_4778),
.Y(n_4840)
);

OR2x2_ASAP7_75t_L g4841 ( 
.A(n_4758),
.B(n_4716),
.Y(n_4841)
);

OR2x2_ASAP7_75t_L g4842 ( 
.A(n_4760),
.B(n_4701),
.Y(n_4842)
);

OR2x2_ASAP7_75t_L g4843 ( 
.A(n_4763),
.B(n_763),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4795),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4801),
.B(n_4673),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4747),
.Y(n_4846)
);

AND2x2_ASAP7_75t_L g4847 ( 
.A(n_4802),
.B(n_4757),
.Y(n_4847)
);

OAI22xp5_ASAP7_75t_L g4848 ( 
.A1(n_4782),
.A2(n_4636),
.B1(n_4697),
.B2(n_4631),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_L g4849 ( 
.A(n_4788),
.B(n_769),
.Y(n_4849)
);

AND2x2_ASAP7_75t_SL g4850 ( 
.A(n_4798),
.B(n_4694),
.Y(n_4850)
);

AND2x2_ASAP7_75t_L g4851 ( 
.A(n_4784),
.B(n_770),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4772),
.B(n_771),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4771),
.B(n_771),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4752),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4756),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4764),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4799),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4773),
.B(n_772),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_L g4859 ( 
.A(n_4792),
.B(n_773),
.Y(n_4859)
);

OR2x2_ASAP7_75t_L g4860 ( 
.A(n_4749),
.B(n_774),
.Y(n_4860)
);

OR2x2_ASAP7_75t_L g4861 ( 
.A(n_4768),
.B(n_775),
.Y(n_4861)
);

AND2x2_ASAP7_75t_L g4862 ( 
.A(n_4789),
.B(n_775),
.Y(n_4862)
);

NAND2x1_ASAP7_75t_L g4863 ( 
.A(n_4765),
.B(n_778),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4775),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4777),
.B(n_780),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4782),
.B(n_781),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4800),
.B(n_782),
.Y(n_4867)
);

NOR2x1_ASAP7_75t_L g4868 ( 
.A(n_4790),
.B(n_783),
.Y(n_4868)
);

OR2x6_ASAP7_75t_L g4869 ( 
.A(n_4776),
.B(n_4779),
.Y(n_4869)
);

AND2x4_ASAP7_75t_L g4870 ( 
.A(n_4781),
.B(n_786),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4787),
.B(n_787),
.Y(n_4871)
);

AND2x2_ASAP7_75t_L g4872 ( 
.A(n_4791),
.B(n_787),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4793),
.B(n_788),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4794),
.B(n_788),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4731),
.Y(n_4875)
);

INVxp67_ASAP7_75t_SL g4876 ( 
.A(n_4735),
.Y(n_4876)
);

HB1xp67_ASAP7_75t_L g4877 ( 
.A(n_4737),
.Y(n_4877)
);

INVx2_ASAP7_75t_SL g4878 ( 
.A(n_4877),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4825),
.B(n_790),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4837),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4876),
.B(n_792),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4834),
.B(n_793),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4805),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4821),
.Y(n_4884)
);

INVxp33_ASAP7_75t_L g4885 ( 
.A(n_4804),
.Y(n_4885)
);

NOR2xp33_ASAP7_75t_SL g4886 ( 
.A(n_4868),
.B(n_1580),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4835),
.Y(n_4887)
);

OAI21xp5_ASAP7_75t_L g4888 ( 
.A1(n_4809),
.A2(n_794),
.B(n_796),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4807),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_L g4890 ( 
.A(n_4829),
.B(n_801),
.Y(n_4890)
);

AOI22xp5_ASAP7_75t_L g4891 ( 
.A1(n_4848),
.A2(n_804),
.B1(n_801),
.B2(n_802),
.Y(n_4891)
);

INVx2_ASAP7_75t_SL g4892 ( 
.A(n_4863),
.Y(n_4892)
);

OAI21xp33_ASAP7_75t_SL g4893 ( 
.A1(n_4875),
.A2(n_4850),
.B(n_4833),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4872),
.Y(n_4894)
);

INVx2_ASAP7_75t_L g4895 ( 
.A(n_4840),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4808),
.Y(n_4896)
);

AO22x1_ASAP7_75t_L g4897 ( 
.A1(n_4828),
.A2(n_807),
.B1(n_805),
.B2(n_806),
.Y(n_4897)
);

OAI33xp33_ASAP7_75t_L g4898 ( 
.A1(n_4845),
.A2(n_809),
.A3(n_811),
.B1(n_806),
.B2(n_808),
.B3(n_810),
.Y(n_4898)
);

AOI21xp33_ASAP7_75t_L g4899 ( 
.A1(n_4831),
.A2(n_809),
.B(n_810),
.Y(n_4899)
);

INVx1_ASAP7_75t_SL g4900 ( 
.A(n_4836),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4838),
.Y(n_4901)
);

NAND3xp33_ASAP7_75t_L g4902 ( 
.A(n_4832),
.B(n_813),
.C(n_814),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4849),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4806),
.B(n_815),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_4847),
.B(n_1563),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4852),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4858),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4857),
.Y(n_4908)
);

INVx1_ASAP7_75t_SL g4909 ( 
.A(n_4822),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4830),
.B(n_817),
.Y(n_4910)
);

AND2x4_ASAP7_75t_SL g4911 ( 
.A(n_4813),
.B(n_818),
.Y(n_4911)
);

AOI221xp5_ASAP7_75t_L g4912 ( 
.A1(n_4817),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.C(n_822),
.Y(n_4912)
);

NAND3xp33_ASAP7_75t_L g4913 ( 
.A(n_4819),
.B(n_820),
.C(n_823),
.Y(n_4913)
);

OR2x2_ASAP7_75t_L g4914 ( 
.A(n_4810),
.B(n_823),
.Y(n_4914)
);

NOR2xp67_ASAP7_75t_L g4915 ( 
.A(n_4826),
.B(n_1561),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4814),
.B(n_4816),
.Y(n_4916)
);

OR2x2_ASAP7_75t_L g4917 ( 
.A(n_4811),
.B(n_827),
.Y(n_4917)
);

OAI32xp33_ASAP7_75t_L g4918 ( 
.A1(n_4861),
.A2(n_4860),
.A3(n_4841),
.B1(n_4842),
.B2(n_4812),
.Y(n_4918)
);

AOI22xp33_ASAP7_75t_L g4919 ( 
.A1(n_4823),
.A2(n_830),
.B1(n_828),
.B2(n_829),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4824),
.B(n_828),
.Y(n_4920)
);

AND2x2_ASAP7_75t_L g4921 ( 
.A(n_4820),
.B(n_1580),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_L g4922 ( 
.A(n_4844),
.B(n_831),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4839),
.B(n_833),
.Y(n_4923)
);

NAND3x2_ASAP7_75t_L g4924 ( 
.A(n_4818),
.B(n_833),
.C(n_836),
.Y(n_4924)
);

INVxp67_ASAP7_75t_L g4925 ( 
.A(n_4866),
.Y(n_4925)
);

INVxp33_ASAP7_75t_L g4926 ( 
.A(n_4865),
.Y(n_4926)
);

INVxp67_ASAP7_75t_L g4927 ( 
.A(n_4869),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4843),
.Y(n_4928)
);

OAI22xp33_ASAP7_75t_SL g4929 ( 
.A1(n_4827),
.A2(n_840),
.B1(n_838),
.B2(n_839),
.Y(n_4929)
);

INVx2_ASAP7_75t_L g4930 ( 
.A(n_4870),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4862),
.Y(n_4931)
);

OAI22xp33_ASAP7_75t_SL g4932 ( 
.A1(n_4846),
.A2(n_844),
.B1(n_841),
.B2(n_843),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4851),
.Y(n_4933)
);

AO22x1_ASAP7_75t_L g4934 ( 
.A1(n_4859),
.A2(n_4855),
.B1(n_4856),
.B2(n_4854),
.Y(n_4934)
);

AOI22xp5_ASAP7_75t_L g4935 ( 
.A1(n_4864),
.A2(n_848),
.B1(n_846),
.B2(n_847),
.Y(n_4935)
);

INVx2_ASAP7_75t_L g4936 ( 
.A(n_4853),
.Y(n_4936)
);

AOI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4871),
.A2(n_853),
.B1(n_850),
.B2(n_852),
.Y(n_4937)
);

AOI22xp5_ASAP7_75t_L g4938 ( 
.A1(n_4873),
.A2(n_856),
.B1(n_854),
.B2(n_855),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4874),
.Y(n_4939)
);

OAI22xp33_ASAP7_75t_L g4940 ( 
.A1(n_4867),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_L g4941 ( 
.A(n_4825),
.B(n_857),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_4815),
.Y(n_4942)
);

A2O1A1Ixp33_ASAP7_75t_L g4943 ( 
.A1(n_4828),
.A2(n_1581),
.B(n_1577),
.C(n_863),
.Y(n_4943)
);

AND2x2_ASAP7_75t_L g4944 ( 
.A(n_4825),
.B(n_1573),
.Y(n_4944)
);

INVx2_ASAP7_75t_SL g4945 ( 
.A(n_4877),
.Y(n_4945)
);

AOI21xp33_ASAP7_75t_L g4946 ( 
.A1(n_4885),
.A2(n_1577),
.B(n_1573),
.Y(n_4946)
);

OAI22xp33_ASAP7_75t_L g4947 ( 
.A1(n_4891),
.A2(n_863),
.B1(n_860),
.B2(n_862),
.Y(n_4947)
);

OAI22xp33_ASAP7_75t_L g4948 ( 
.A1(n_4902),
.A2(n_865),
.B1(n_862),
.B2(n_864),
.Y(n_4948)
);

AOI211x1_ASAP7_75t_L g4949 ( 
.A1(n_4934),
.A2(n_866),
.B(n_864),
.C(n_865),
.Y(n_4949)
);

OA21x2_ASAP7_75t_L g4950 ( 
.A1(n_4910),
.A2(n_868),
.B(n_872),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4878),
.Y(n_4951)
);

AND2x2_ASAP7_75t_L g4952 ( 
.A(n_4916),
.B(n_872),
.Y(n_4952)
);

AOI32xp33_ASAP7_75t_L g4953 ( 
.A1(n_4893),
.A2(n_875),
.A3(n_873),
.B1(n_874),
.B2(n_876),
.Y(n_4953)
);

O2A1O1Ixp33_ASAP7_75t_L g4954 ( 
.A1(n_4943),
.A2(n_880),
.B(n_876),
.C(n_878),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4945),
.Y(n_4955)
);

INVx1_ASAP7_75t_SL g4956 ( 
.A(n_4911),
.Y(n_4956)
);

AOI21xp33_ASAP7_75t_L g4957 ( 
.A1(n_4900),
.A2(n_4926),
.B(n_4927),
.Y(n_4957)
);

NOR3xp33_ASAP7_75t_L g4958 ( 
.A(n_4925),
.B(n_881),
.C(n_882),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4880),
.Y(n_4959)
);

XNOR2x1_ASAP7_75t_L g4960 ( 
.A(n_4924),
.B(n_4897),
.Y(n_4960)
);

OAI221xp5_ASAP7_75t_L g4961 ( 
.A1(n_4888),
.A2(n_885),
.B1(n_883),
.B2(n_884),
.C(n_886),
.Y(n_4961)
);

OAI321xp33_ASAP7_75t_L g4962 ( 
.A1(n_4889),
.A2(n_887),
.A3(n_889),
.B1(n_885),
.B2(n_886),
.C(n_888),
.Y(n_4962)
);

OAI22xp33_ASAP7_75t_L g4963 ( 
.A1(n_4914),
.A2(n_890),
.B1(n_888),
.B2(n_889),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4879),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4881),
.Y(n_4965)
);

NAND2x1_ASAP7_75t_L g4966 ( 
.A(n_4930),
.B(n_1555),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4941),
.Y(n_4967)
);

XOR2x2_ASAP7_75t_L g4968 ( 
.A(n_4912),
.B(n_890),
.Y(n_4968)
);

OAI22xp5_ASAP7_75t_L g4969 ( 
.A1(n_4909),
.A2(n_893),
.B1(n_891),
.B2(n_892),
.Y(n_4969)
);

NAND2xp33_ASAP7_75t_L g4970 ( 
.A(n_4928),
.B(n_894),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_4905),
.B(n_894),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4942),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4921),
.B(n_896),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4896),
.Y(n_4974)
);

OAI21xp33_ASAP7_75t_L g4975 ( 
.A1(n_4895),
.A2(n_897),
.B(n_898),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4931),
.B(n_898),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4933),
.B(n_899),
.Y(n_4977)
);

INVxp67_ASAP7_75t_SL g4978 ( 
.A(n_4932),
.Y(n_4978)
);

OAI221xp5_ASAP7_75t_L g4979 ( 
.A1(n_4919),
.A2(n_904),
.B1(n_901),
.B2(n_902),
.C(n_906),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4899),
.A2(n_901),
.B(n_906),
.Y(n_4980)
);

AOI211xp5_ASAP7_75t_L g4981 ( 
.A1(n_4929),
.A2(n_910),
.B(n_908),
.C(n_909),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4936),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4890),
.Y(n_4983)
);

AOI322xp5_ASAP7_75t_L g4984 ( 
.A1(n_4883),
.A2(n_916),
.A3(n_915),
.B1(n_913),
.B2(n_911),
.C1(n_912),
.C2(n_914),
.Y(n_4984)
);

OAI22xp5_ASAP7_75t_L g4985 ( 
.A1(n_4913),
.A2(n_914),
.B1(n_912),
.B2(n_913),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4894),
.Y(n_4986)
);

NOR2xp33_ASAP7_75t_L g4987 ( 
.A(n_4898),
.B(n_917),
.Y(n_4987)
);

AOI22xp5_ASAP7_75t_L g4988 ( 
.A1(n_4901),
.A2(n_922),
.B1(n_918),
.B2(n_921),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4908),
.B(n_924),
.Y(n_4989)
);

AOI22xp33_ASAP7_75t_L g4990 ( 
.A1(n_4939),
.A2(n_927),
.B1(n_925),
.B2(n_926),
.Y(n_4990)
);

AOI22xp33_ASAP7_75t_L g4991 ( 
.A1(n_4903),
.A2(n_929),
.B1(n_927),
.B2(n_928),
.Y(n_4991)
);

OAI21xp5_ASAP7_75t_SL g4992 ( 
.A1(n_4884),
.A2(n_1572),
.B(n_928),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4887),
.B(n_929),
.Y(n_4993)
);

OR2x2_ASAP7_75t_L g4994 ( 
.A(n_4917),
.B(n_930),
.Y(n_4994)
);

OAI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4882),
.A2(n_931),
.B(n_932),
.Y(n_4995)
);

AOI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4940),
.A2(n_934),
.B(n_935),
.Y(n_4996)
);

OAI211xp5_ASAP7_75t_SL g4997 ( 
.A1(n_4906),
.A2(n_938),
.B(n_936),
.C(n_937),
.Y(n_4997)
);

OAI21xp5_ASAP7_75t_L g4998 ( 
.A1(n_4935),
.A2(n_939),
.B(n_940),
.Y(n_4998)
);

AOI22xp33_ASAP7_75t_L g4999 ( 
.A1(n_4907),
.A2(n_942),
.B1(n_940),
.B2(n_941),
.Y(n_4999)
);

OR2x2_ASAP7_75t_L g5000 ( 
.A(n_4904),
.B(n_943),
.Y(n_5000)
);

AOI22xp5_ASAP7_75t_L g5001 ( 
.A1(n_4922),
.A2(n_946),
.B1(n_944),
.B2(n_945),
.Y(n_5001)
);

OAI32xp33_ASAP7_75t_L g5002 ( 
.A1(n_4923),
.A2(n_947),
.A3(n_949),
.B1(n_946),
.B2(n_948),
.Y(n_5002)
);

AND2x4_ASAP7_75t_L g5003 ( 
.A(n_4920),
.B(n_944),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4937),
.B(n_950),
.Y(n_5004)
);

INVxp67_ASAP7_75t_SL g5005 ( 
.A(n_4938),
.Y(n_5005)
);

NAND2xp33_ASAP7_75t_SL g5006 ( 
.A(n_4892),
.B(n_951),
.Y(n_5006)
);

INVx2_ASAP7_75t_L g5007 ( 
.A(n_4892),
.Y(n_5007)
);

AND2x2_ASAP7_75t_L g5008 ( 
.A(n_4916),
.B(n_954),
.Y(n_5008)
);

AOI221xp5_ASAP7_75t_L g5009 ( 
.A1(n_4918),
.A2(n_969),
.B1(n_975),
.B2(n_962),
.C(n_954),
.Y(n_5009)
);

AOI22xp33_ASAP7_75t_SL g5010 ( 
.A1(n_4886),
.A2(n_958),
.B1(n_956),
.B2(n_957),
.Y(n_5010)
);

A2O1A1Ixp33_ASAP7_75t_L g5011 ( 
.A1(n_4891),
.A2(n_960),
.B(n_958),
.C(n_959),
.Y(n_5011)
);

AND2x2_ASAP7_75t_L g5012 ( 
.A(n_4916),
.B(n_959),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_4944),
.B(n_962),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_L g5014 ( 
.A(n_4944),
.B(n_963),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4892),
.Y(n_5015)
);

BUFx2_ASAP7_75t_L g5016 ( 
.A(n_4892),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4944),
.Y(n_5017)
);

AOI33xp33_ASAP7_75t_L g5018 ( 
.A1(n_4900),
.A2(n_968),
.A3(n_970),
.B1(n_964),
.B2(n_966),
.B3(n_969),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4944),
.Y(n_5019)
);

OAI21xp5_ASAP7_75t_L g5020 ( 
.A1(n_4891),
.A2(n_970),
.B(n_971),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4944),
.B(n_972),
.Y(n_5021)
);

HB1xp67_ASAP7_75t_L g5022 ( 
.A(n_4915),
.Y(n_5022)
);

OA21x2_ASAP7_75t_L g5023 ( 
.A1(n_4891),
.A2(n_973),
.B(n_974),
.Y(n_5023)
);

OAI211xp5_ASAP7_75t_SL g5024 ( 
.A1(n_4891),
.A2(n_979),
.B(n_977),
.C(n_978),
.Y(n_5024)
);

OAI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_4891),
.A2(n_980),
.B(n_981),
.Y(n_5025)
);

AOI211xp5_ASAP7_75t_SL g5026 ( 
.A1(n_4957),
.A2(n_988),
.B(n_991),
.C(n_981),
.Y(n_5026)
);

AND2x4_ASAP7_75t_L g5027 ( 
.A(n_5016),
.B(n_1566),
.Y(n_5027)
);

INVxp67_ASAP7_75t_L g5028 ( 
.A(n_5022),
.Y(n_5028)
);

AOI221xp5_ASAP7_75t_L g5029 ( 
.A1(n_4978),
.A2(n_1571),
.B1(n_985),
.B2(n_982),
.C(n_984),
.Y(n_5029)
);

INVxp67_ASAP7_75t_L g5030 ( 
.A(n_5006),
.Y(n_5030)
);

AOI22xp33_ASAP7_75t_L g5031 ( 
.A1(n_5005),
.A2(n_4960),
.B1(n_4955),
.B2(n_4951),
.Y(n_5031)
);

A2O1A1Ixp33_ASAP7_75t_L g5032 ( 
.A1(n_4953),
.A2(n_987),
.B(n_985),
.C(n_986),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4956),
.B(n_986),
.Y(n_5033)
);

INVx2_ASAP7_75t_L g5034 ( 
.A(n_5007),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_5015),
.Y(n_5035)
);

HB1xp67_ASAP7_75t_L g5036 ( 
.A(n_4966),
.Y(n_5036)
);

OAI32xp33_ASAP7_75t_L g5037 ( 
.A1(n_4987),
.A2(n_1007),
.A3(n_1016),
.B1(n_998),
.B2(n_992),
.Y(n_5037)
);

AND2x2_ASAP7_75t_L g5038 ( 
.A(n_5017),
.B(n_993),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_5019),
.B(n_994),
.Y(n_5039)
);

AOI222xp33_ASAP7_75t_L g5040 ( 
.A1(n_5009),
.A2(n_1002),
.B1(n_1004),
.B2(n_999),
.C1(n_1000),
.C2(n_1003),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4952),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_5008),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_5012),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4994),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_L g5045 ( 
.A(n_4949),
.B(n_1005),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4973),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4981),
.B(n_1009),
.Y(n_5047)
);

OR2x2_ASAP7_75t_L g5048 ( 
.A(n_4972),
.B(n_1012),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4971),
.Y(n_5049)
);

O2A1O1Ixp5_ASAP7_75t_L g5050 ( 
.A1(n_4959),
.A2(n_1015),
.B(n_1013),
.C(n_1014),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_5003),
.B(n_1018),
.Y(n_5051)
);

OAI31xp33_ASAP7_75t_SL g5052 ( 
.A1(n_5024),
.A2(n_4948),
.A3(n_4997),
.B(n_5010),
.Y(n_5052)
);

AND2x2_ASAP7_75t_L g5053 ( 
.A(n_4982),
.B(n_1019),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4989),
.Y(n_5054)
);

AOI21xp33_ASAP7_75t_SL g5055 ( 
.A1(n_5023),
.A2(n_1556),
.B(n_1554),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_5018),
.B(n_1020),
.Y(n_5056)
);

AOI22xp5_ASAP7_75t_L g5057 ( 
.A1(n_4968),
.A2(n_1559),
.B1(n_1560),
.B2(n_1558),
.Y(n_5057)
);

A2O1A1Ixp33_ASAP7_75t_L g5058 ( 
.A1(n_4954),
.A2(n_1027),
.B(n_1024),
.C(n_1025),
.Y(n_5058)
);

AOI22xp5_ASAP7_75t_L g5059 ( 
.A1(n_4970),
.A2(n_1543),
.B1(n_1544),
.B2(n_1542),
.Y(n_5059)
);

AND2x2_ASAP7_75t_L g5060 ( 
.A(n_4964),
.B(n_4965),
.Y(n_5060)
);

AND2x2_ASAP7_75t_L g5061 ( 
.A(n_4967),
.B(n_1030),
.Y(n_5061)
);

A2O1A1Ixp33_ASAP7_75t_L g5062 ( 
.A1(n_4962),
.A2(n_4996),
.B(n_4980),
.C(n_4984),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_5013),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_5014),
.Y(n_5064)
);

OA22x2_ASAP7_75t_L g5065 ( 
.A1(n_4992),
.A2(n_4986),
.B1(n_4974),
.B2(n_5020),
.Y(n_5065)
);

OAI22xp5_ASAP7_75t_L g5066 ( 
.A1(n_5011),
.A2(n_1036),
.B1(n_1034),
.B2(n_1035),
.Y(n_5066)
);

INVx2_ASAP7_75t_L g5067 ( 
.A(n_5000),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_4963),
.B(n_1036),
.Y(n_5068)
);

OAI21xp5_ASAP7_75t_SL g5069 ( 
.A1(n_5025),
.A2(n_1037),
.B(n_1038),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4947),
.B(n_1037),
.Y(n_5070)
);

AOI211xp5_ASAP7_75t_SL g5071 ( 
.A1(n_4983),
.A2(n_1044),
.B(n_1053),
.C(n_1038),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_5021),
.Y(n_5072)
);

NAND3xp33_ASAP7_75t_SL g5073 ( 
.A(n_4958),
.B(n_1039),
.C(n_1040),
.Y(n_5073)
);

INVx1_ASAP7_75t_SL g5074 ( 
.A(n_4950),
.Y(n_5074)
);

AOI21xp33_ASAP7_75t_SL g5075 ( 
.A1(n_4950),
.A2(n_4969),
.B(n_4985),
.Y(n_5075)
);

O2A1O1Ixp33_ASAP7_75t_L g5076 ( 
.A1(n_5002),
.A2(n_1043),
.B(n_1041),
.C(n_1042),
.Y(n_5076)
);

AOI21xp5_ASAP7_75t_L g5077 ( 
.A1(n_5004),
.A2(n_1043),
.B(n_1044),
.Y(n_5077)
);

NOR2xp33_ASAP7_75t_L g5078 ( 
.A(n_4975),
.B(n_1045),
.Y(n_5078)
);

NAND4xp25_ASAP7_75t_L g5079 ( 
.A(n_4998),
.B(n_1049),
.C(n_1046),
.D(n_1047),
.Y(n_5079)
);

INVx2_ASAP7_75t_SL g5080 ( 
.A(n_5027),
.Y(n_5080)
);

OAI211xp5_ASAP7_75t_SL g5081 ( 
.A1(n_5031),
.A2(n_4961),
.B(n_4995),
.C(n_4946),
.Y(n_5081)
);

OAI221xp5_ASAP7_75t_L g5082 ( 
.A1(n_5052),
.A2(n_4979),
.B1(n_4990),
.B2(n_4999),
.C(n_4991),
.Y(n_5082)
);

OAI21xp5_ASAP7_75t_L g5083 ( 
.A1(n_5062),
.A2(n_4977),
.B(n_4976),
.Y(n_5083)
);

NAND2x1p5_ASAP7_75t_L g5084 ( 
.A(n_5027),
.B(n_4988),
.Y(n_5084)
);

O2A1O1Ixp33_ASAP7_75t_L g5085 ( 
.A1(n_5032),
.A2(n_4993),
.B(n_5001),
.C(n_1053),
.Y(n_5085)
);

OAI21xp5_ASAP7_75t_L g5086 ( 
.A1(n_5028),
.A2(n_1051),
.B(n_1054),
.Y(n_5086)
);

AOI221xp5_ASAP7_75t_L g5087 ( 
.A1(n_5037),
.A2(n_1057),
.B1(n_1055),
.B2(n_1056),
.C(n_1058),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_5033),
.Y(n_5088)
);

OAI22xp5_ASAP7_75t_L g5089 ( 
.A1(n_5057),
.A2(n_1063),
.B1(n_1061),
.B2(n_1062),
.Y(n_5089)
);

O2A1O1Ixp33_ASAP7_75t_L g5090 ( 
.A1(n_5058),
.A2(n_1066),
.B(n_1064),
.C(n_1065),
.Y(n_5090)
);

OAI221xp5_ASAP7_75t_L g5091 ( 
.A1(n_5029),
.A2(n_1069),
.B1(n_1067),
.B2(n_1068),
.C(n_1070),
.Y(n_5091)
);

OAI222xp33_ASAP7_75t_L g5092 ( 
.A1(n_5065),
.A2(n_1553),
.B1(n_1551),
.B2(n_1552),
.C1(n_1546),
.C2(n_1074),
.Y(n_5092)
);

AOI22xp5_ASAP7_75t_L g5093 ( 
.A1(n_5034),
.A2(n_1075),
.B1(n_1072),
.B2(n_1073),
.Y(n_5093)
);

AOI221xp5_ASAP7_75t_L g5094 ( 
.A1(n_5076),
.A2(n_1078),
.B1(n_1075),
.B2(n_1077),
.C(n_1079),
.Y(n_5094)
);

AOI22xp5_ASAP7_75t_L g5095 ( 
.A1(n_5035),
.A2(n_1080),
.B1(n_1077),
.B2(n_1079),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_5077),
.A2(n_1080),
.B(n_1081),
.Y(n_5096)
);

AOI21xp5_ASAP7_75t_L g5097 ( 
.A1(n_5045),
.A2(n_1082),
.B(n_1083),
.Y(n_5097)
);

AOI21xp33_ASAP7_75t_L g5098 ( 
.A1(n_5041),
.A2(n_1083),
.B(n_1084),
.Y(n_5098)
);

NOR2xp33_ASAP7_75t_L g5099 ( 
.A(n_5042),
.B(n_5043),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_5071),
.B(n_1088),
.Y(n_5100)
);

NAND3xp33_ASAP7_75t_SL g5101 ( 
.A(n_5026),
.B(n_1091),
.C(n_1090),
.Y(n_5101)
);

OAI211xp5_ASAP7_75t_L g5102 ( 
.A1(n_5040),
.A2(n_1093),
.B(n_1089),
.C(n_1092),
.Y(n_5102)
);

A2O1A1Ixp33_ASAP7_75t_L g5103 ( 
.A1(n_5050),
.A2(n_1103),
.B(n_1110),
.C(n_1094),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_5038),
.Y(n_5104)
);

AOI222xp33_ASAP7_75t_L g5105 ( 
.A1(n_5073),
.A2(n_1097),
.B1(n_1100),
.B2(n_1095),
.C1(n_1096),
.C2(n_1099),
.Y(n_5105)
);

NOR2xp33_ASAP7_75t_L g5106 ( 
.A(n_5079),
.B(n_1100),
.Y(n_5106)
);

OAI221xp5_ASAP7_75t_L g5107 ( 
.A1(n_5069),
.A2(n_1104),
.B1(n_1101),
.B2(n_1102),
.C(n_1105),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5039),
.Y(n_5108)
);

NOR3xp33_ASAP7_75t_L g5109 ( 
.A(n_5044),
.B(n_1104),
.C(n_1107),
.Y(n_5109)
);

AOI22xp5_ASAP7_75t_L g5110 ( 
.A1(n_5054),
.A2(n_1110),
.B1(n_1108),
.B2(n_1109),
.Y(n_5110)
);

AOI21xp5_ASAP7_75t_L g5111 ( 
.A1(n_5047),
.A2(n_1112),
.B(n_1113),
.Y(n_5111)
);

AOI221xp5_ASAP7_75t_L g5112 ( 
.A1(n_5066),
.A2(n_1119),
.B1(n_1117),
.B2(n_1118),
.C(n_1120),
.Y(n_5112)
);

AOI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_5056),
.A2(n_5068),
.B(n_5070),
.Y(n_5113)
);

AND2x2_ASAP7_75t_L g5114 ( 
.A(n_5067),
.B(n_1127),
.Y(n_5114)
);

AOI222xp33_ASAP7_75t_L g5115 ( 
.A1(n_5060),
.A2(n_1129),
.B1(n_1131),
.B2(n_1127),
.C1(n_1128),
.C2(n_1130),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_5053),
.B(n_1132),
.Y(n_5116)
);

NAND4xp25_ASAP7_75t_L g5117 ( 
.A(n_5063),
.B(n_1137),
.C(n_1135),
.D(n_1136),
.Y(n_5117)
);

AOI22xp33_ASAP7_75t_L g5118 ( 
.A1(n_5046),
.A2(n_5049),
.B1(n_5072),
.B2(n_5064),
.Y(n_5118)
);

INVxp67_ASAP7_75t_SL g5119 ( 
.A(n_5051),
.Y(n_5119)
);

OAI22xp5_ASAP7_75t_L g5120 ( 
.A1(n_5059),
.A2(n_1140),
.B1(n_1138),
.B2(n_1139),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_5061),
.B(n_1141),
.Y(n_5121)
);

NOR2x1_ASAP7_75t_L g5122 ( 
.A(n_5048),
.B(n_1142),
.Y(n_5122)
);

AOI21xp5_ASAP7_75t_L g5123 ( 
.A1(n_5078),
.A2(n_1145),
.B(n_1146),
.Y(n_5123)
);

AOI221xp5_ASAP7_75t_L g5124 ( 
.A1(n_5075),
.A2(n_1149),
.B1(n_1147),
.B2(n_1148),
.C(n_1150),
.Y(n_5124)
);

A2O1A1Ixp33_ASAP7_75t_L g5125 ( 
.A1(n_5076),
.A2(n_1158),
.B(n_1166),
.C(n_1147),
.Y(n_5125)
);

AOI221xp5_ASAP7_75t_L g5126 ( 
.A1(n_5075),
.A2(n_1152),
.B1(n_1150),
.B2(n_1151),
.C(n_1153),
.Y(n_5126)
);

AOI221xp5_ASAP7_75t_L g5127 ( 
.A1(n_5075),
.A2(n_1162),
.B1(n_1160),
.B2(n_1161),
.C(n_1163),
.Y(n_5127)
);

O2A1O1Ixp33_ASAP7_75t_L g5128 ( 
.A1(n_5055),
.A2(n_1163),
.B(n_1161),
.C(n_1162),
.Y(n_5128)
);

A2O1A1Ixp33_ASAP7_75t_L g5129 ( 
.A1(n_5076),
.A2(n_1175),
.B(n_1184),
.C(n_1165),
.Y(n_5129)
);

OAI321xp33_ASAP7_75t_L g5130 ( 
.A1(n_5028),
.A2(n_1168),
.A3(n_1170),
.B1(n_1165),
.B2(n_1167),
.C(n_1169),
.Y(n_5130)
);

NOR2xp33_ASAP7_75t_L g5131 ( 
.A(n_5036),
.B(n_1171),
.Y(n_5131)
);

NOR2xp33_ASAP7_75t_L g5132 ( 
.A(n_5036),
.B(n_1172),
.Y(n_5132)
);

OAI21xp5_ASAP7_75t_SL g5133 ( 
.A1(n_5031),
.A2(n_1176),
.B(n_1177),
.Y(n_5133)
);

AOI221xp5_ASAP7_75t_L g5134 ( 
.A1(n_5075),
.A2(n_1187),
.B1(n_1185),
.B2(n_1186),
.C(n_1188),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_5036),
.B(n_1186),
.Y(n_5135)
);

AOI31xp33_ASAP7_75t_L g5136 ( 
.A1(n_5036),
.A2(n_1191),
.A3(n_1189),
.B(n_1190),
.Y(n_5136)
);

NOR2xp33_ASAP7_75t_L g5137 ( 
.A(n_5036),
.B(n_1192),
.Y(n_5137)
);

OAI32xp33_ASAP7_75t_L g5138 ( 
.A1(n_5074),
.A2(n_1195),
.A3(n_1197),
.B1(n_1194),
.B2(n_1196),
.Y(n_5138)
);

OAI221xp5_ASAP7_75t_L g5139 ( 
.A1(n_5052),
.A2(n_1196),
.B1(n_1193),
.B2(n_1194),
.C(n_1197),
.Y(n_5139)
);

AOI21xp33_ASAP7_75t_SL g5140 ( 
.A1(n_5036),
.A2(n_1201),
.B(n_1199),
.Y(n_5140)
);

AOI211xp5_ASAP7_75t_SL g5141 ( 
.A1(n_5030),
.A2(n_1204),
.B(n_1202),
.C(n_1203),
.Y(n_5141)
);

AOI221xp5_ASAP7_75t_L g5142 ( 
.A1(n_5075),
.A2(n_1206),
.B1(n_1203),
.B2(n_1205),
.C(n_1207),
.Y(n_5142)
);

INVx1_ASAP7_75t_SL g5143 ( 
.A(n_5036),
.Y(n_5143)
);

OAI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_5031),
.A2(n_1207),
.B1(n_1205),
.B2(n_1206),
.Y(n_5144)
);

OAI21xp5_ASAP7_75t_SL g5145 ( 
.A1(n_5133),
.A2(n_5143),
.B(n_5092),
.Y(n_5145)
);

OAI22xp33_ASAP7_75t_L g5146 ( 
.A1(n_5080),
.A2(n_1218),
.B1(n_1215),
.B2(n_1217),
.Y(n_5146)
);

AOI221xp5_ASAP7_75t_L g5147 ( 
.A1(n_5144),
.A2(n_1220),
.B1(n_1222),
.B2(n_1219),
.C(n_1221),
.Y(n_5147)
);

AOI21xp33_ASAP7_75t_L g5148 ( 
.A1(n_5085),
.A2(n_1224),
.B(n_1223),
.Y(n_5148)
);

AOI221xp5_ASAP7_75t_L g5149 ( 
.A1(n_5082),
.A2(n_1226),
.B1(n_1228),
.B2(n_1225),
.C(n_1227),
.Y(n_5149)
);

OAI211xp5_ASAP7_75t_SL g5150 ( 
.A1(n_5083),
.A2(n_1233),
.B(n_1231),
.C(n_1232),
.Y(n_5150)
);

OAI211xp5_ASAP7_75t_SL g5151 ( 
.A1(n_5118),
.A2(n_1234),
.B(n_1231),
.C(n_1232),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5135),
.Y(n_5152)
);

AOI21xp33_ASAP7_75t_L g5153 ( 
.A1(n_5099),
.A2(n_1237),
.B(n_1236),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_5141),
.B(n_1235),
.Y(n_5154)
);

AOI21xp5_ASAP7_75t_L g5155 ( 
.A1(n_5096),
.A2(n_1238),
.B(n_1240),
.Y(n_5155)
);

A2O1A1Ixp33_ASAP7_75t_SL g5156 ( 
.A1(n_5131),
.A2(n_1242),
.B(n_1240),
.C(n_1241),
.Y(n_5156)
);

AOI22xp5_ASAP7_75t_L g5157 ( 
.A1(n_5081),
.A2(n_1245),
.B1(n_1243),
.B2(n_1244),
.Y(n_5157)
);

NOR3xp33_ASAP7_75t_L g5158 ( 
.A(n_5139),
.B(n_1252),
.C(n_1245),
.Y(n_5158)
);

BUFx2_ASAP7_75t_L g5159 ( 
.A(n_5122),
.Y(n_5159)
);

A2O1A1Ixp33_ASAP7_75t_L g5160 ( 
.A1(n_5128),
.A2(n_1248),
.B(n_1249),
.C(n_1247),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_5132),
.B(n_1246),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_5137),
.B(n_1248),
.Y(n_5162)
);

INVx1_ASAP7_75t_SL g5163 ( 
.A(n_5114),
.Y(n_5163)
);

O2A1O1Ixp33_ASAP7_75t_L g5164 ( 
.A1(n_5136),
.A2(n_5103),
.B(n_5129),
.C(n_5125),
.Y(n_5164)
);

AOI322xp5_ASAP7_75t_L g5165 ( 
.A1(n_5101),
.A2(n_1258),
.A3(n_1257),
.B1(n_1254),
.B2(n_1250),
.C1(n_1251),
.C2(n_1255),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_5084),
.Y(n_5166)
);

OAI21xp5_ASAP7_75t_SL g5167 ( 
.A1(n_5102),
.A2(n_1259),
.B(n_1260),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5088),
.B(n_1263),
.Y(n_5168)
);

OAI32xp33_ASAP7_75t_L g5169 ( 
.A1(n_5104),
.A2(n_1266),
.A3(n_1263),
.B1(n_1265),
.B2(n_1267),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_5116),
.Y(n_5170)
);

AOI22xp33_ASAP7_75t_SL g5171 ( 
.A1(n_5108),
.A2(n_1271),
.B1(n_1269),
.B2(n_1270),
.Y(n_5171)
);

OAI221xp5_ASAP7_75t_L g5172 ( 
.A1(n_5094),
.A2(n_5126),
.B1(n_5134),
.B2(n_5127),
.C(n_5124),
.Y(n_5172)
);

AOI211x1_ASAP7_75t_L g5173 ( 
.A1(n_5097),
.A2(n_1275),
.B(n_1272),
.C(n_1274),
.Y(n_5173)
);

OAI211xp5_ASAP7_75t_L g5174 ( 
.A1(n_5142),
.A2(n_1276),
.B(n_1274),
.C(n_1275),
.Y(n_5174)
);

AOI211xp5_ASAP7_75t_SL g5175 ( 
.A1(n_5113),
.A2(n_1278),
.B(n_1276),
.C(n_1277),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_SL g5176 ( 
.A(n_5140),
.B(n_1277),
.Y(n_5176)
);

OAI22xp5_ASAP7_75t_L g5177 ( 
.A1(n_5107),
.A2(n_1284),
.B1(n_1280),
.B2(n_1281),
.Y(n_5177)
);

AOI22xp5_ASAP7_75t_L g5178 ( 
.A1(n_5106),
.A2(n_1295),
.B1(n_1292),
.B2(n_1294),
.Y(n_5178)
);

NAND3x1_ASAP7_75t_L g5179 ( 
.A(n_5100),
.B(n_1295),
.C(n_1296),
.Y(n_5179)
);

OAI21xp33_ASAP7_75t_SL g5180 ( 
.A1(n_5119),
.A2(n_1297),
.B(n_1298),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_5121),
.Y(n_5181)
);

OAI311xp33_ASAP7_75t_L g5182 ( 
.A1(n_5087),
.A2(n_1301),
.A3(n_1299),
.B1(n_1300),
.C1(n_1302),
.Y(n_5182)
);

A2O1A1Ixp33_ASAP7_75t_L g5183 ( 
.A1(n_5090),
.A2(n_1304),
.B(n_1305),
.C(n_1303),
.Y(n_5183)
);

O2A1O1Ixp33_ASAP7_75t_L g5184 ( 
.A1(n_5156),
.A2(n_5138),
.B(n_5130),
.C(n_5091),
.Y(n_5184)
);

AOI211xp5_ASAP7_75t_SL g5185 ( 
.A1(n_5148),
.A2(n_5111),
.B(n_5098),
.C(n_5123),
.Y(n_5185)
);

AOI21xp33_ASAP7_75t_L g5186 ( 
.A1(n_5166),
.A2(n_5105),
.B(n_5089),
.Y(n_5186)
);

O2A1O1Ixp33_ASAP7_75t_L g5187 ( 
.A1(n_5182),
.A2(n_5109),
.B(n_5086),
.C(n_5120),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_5159),
.Y(n_5188)
);

AO22x2_ASAP7_75t_L g5189 ( 
.A1(n_5173),
.A2(n_5117),
.B1(n_5115),
.B2(n_5112),
.Y(n_5189)
);

NAND2xp5_ASAP7_75t_L g5190 ( 
.A(n_5175),
.B(n_5110),
.Y(n_5190)
);

OAI211xp5_ASAP7_75t_SL g5191 ( 
.A1(n_5145),
.A2(n_5095),
.B(n_5093),
.C(n_1304),
.Y(n_5191)
);

INVx2_ASAP7_75t_L g5192 ( 
.A(n_5168),
.Y(n_5192)
);

AOI221xp5_ASAP7_75t_L g5193 ( 
.A1(n_5164),
.A2(n_1309),
.B1(n_1306),
.B2(n_1307),
.C(n_1310),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_5154),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5161),
.Y(n_5195)
);

O2A1O1Ixp33_ASAP7_75t_L g5196 ( 
.A1(n_5183),
.A2(n_1315),
.B(n_1312),
.C(n_1314),
.Y(n_5196)
);

AOI21xp5_ASAP7_75t_L g5197 ( 
.A1(n_5176),
.A2(n_1316),
.B(n_1318),
.Y(n_5197)
);

AOI322xp5_ASAP7_75t_L g5198 ( 
.A1(n_5149),
.A2(n_1324),
.A3(n_1323),
.B1(n_1320),
.B2(n_1316),
.C1(n_1319),
.C2(n_1322),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_5162),
.Y(n_5199)
);

INVx1_ASAP7_75t_SL g5200 ( 
.A(n_5163),
.Y(n_5200)
);

AOI22xp5_ASAP7_75t_L g5201 ( 
.A1(n_5158),
.A2(n_1539),
.B1(n_1541),
.B2(n_1538),
.Y(n_5201)
);

AOI221xp5_ASAP7_75t_L g5202 ( 
.A1(n_5172),
.A2(n_1327),
.B1(n_1325),
.B2(n_1326),
.C(n_1328),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5179),
.Y(n_5203)
);

OAI22xp5_ASAP7_75t_L g5204 ( 
.A1(n_5157),
.A2(n_1329),
.B1(n_1325),
.B2(n_1326),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_5165),
.B(n_5171),
.Y(n_5205)
);

AOI222xp33_ASAP7_75t_L g5206 ( 
.A1(n_5167),
.A2(n_1331),
.B1(n_1333),
.B2(n_1329),
.C1(n_1330),
.C2(n_1332),
.Y(n_5206)
);

OAI32xp33_ASAP7_75t_L g5207 ( 
.A1(n_5180),
.A2(n_1334),
.A3(n_1330),
.B1(n_1332),
.B2(n_1335),
.Y(n_5207)
);

O2A1O1Ixp33_ASAP7_75t_L g5208 ( 
.A1(n_5160),
.A2(n_1340),
.B(n_1338),
.C(n_1339),
.Y(n_5208)
);

XOR2xp5_ASAP7_75t_L g5209 ( 
.A(n_5177),
.B(n_5178),
.Y(n_5209)
);

NAND2xp5_ASAP7_75t_L g5210 ( 
.A(n_5146),
.B(n_1341),
.Y(n_5210)
);

AOI22xp5_ASAP7_75t_L g5211 ( 
.A1(n_5151),
.A2(n_1345),
.B1(n_1343),
.B2(n_1344),
.Y(n_5211)
);

OAI211xp5_ASAP7_75t_L g5212 ( 
.A1(n_5186),
.A2(n_5174),
.B(n_5147),
.C(n_5155),
.Y(n_5212)
);

O2A1O1Ixp33_ASAP7_75t_L g5213 ( 
.A1(n_5207),
.A2(n_5150),
.B(n_5169),
.C(n_5153),
.Y(n_5213)
);

OAI22xp5_ASAP7_75t_L g5214 ( 
.A1(n_5211),
.A2(n_5152),
.B1(n_5181),
.B2(n_5170),
.Y(n_5214)
);

XNOR2x1_ASAP7_75t_L g5215 ( 
.A(n_5200),
.B(n_1346),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_5203),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_5210),
.Y(n_5217)
);

OAI22xp5_ASAP7_75t_L g5218 ( 
.A1(n_5201),
.A2(n_1351),
.B1(n_1349),
.B2(n_1350),
.Y(n_5218)
);

AOI211x1_ASAP7_75t_SL g5219 ( 
.A1(n_5191),
.A2(n_1351),
.B(n_1349),
.C(n_1350),
.Y(n_5219)
);

OAI211xp5_ASAP7_75t_SL g5220 ( 
.A1(n_5185),
.A2(n_1357),
.B(n_1354),
.C(n_1356),
.Y(n_5220)
);

OAI21xp5_ASAP7_75t_SL g5221 ( 
.A1(n_5184),
.A2(n_1358),
.B(n_1359),
.Y(n_5221)
);

NAND2xp33_ASAP7_75t_SL g5222 ( 
.A(n_5190),
.B(n_1360),
.Y(n_5222)
);

OAI32xp33_ASAP7_75t_L g5223 ( 
.A1(n_5188),
.A2(n_1364),
.A3(n_1362),
.B1(n_1363),
.B2(n_1365),
.Y(n_5223)
);

AOI22xp5_ASAP7_75t_L g5224 ( 
.A1(n_5189),
.A2(n_1365),
.B1(n_1363),
.B2(n_1364),
.Y(n_5224)
);

INVx2_ASAP7_75t_SL g5225 ( 
.A(n_5192),
.Y(n_5225)
);

AOI22xp5_ASAP7_75t_L g5226 ( 
.A1(n_5189),
.A2(n_1368),
.B1(n_1366),
.B2(n_1367),
.Y(n_5226)
);

AOI22xp33_ASAP7_75t_L g5227 ( 
.A1(n_5194),
.A2(n_1371),
.B1(n_1369),
.B2(n_1370),
.Y(n_5227)
);

O2A1O1Ixp33_ASAP7_75t_L g5228 ( 
.A1(n_5196),
.A2(n_1372),
.B(n_1370),
.C(n_1371),
.Y(n_5228)
);

AOI22xp5_ASAP7_75t_L g5229 ( 
.A1(n_5225),
.A2(n_5205),
.B1(n_5209),
.B2(n_5206),
.Y(n_5229)
);

HB1xp67_ASAP7_75t_L g5230 ( 
.A(n_5215),
.Y(n_5230)
);

NOR2x1_ASAP7_75t_L g5231 ( 
.A(n_5221),
.B(n_5195),
.Y(n_5231)
);

NOR2x1_ASAP7_75t_L g5232 ( 
.A(n_5220),
.B(n_5199),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5224),
.Y(n_5233)
);

AOI22xp5_ASAP7_75t_L g5234 ( 
.A1(n_5216),
.A2(n_5212),
.B1(n_5222),
.B2(n_5214),
.Y(n_5234)
);

NOR2xp67_ASAP7_75t_L g5235 ( 
.A(n_5226),
.B(n_5197),
.Y(n_5235)
);

AOI22xp33_ASAP7_75t_L g5236 ( 
.A1(n_5217),
.A2(n_5204),
.B1(n_5202),
.B2(n_5193),
.Y(n_5236)
);

OR3x1_ASAP7_75t_L g5237 ( 
.A(n_5223),
.B(n_5187),
.C(n_5208),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_5219),
.B(n_5198),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5230),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_5237),
.Y(n_5240)
);

INVxp67_ASAP7_75t_SL g5241 ( 
.A(n_5232),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_5233),
.Y(n_5242)
);

CKINVDCx20_ASAP7_75t_R g5243 ( 
.A(n_5229),
.Y(n_5243)
);

AND2x4_ASAP7_75t_L g5244 ( 
.A(n_5231),
.B(n_5227),
.Y(n_5244)
);

XOR2x1_ASAP7_75t_L g5245 ( 
.A(n_5234),
.B(n_5218),
.Y(n_5245)
);

AOI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_5241),
.A2(n_5228),
.B(n_5238),
.Y(n_5246)
);

OAI22xp5_ASAP7_75t_L g5247 ( 
.A1(n_5243),
.A2(n_5236),
.B1(n_5235),
.B2(n_5213),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_5245),
.Y(n_5248)
);

AOI221x1_ASAP7_75t_L g5249 ( 
.A1(n_5240),
.A2(n_1381),
.B1(n_1377),
.B2(n_1380),
.C(n_1382),
.Y(n_5249)
);

AOI221xp5_ASAP7_75t_L g5250 ( 
.A1(n_5242),
.A2(n_1385),
.B1(n_1383),
.B2(n_1384),
.C(n_1386),
.Y(n_5250)
);

XNOR2xp5_ASAP7_75t_L g5251 ( 
.A(n_5247),
.B(n_5239),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_5248),
.Y(n_5252)
);

AOI21xp5_ASAP7_75t_L g5253 ( 
.A1(n_5251),
.A2(n_5246),
.B(n_5244),
.Y(n_5253)
);

INVx2_ASAP7_75t_L g5254 ( 
.A(n_5252),
.Y(n_5254)
);

BUFx2_ASAP7_75t_L g5255 ( 
.A(n_5254),
.Y(n_5255)
);

INVx4_ASAP7_75t_L g5256 ( 
.A(n_5255),
.Y(n_5256)
);

OAI22xp33_ASAP7_75t_L g5257 ( 
.A1(n_5256),
.A2(n_5253),
.B1(n_5249),
.B2(n_5250),
.Y(n_5257)
);

OAI21x1_ASAP7_75t_L g5258 ( 
.A1(n_5257),
.A2(n_1385),
.B(n_1387),
.Y(n_5258)
);

NAND2x1p5_ASAP7_75t_L g5259 ( 
.A(n_5258),
.B(n_1387),
.Y(n_5259)
);

AOI22xp33_ASAP7_75t_L g5260 ( 
.A1(n_5259),
.A2(n_1390),
.B1(n_1388),
.B2(n_1389),
.Y(n_5260)
);

AOI22xp5_ASAP7_75t_L g5261 ( 
.A1(n_5260),
.A2(n_1395),
.B1(n_1393),
.B2(n_1394),
.Y(n_5261)
);

OR2x2_ASAP7_75t_L g5262 ( 
.A(n_5261),
.B(n_1396),
.Y(n_5262)
);

A2O1A1Ixp33_ASAP7_75t_L g5263 ( 
.A1(n_5262),
.A2(n_1399),
.B(n_1397),
.C(n_1398),
.Y(n_5263)
);

AOI211xp5_ASAP7_75t_L g5264 ( 
.A1(n_5263),
.A2(n_1545),
.B(n_1401),
.C(n_1400),
.Y(n_5264)
);


endmodule