module fake_jpeg_31705_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_52),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_54),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_0),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_0),
.C(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_50),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_50),
.B1(n_54),
.B2(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_53),
.B1(n_40),
.B2(n_51),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_53),
.B1(n_49),
.B2(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_45),
.B1(n_52),
.B2(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_3),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_2),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_39),
.B(n_22),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_95),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_4),
.B1(n_8),
.B2(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_89),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_13),
.C(n_14),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_29),
.C(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_36),
.Y(n_110)
);

AOI21x1_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_27),
.B(n_28),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_108),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_32),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_97),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_116),
.B(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_96),
.C(n_106),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_113),
.C(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_118),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_104),
.Y(n_124)
);


endmodule