module fake_jpeg_18098_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_68),
.B(n_86),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_17),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_78),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_14),
.B(n_15),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_35),
.B(n_43),
.C(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_74),
.B(n_76),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_80),
.B1(n_92),
.B2(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_33),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_26),
.B(n_28),
.C(n_22),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_32),
.B1(n_22),
.B2(n_34),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_88),
.B1(n_94),
.B2(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_32),
.B1(n_34),
.B2(n_22),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_48),
.C(n_41),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_32),
.B1(n_22),
.B2(n_34),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_42),
.B1(n_44),
.B2(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_28),
.B1(n_33),
.B2(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_96),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_44),
.A3(n_41),
.B1(n_46),
.B2(n_28),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_47),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_101)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_68),
.B1(n_7),
.B2(n_15),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_30),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_112),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_21),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_18),
.B1(n_20),
.B2(n_36),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_36),
.B1(n_27),
.B2(n_21),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_125),
.Y(n_143)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_116),
.A2(n_70),
.B1(n_29),
.B2(n_21),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_29),
.B1(n_40),
.B2(n_47),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_86),
.B(n_70),
.C(n_99),
.Y(n_148)
);

BUFx2_ASAP7_75t_SL g120 ( 
.A(n_81),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_36),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_36),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_36),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_83),
.B1(n_95),
.B2(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_40),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_105),
.B(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_89),
.B1(n_77),
.B2(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_147),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_92),
.C(n_72),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_115),
.B(n_113),
.C(n_117),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_93),
.B1(n_87),
.B2(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_158),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_87),
.B1(n_85),
.B2(n_72),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_155),
.B1(n_116),
.B2(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_110),
.C(n_123),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_107),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_21),
.B1(n_27),
.B2(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_108),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_164),
.A2(n_167),
.B(n_173),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_170),
.Y(n_205)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_171),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_153),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_140),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_144),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_123),
.B1(n_109),
.B2(n_125),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_176),
.B1(n_183),
.B2(n_146),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_118),
.B(n_117),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_118),
.B(n_128),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_189),
.B(n_27),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_124),
.B1(n_119),
.B2(n_129),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_148),
.B1(n_137),
.B2(n_149),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_119),
.B1(n_129),
.B2(n_108),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_29),
.B(n_27),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_148),
.B(n_156),
.Y(n_196)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_30),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_159),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_148),
.A2(n_132),
.B(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_167),
.A2(n_178),
.B1(n_184),
.B2(n_192),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_197),
.B1(n_224),
.B2(n_199),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_162),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_194),
.B(n_202),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_153),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_25),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_198),
.A2(n_191),
.B1(n_182),
.B2(n_170),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_208),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_164),
.C(n_168),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_207),
.C(n_209),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_182),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_134),
.B1(n_160),
.B2(n_135),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_213),
.B(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_132),
.C(n_135),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_154),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_132),
.C(n_107),
.Y(n_209)
);

AOI32xp33_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_154),
.A3(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_175),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_0),
.B(n_1),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_30),
.Y(n_217)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_179),
.A2(n_176),
.B1(n_183),
.B2(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_177),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_169),
.B(n_163),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_246),
.B(n_216),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_228),
.A2(n_240),
.B1(n_211),
.B2(n_2),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_222),
.B(n_196),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_193),
.B(n_195),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_218),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_243),
.C(n_244),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_204),
.B1(n_218),
.B2(n_217),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_175),
.B1(n_166),
.B2(n_171),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_198),
.A2(n_186),
.B1(n_25),
.B2(n_24),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_25),
.B1(n_24),
.B2(n_8),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_240),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_242),
.B(n_248),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_7),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_200),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_261),
.B1(n_264),
.B2(n_267),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_262),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_237),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_10),
.B1(n_9),
.B2(n_3),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_201),
.B(n_206),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_3),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_223),
.B(n_224),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_211),
.B(n_220),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_246),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_266),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_229),
.B1(n_245),
.B2(n_243),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_235),
.B(n_9),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_269),
.B(n_5),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_236),
.A2(n_9),
.B(n_15),
.C(n_13),
.D(n_12),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_4),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_231),
.B1(n_228),
.B2(n_234),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_272),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_275),
.B(n_265),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_245),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_282),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_229),
.B1(n_235),
.B2(n_232),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_244),
.B1(n_16),
.B2(n_12),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_10),
.C(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_289),
.C(n_251),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_1),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_284),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_268),
.Y(n_299)
);

OAI21x1_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_288),
.B(n_270),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_6),
.C(n_4),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_260),
.C(n_262),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_299),
.Y(n_307)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

XNOR2x2_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_255),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_297),
.A2(n_271),
.B1(n_283),
.B2(n_286),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_281),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_275),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_258),
.C(n_261),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_295),
.C(n_293),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_288),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_297),
.A2(n_252),
.B(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_312),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_272),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_316),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_292),
.B(n_252),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_286),
.B1(n_278),
.B2(n_253),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_299),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_303),
.C(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_321),
.C(n_316),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_294),
.C(n_296),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_324),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_307),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_330),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_253),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_334),
.B(n_322),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_319),
.B(n_321),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_332),
.B(n_301),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_335),
.B(n_336),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_266),
.B(n_312),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_269),
.B(n_298),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_313),
.B(n_285),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_5),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_6),
.B(n_250),
.Y(n_345)
);


endmodule