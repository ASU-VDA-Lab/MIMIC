module real_aes_17263_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_635;
wire n_357;
wire n_673;
wire n_386;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_889;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_602;
wire n_139;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_0), .Y(n_222) );
AND2x4_ASAP7_75t_L g109 ( .A(n_1), .B(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g153 ( .A(n_2), .Y(n_153) );
INVx1_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_4), .B(n_162), .Y(n_161) );
OR2x2_ASAP7_75t_L g117 ( .A(n_5), .B(n_21), .Y(n_117) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_6), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_7), .A2(n_52), .B1(n_528), .B2(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_7), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_8), .B(n_142), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_9), .B(n_142), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_10), .B(n_190), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_11), .A2(n_82), .B1(n_142), .B2(n_144), .Y(n_241) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_12), .A2(n_35), .B(n_136), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_13), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_13), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_14), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_15), .B(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g639 ( .A(n_16), .Y(n_639) );
AO32x2_ASAP7_75t_L g238 ( .A1(n_17), .A2(n_133), .A3(n_134), .B1(n_239), .B2(n_242), .Y(n_238) );
AO32x1_ASAP7_75t_L g260 ( .A1(n_17), .A2(n_133), .A3(n_134), .B1(n_239), .B2(n_242), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_18), .B(n_602), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_19), .B(n_133), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_20), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_22), .A2(n_41), .B1(n_149), .B2(n_180), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_23), .A2(n_90), .B1(n_144), .B2(n_150), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_24), .B(n_164), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_25), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_26), .B(n_197), .Y(n_251) );
OAI211xp5_ASAP7_75t_L g120 ( .A1(n_27), .A2(n_121), .B(n_497), .C(n_503), .Y(n_120) );
INVx1_ASAP7_75t_L g507 ( .A(n_27), .Y(n_507) );
OAI31xp33_ASAP7_75t_SL g509 ( .A1(n_27), .A2(n_506), .A3(n_507), .B(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_27), .A2(n_122), .B1(n_507), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_28), .A2(n_64), .B1(n_150), .B2(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_29), .B(n_142), .Y(n_591) );
INVx2_ASAP7_75t_L g511 ( .A(n_30), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_31), .B(n_146), .Y(n_612) );
INVx1_ASAP7_75t_L g115 ( .A(n_32), .Y(n_115) );
BUFx3_ASAP7_75t_L g523 ( .A(n_32), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_33), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_34), .B(n_569), .Y(n_618) );
AND2x2_ASAP7_75t_L g644 ( .A(n_36), .B(n_569), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_37), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_38), .B(n_196), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_39), .B(n_602), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_40), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_42), .B(n_581), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_43), .A2(n_77), .B1(n_196), .B2(n_197), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_44), .B(n_231), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_45), .A2(n_181), .B(n_220), .C(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_46), .A2(n_79), .B1(n_142), .B2(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g136 ( .A(n_47), .Y(n_136) );
AND2x4_ASAP7_75t_L g138 ( .A(n_48), .B(n_139), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_49), .A2(n_51), .B1(n_149), .B2(n_150), .Y(n_604) );
AOI22xp5_ASAP7_75t_SL g515 ( .A1(n_50), .A2(n_92), .B1(n_516), .B2(n_517), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_50), .Y(n_516) );
INVxp67_ASAP7_75t_SL g529 ( .A(n_52), .Y(n_529) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_53), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_53), .B(n_133), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_54), .B(n_569), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_55), .Y(n_643) );
CKINVDCx14_ASAP7_75t_R g894 ( .A(n_56), .Y(n_894) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_57), .B(n_150), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_58), .B(n_144), .Y(n_160) );
INVx1_ASAP7_75t_L g139 ( .A(n_59), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_60), .B(n_133), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_61), .A2(n_220), .B(n_221), .C(n_223), .Y(n_219) );
INVx1_ASAP7_75t_SL g498 ( .A(n_62), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g168 ( .A(n_63), .B(n_144), .C(n_166), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_65), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_66), .B(n_133), .Y(n_595) );
AND2x2_ASAP7_75t_L g225 ( .A(n_67), .B(n_226), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_68), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_69), .B(n_550), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_70), .B(n_146), .C(n_180), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_71), .A2(n_94), .B1(n_142), .B2(n_196), .Y(n_200) );
INVx2_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_73), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_74), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_75), .B(n_199), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_76), .B(n_142), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_78), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_80), .B(n_184), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_81), .A2(n_89), .B1(n_601), .B2(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_83), .B(n_142), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_84), .B(n_166), .Y(n_165) );
NAND2xp33_ASAP7_75t_SL g567 ( .A(n_85), .B(n_162), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_86), .B(n_178), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_87), .A2(n_102), .B1(n_149), .B2(n_150), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_88), .B(n_197), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_91), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g535 ( .A(n_91), .Y(n_535) );
INVx1_ASAP7_75t_L g517 ( .A(n_92), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_93), .B(n_190), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_95), .Y(n_897) );
NAND2xp33_ASAP7_75t_L g551 ( .A(n_96), .B(n_162), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_97), .B(n_569), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_98), .B(n_162), .C(n_199), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_99), .B(n_550), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_100), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_101), .B(n_602), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_118), .B(n_904), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx2_ASAP7_75t_SL g917 ( .A(n_109), .Y(n_917) );
AND2x2_ASAP7_75t_L g510 ( .A(n_111), .B(n_511), .Y(n_510) );
INVx5_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx4_ASAP7_75t_L g896 ( .A(n_112), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_112), .Y(n_911) );
INVx3_ASAP7_75t_L g918 ( .A(n_112), .Y(n_918) );
AND2x6_ASAP7_75t_SL g112 ( .A(n_113), .B(n_116), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_116), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2x1_ASAP7_75t_L g903 ( .A(n_117), .B(n_523), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_512), .C(n_889), .Y(n_118) );
NAND3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_504), .C(n_508), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_122), .B(n_506), .Y(n_505) );
AOI31xp33_ASAP7_75t_L g508 ( .A1(n_122), .A2(n_506), .A3(n_507), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g908 ( .A(n_122), .Y(n_908) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp33_ASAP7_75t_R g503 ( .A(n_123), .B(n_497), .Y(n_503) );
OAI22x1_ASAP7_75t_L g530 ( .A1(n_123), .A2(n_531), .B1(n_536), .B2(n_887), .Y(n_530) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_398), .Y(n_123) );
AND4x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_320), .C(n_353), .D(n_384), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_287), .Y(n_125) );
OAI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_206), .B1(n_255), .B2(n_265), .C(n_274), .Y(n_126) );
AOI21xp33_ASAP7_75t_L g392 ( .A1(n_127), .A2(n_377), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_170), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_154), .Y(n_129) );
INVx2_ASAP7_75t_L g273 ( .A(n_130), .Y(n_273) );
AND2x2_ASAP7_75t_L g283 ( .A(n_130), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g319 ( .A(n_130), .B(n_192), .Y(n_319) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g308 ( .A(n_131), .Y(n_308) );
AOI31xp67_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_137), .A3(n_140), .B(n_151), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_134), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
BUFx3_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_134), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_SL g245 ( .A(n_134), .Y(n_245) );
AND2x4_ASAP7_75t_SL g556 ( .A(n_134), .B(n_137), .Y(n_556) );
INVx1_ASAP7_75t_SL g560 ( .A(n_134), .Y(n_560) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g157 ( .A(n_135), .Y(n_157) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_137), .A2(n_159), .B(n_163), .Y(n_158) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_137), .A2(n_175), .B(n_182), .Y(n_174) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_137), .A2(n_562), .B(n_565), .Y(n_561) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_137), .A2(n_575), .B(n_578), .Y(n_574) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_137), .A2(n_589), .B(n_592), .Y(n_588) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_137), .A2(n_611), .B(n_614), .Y(n_610) );
OAI21x1_ASAP7_75t_L g667 ( .A1(n_137), .A2(n_668), .B(n_671), .Y(n_667) );
BUFx10_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g202 ( .A(n_138), .Y(n_202) );
INVx1_ASAP7_75t_L g224 ( .A(n_138), .Y(n_224) );
AO31x2_ASAP7_75t_L g228 ( .A1(n_138), .A2(n_193), .A3(n_229), .B(n_234), .Y(n_228) );
BUFx10_ASAP7_75t_L g606 ( .A(n_138), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B1(n_146), .B2(n_148), .Y(n_140) );
INVx3_ASAP7_75t_L g253 ( .A(n_142), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_142), .A2(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g617 ( .A(n_142), .Y(n_617) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_143), .Y(n_144) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_143), .Y(n_150) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
INVx1_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVx1_ASAP7_75t_L g196 ( .A(n_143), .Y(n_196) );
INVx1_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
INVx3_ASAP7_75t_L g550 ( .A(n_143), .Y(n_550) );
INVx1_ASAP7_75t_L g603 ( .A(n_143), .Y(n_603) );
INVx2_ASAP7_75t_SL g197 ( .A(n_144), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_144), .B(n_639), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_145), .A2(n_195), .B1(n_198), .B2(n_200), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_145), .A2(n_230), .B1(n_232), .B2(n_233), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_145), .A2(n_251), .B(n_252), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_145), .A2(n_600), .B1(n_604), .B2(n_605), .Y(n_599) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_146), .A2(n_160), .B(n_161), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_146), .A2(n_181), .B1(n_240), .B2(n_241), .Y(n_239) );
O2A1O1Ixp5_ASAP7_75t_L g575 ( .A1(n_146), .A2(n_177), .B(n_576), .C(n_577), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_146), .A2(n_593), .B(n_594), .Y(n_592) );
BUFx8_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
INVx2_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
INVx1_ASAP7_75t_L g199 ( .A(n_147), .Y(n_199) );
INVx1_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_149), .A2(n_180), .B1(n_216), .B2(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
INVx2_ASAP7_75t_L g601 ( .A(n_150), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_150), .A2(n_612), .B(n_613), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_150), .A2(n_550), .B1(n_642), .B2(n_643), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g294 ( .A(n_154), .B(n_284), .Y(n_294) );
OR2x2_ASAP7_75t_L g403 ( .A(n_154), .B(n_172), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B(n_169), .Y(n_154) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_155), .A2(n_158), .B(n_169), .Y(n_272) );
OAI21x1_ASAP7_75t_L g573 ( .A1(n_155), .A2(n_574), .B(n_582), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_155), .A2(n_574), .B(n_582), .Y(n_655) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_155), .A2(n_667), .B(n_674), .Y(n_666) );
OAI21xp33_ASAP7_75t_SL g692 ( .A1(n_155), .A2(n_667), .B(n_674), .Y(n_692) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g569 ( .A(n_156), .Y(n_569) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
INVx2_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
INVx2_ASAP7_75t_L g581 ( .A(n_162), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_168), .Y(n_163) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_167), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_170), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_192), .Y(n_171) );
INVx1_ASAP7_75t_L g268 ( .A(n_172), .Y(n_268) );
INVx2_ASAP7_75t_SL g345 ( .A(n_172), .Y(n_345) );
BUFx2_ASAP7_75t_L g375 ( .A(n_172), .Y(n_375) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_189), .Y(n_172) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_173), .A2(n_174), .B(n_189), .Y(n_284) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_173), .A2(n_588), .B(n_595), .Y(n_587) );
OA21x2_ASAP7_75t_L g609 ( .A1(n_173), .A2(n_610), .B(n_618), .Y(n_609) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_173), .A2(n_588), .B(n_595), .Y(n_625) );
OAI21x1_ASAP7_75t_L g654 ( .A1(n_173), .A2(n_610), .B(n_618), .Y(n_654) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_179), .C(n_181), .Y(n_175) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g231 ( .A(n_180), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_181), .A2(n_549), .B(n_551), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_181), .A2(n_566), .B(n_567), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_181), .A2(n_590), .B(n_591), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_181), .A2(n_669), .B(n_670), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B1(n_187), .B2(n_188), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_184), .A2(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_185), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_552) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx3_ASAP7_75t_L g223 ( .A(n_186), .Y(n_223) );
INVx2_ASAP7_75t_L g212 ( .A(n_190), .Y(n_212) );
NOR2xp67_ASAP7_75t_SL g634 ( .A(n_190), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AO31x2_ASAP7_75t_L g598 ( .A1(n_191), .A2(n_599), .A3(n_606), .B(n_607), .Y(n_598) );
AND2x2_ASAP7_75t_L g267 ( .A(n_192), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g286 ( .A(n_192), .Y(n_286) );
OR2x2_ASAP7_75t_L g306 ( .A(n_192), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g347 ( .A(n_192), .Y(n_347) );
INVx1_ASAP7_75t_L g358 ( .A(n_192), .Y(n_358) );
AND2x2_ASAP7_75t_L g365 ( .A(n_192), .B(n_307), .Y(n_365) );
AO31x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .A3(n_201), .B(n_203), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_196), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g218 ( .A(n_199), .Y(n_218) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_SL g242 ( .A(n_202), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx2_ASAP7_75t_L g226 ( .A(n_205), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_205), .B(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_208), .B(n_236), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_227), .Y(n_208) );
INVx1_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_210), .Y(n_291) );
INVx1_ASAP7_75t_L g300 ( .A(n_210), .Y(n_300) );
INVx1_ASAP7_75t_L g339 ( .A(n_210), .Y(n_339) );
AND2x2_ASAP7_75t_L g369 ( .A(n_210), .B(n_228), .Y(n_369) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g263 ( .A(n_211), .Y(n_263) );
AOI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_225), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_219), .B(n_224), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_215), .B(n_218), .Y(n_214) );
AOI21x1_ASAP7_75t_L g614 ( .A1(n_218), .A2(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g554 ( .A(n_220), .Y(n_554) );
INVx2_ASAP7_75t_L g233 ( .A(n_223), .Y(n_233) );
INVx2_ASAP7_75t_L g605 ( .A(n_223), .Y(n_605) );
INVx1_ASAP7_75t_L g275 ( .A(n_227), .Y(n_275) );
AND2x4_ASAP7_75t_L g324 ( .A(n_227), .B(n_238), .Y(n_324) );
AND2x2_ASAP7_75t_L g334 ( .A(n_227), .B(n_263), .Y(n_334) );
INVx1_ASAP7_75t_L g395 ( .A(n_227), .Y(n_395) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g281 ( .A(n_228), .B(n_260), .Y(n_281) );
AND2x2_ASAP7_75t_L g299 ( .A(n_228), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g315 ( .A(n_228), .B(n_260), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_228), .B(n_243), .Y(n_424) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_233), .A2(n_248), .B(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_233), .A2(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_236), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
OR2x2_ASAP7_75t_L g441 ( .A(n_237), .B(n_243), .Y(n_441) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g388 ( .A(n_238), .Y(n_388) );
AND2x2_ASAP7_75t_L g413 ( .A(n_238), .B(n_243), .Y(n_413) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_242), .A2(n_247), .B(n_250), .Y(n_246) );
INVx3_ASAP7_75t_L g264 ( .A(n_243), .Y(n_264) );
AND2x2_ASAP7_75t_L g290 ( .A(n_243), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g312 ( .A(n_243), .Y(n_312) );
INVx1_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
INVx1_ASAP7_75t_L g336 ( .A(n_243), .Y(n_336) );
BUFx2_ASAP7_75t_L g431 ( .A(n_243), .Y(n_431) );
OR2x2_ASAP7_75t_L g459 ( .A(n_243), .B(n_263), .Y(n_459) );
INVxp67_ASAP7_75t_L g476 ( .A(n_243), .Y(n_476) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_254), .Y(n_244) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_261), .Y(n_256) );
AND2x4_ASAP7_75t_L g289 ( .A(n_257), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_257), .B(n_369), .Y(n_450) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g277 ( .A(n_259), .B(n_264), .Y(n_277) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_259), .Y(n_301) );
INVx1_ASAP7_75t_L g425 ( .A(n_259), .Y(n_425) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g338 ( .A(n_260), .Y(n_338) );
AND2x2_ASAP7_75t_L g352 ( .A(n_261), .B(n_315), .Y(n_352) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g314 ( .A(n_263), .Y(n_314) );
OR2x2_ASAP7_75t_L g372 ( .A(n_263), .B(n_338), .Y(n_372) );
INVx1_ASAP7_75t_L g435 ( .A(n_263), .Y(n_435) );
AND2x2_ASAP7_75t_L g378 ( .A(n_264), .B(n_324), .Y(n_378) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
AND2x2_ASAP7_75t_L g381 ( .A(n_267), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
AND2x2_ASAP7_75t_L g285 ( .A(n_270), .B(n_286), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_270), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g304 ( .A(n_271), .Y(n_304) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g383 ( .A(n_272), .B(n_308), .Y(n_383) );
AND2x2_ASAP7_75t_L g346 ( .A(n_273), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g417 ( .A(n_273), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_278), .C(n_282), .Y(n_274) );
INVx1_ASAP7_75t_L g409 ( .A(n_276), .Y(n_409) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g405 ( .A(n_277), .B(n_369), .Y(n_405) );
INVx1_ASAP7_75t_L g496 ( .A(n_277), .Y(n_496) );
INVx1_ASAP7_75t_L g461 ( .A(n_278), .Y(n_461) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g494 ( .A(n_279), .B(n_413), .Y(n_494) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g311 ( .A(n_281), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g466 ( .A(n_281), .B(n_431), .Y(n_466) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVxp67_ASAP7_75t_L g356 ( .A(n_283), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_283), .B(n_318), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_283), .B(n_285), .Y(n_448) );
INVx1_ASAP7_75t_L g331 ( .A(n_284), .Y(n_331) );
INVx2_ASAP7_75t_SL g296 ( .A(n_286), .Y(n_296) );
OR2x2_ASAP7_75t_L g325 ( .A(n_286), .B(n_326), .Y(n_325) );
OAI221xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B1(n_297), .B2(n_302), .C(n_309), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_289), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g361 ( .A(n_291), .Y(n_361) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g418 ( .A(n_294), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_294), .B(n_296), .Y(n_456) );
OR2x2_ASAP7_75t_L g438 ( .A(n_295), .B(n_428), .Y(n_438) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g407 ( .A(n_296), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g454 ( .A(n_296), .B(n_383), .Y(n_454) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g389 ( .A(n_299), .B(n_312), .Y(n_389) );
BUFx2_ASAP7_75t_L g415 ( .A(n_299), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_303), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g391 ( .A(n_306), .Y(n_391) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .B(n_316), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g368 ( .A(n_312), .Y(n_368) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_312), .Y(n_371) );
OR2x2_ASAP7_75t_L g481 ( .A(n_312), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g442 ( .A(n_313), .Y(n_442) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g350 ( .A(n_314), .Y(n_350) );
AND2x2_ASAP7_75t_L g477 ( .A(n_315), .B(n_350), .Y(n_477) );
INVx2_ASAP7_75t_SL g482 ( .A(n_315), .Y(n_482) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g364 ( .A(n_318), .Y(n_364) );
AND2x4_ASAP7_75t_L g340 ( .A(n_319), .B(n_329), .Y(n_340) );
INVx2_ASAP7_75t_L g404 ( .A(n_319), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_319), .B(n_345), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_319), .B(n_375), .Y(n_491) );
AOI221x1_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_327), .B1(n_332), .B2(n_340), .C(n_341), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx2_ASAP7_75t_L g460 ( .A(n_323), .Y(n_460) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_323), .A2(n_468), .B(n_470), .Y(n_467) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g349 ( .A(n_324), .B(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
AND2x4_ASAP7_75t_L g434 ( .A(n_324), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g394 ( .A(n_326), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI32xp33_ASAP7_75t_L g439 ( .A1(n_328), .A2(n_437), .A3(n_440), .B1(n_442), .B2(n_443), .Y(n_439) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_329), .B(n_346), .Y(n_462) );
AND2x2_ASAP7_75t_L g478 ( .A(n_329), .B(n_358), .Y(n_478) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_333), .B(n_335), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_334), .B(n_476), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g410 ( .A1(n_335), .A2(n_411), .B(n_414), .C(n_416), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_348), .B(n_351), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g376 ( .A1(n_342), .A2(n_377), .B(n_379), .Y(n_376) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_345), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_349), .A2(n_422), .B1(n_426), .B2(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g488 ( .A(n_349), .B(n_476), .Y(n_488) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_376), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_359), .B1(n_360), .B2(n_362), .C(n_366), .Y(n_354) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_355), .A2(n_465), .B(n_466), .Y(n_464) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g447 ( .A(n_361), .B(n_413), .Y(n_447) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AOI31xp33_ASAP7_75t_L g384 ( .A1(n_364), .A2(n_385), .A3(n_390), .B(n_392), .Y(n_384) );
AND2x2_ASAP7_75t_L g484 ( .A(n_364), .B(n_391), .Y(n_484) );
AND2x2_ASAP7_75t_L g373 ( .A(n_365), .B(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_365), .Y(n_437) );
INVx1_ASAP7_75t_L g471 ( .A(n_365), .Y(n_471) );
OAI21xp33_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_370), .B(n_373), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g397 ( .A(n_369), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_369), .B(n_496), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_370), .A2(n_453), .B(n_455), .Y(n_452) );
NOR2x1p5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_372), .A2(n_387), .B(n_394), .C(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g406 ( .A(n_375), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g426 ( .A(n_375), .B(n_382), .Y(n_426) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
INVx1_ASAP7_75t_L g444 ( .A(n_383), .Y(n_444) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_389), .A2(n_406), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g465 ( .A(n_389), .Y(n_465) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_451), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_419), .C(n_429), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_405), .B1(n_406), .B2(n_409), .C(n_410), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_407), .A2(n_474), .B1(n_477), .B2(n_478), .Y(n_473) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g470 ( .A(n_418), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g469 ( .A(n_424), .Y(n_469) );
INVx2_ASAP7_75t_L g449 ( .A(n_426), .Y(n_449) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI211xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B(n_439), .C(n_445), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_438), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g440 ( .A(n_435), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B1(n_449), .B2(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND4xp75_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .C(n_472), .D(n_485), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_461), .B2(n_462), .Y(n_455) );
NAND2x1_ASAP7_75t_SL g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_479), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B(n_484), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_488), .B1(n_489), .B2(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVxp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g506 ( .A(n_497), .Y(n_506) );
XOR2xp5_ASAP7_75t_L g906 ( .A(n_497), .B(n_907), .Y(n_906) );
XNOR2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_500), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_502), .A2(n_905), .B1(n_912), .B2(n_919), .Y(n_904) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g520 ( .A(n_511), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_511), .B(n_901), .Y(n_900) );
INVx3_ASAP7_75t_L g915 ( .A(n_511), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_511), .B(n_918), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
NOR2xp67_ASAP7_75t_R g513 ( .A(n_514), .B(n_518), .Y(n_513) );
AOI31xp33_ASAP7_75t_L g889 ( .A1(n_514), .A2(n_519), .A3(n_525), .B(n_890), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
INVx5_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x6_ASAP7_75t_SL g519 ( .A(n_520), .B(n_521), .Y(n_519) );
BUFx3_ASAP7_75t_L g891 ( .A(n_520), .Y(n_891) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
XNOR2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
BUFx8_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_534), .Y(n_888) );
AND2x2_ASAP7_75t_L g902 ( .A(n_534), .B(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_819), .Y(n_537) );
NAND4xp25_ASAP7_75t_L g538 ( .A(n_539), .B(n_694), .C(n_734), .D(n_783), .Y(n_538) );
NOR2xp67_ASAP7_75t_L g539 ( .A(n_540), .B(n_645), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_570), .B1(n_619), .B2(n_628), .Y(n_540) );
INVx1_ASAP7_75t_L g815 ( .A(n_541), .Y(n_815) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_542), .B(n_664), .Y(n_731) );
AND2x2_ASAP7_75t_L g762 ( .A(n_542), .B(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_557), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_543), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g686 ( .A(n_543), .Y(n_686) );
AND2x2_ASAP7_75t_L g861 ( .A(n_543), .B(n_729), .Y(n_861) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g630 ( .A(n_544), .Y(n_630) );
AND2x2_ASAP7_75t_L g714 ( .A(n_544), .B(n_676), .Y(n_714) );
AND2x2_ASAP7_75t_L g758 ( .A(n_544), .B(n_665), .Y(n_758) );
OR2x2_ASAP7_75t_L g776 ( .A(n_544), .B(n_777), .Y(n_776) );
INVx4_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g680 ( .A(n_545), .B(n_665), .Y(n_680) );
BUFx2_ASAP7_75t_L g737 ( .A(n_545), .Y(n_737) );
OR2x2_ASAP7_75t_L g745 ( .A(n_545), .B(n_703), .Y(n_745) );
INVx1_ASAP7_75t_L g800 ( .A(n_545), .Y(n_800) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
OAI21x1_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_552), .B(n_556), .Y(n_547) );
AND2x2_ASAP7_75t_L g631 ( .A(n_557), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g739 ( .A(n_557), .B(n_716), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_557), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g777 ( .A(n_558), .Y(n_777) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_558), .Y(n_782) );
AND2x2_ASAP7_75t_L g799 ( .A(n_558), .B(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g689 ( .A(n_559), .B(n_633), .Y(n_689) );
INVx1_ASAP7_75t_L g703 ( .A(n_559), .Y(n_703) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_568), .Y(n_559) );
NAND2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_583), .Y(n_570) );
AND2x4_ASAP7_75t_L g864 ( .A(n_571), .B(n_792), .Y(n_864) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_572), .Y(n_627) );
BUFx3_ASAP7_75t_L g660 ( .A(n_572), .Y(n_660) );
INVx1_ASAP7_75t_L g724 ( .A(n_572), .Y(n_724) );
AND2x2_ASAP7_75t_L g727 ( .A(n_572), .B(n_586), .Y(n_727) );
AND2x2_ASAP7_75t_L g752 ( .A(n_572), .B(n_609), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_572), .Y(n_755) );
AND2x2_ASAP7_75t_L g787 ( .A(n_572), .B(n_654), .Y(n_787) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_596), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g696 ( .A(n_585), .B(n_682), .Y(n_696) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g722 ( .A(n_587), .B(n_709), .Y(n_722) );
AND2x2_ASAP7_75t_L g751 ( .A(n_587), .B(n_598), .Y(n_751) );
OR2x2_ASAP7_75t_L g847 ( .A(n_587), .B(n_598), .Y(n_847) );
AND2x2_ASAP7_75t_L g726 ( .A(n_596), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g875 ( .A(n_596), .Y(n_875) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_597), .Y(n_621) );
OR2x2_ASAP7_75t_L g809 ( .A(n_597), .B(n_623), .Y(n_809) );
INVx1_ASAP7_75t_L g831 ( .A(n_597), .Y(n_831) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_609), .Y(n_597) );
AND2x2_ASAP7_75t_L g649 ( .A(n_598), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g682 ( .A(n_598), .B(n_654), .Y(n_682) );
INVx1_ASAP7_75t_L g709 ( .A(n_598), .Y(n_709) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_598), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_598), .B(n_609), .Y(n_796) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_605), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g635 ( .A(n_606), .Y(n_635) );
AND2x2_ASAP7_75t_L g733 ( .A(n_609), .B(n_655), .Y(n_733) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR3x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .C(n_626), .Y(n_620) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_623), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g681 ( .A(n_623), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g732 ( .A(n_623), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g772 ( .A(n_623), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_623), .B(n_795), .Y(n_827) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp67_ASAP7_75t_L g768 ( .A(n_624), .B(n_708), .Y(n_768) );
AND2x2_ASAP7_75t_L g792 ( .A(n_624), .B(n_654), .Y(n_792) );
BUFx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g650 ( .A(n_625), .Y(n_650) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g803 ( .A(n_627), .B(n_682), .Y(n_803) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_630), .B(n_689), .Y(n_868) );
AND2x4_ASAP7_75t_L g860 ( .A(n_631), .B(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_631), .B(n_680), .Y(n_874) );
INVx2_ASAP7_75t_L g676 ( .A(n_632), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_632), .Y(n_679) );
INVx2_ASAP7_75t_L g764 ( .A(n_632), .Y(n_764) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g748 ( .A(n_633), .Y(n_748) );
AOI21x1_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_644), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_640), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_683), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_661), .B1(n_677), .B2(n_681), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_656), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g711 ( .A(n_649), .B(n_660), .Y(n_711) );
AND2x2_ASAP7_75t_L g871 ( .A(n_649), .B(n_752), .Y(n_871) );
BUFx2_ASAP7_75t_L g742 ( .A(n_650), .Y(n_742) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g741 ( .A(n_653), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_654), .Y(n_658) );
INVx1_ASAP7_75t_L g708 ( .A(n_654), .Y(n_708) );
INVx1_ASAP7_75t_L g833 ( .A(n_655), .Y(n_833) );
AOI31xp33_ASAP7_75t_L g851 ( .A1(n_656), .A2(n_852), .A3(n_853), .B(n_854), .Y(n_851) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_657), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_658), .B(n_751), .Y(n_850) );
INVx2_ASAP7_75t_L g878 ( .A(n_658), .Y(n_878) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_659), .Y(n_693) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g706 ( .A(n_660), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_660), .B(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g836 ( .A(n_660), .B(n_796), .Y(n_836) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_675), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g747 ( .A(n_665), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g716 ( .A(n_666), .Y(n_716) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_679), .Y(n_700) );
INVx1_ASAP7_75t_L g740 ( .A(n_679), .Y(n_740) );
INVx1_ASAP7_75t_L g720 ( .A(n_680), .Y(n_720) );
AND2x2_ASAP7_75t_L g781 ( .A(n_680), .B(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g837 ( .A(n_680), .B(n_764), .Y(n_837) );
OAI21xp5_ASAP7_75t_L g753 ( .A1(n_681), .A2(n_754), .B(n_756), .Y(n_753) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_693), .Y(n_683) );
NAND3x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .C(n_690), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g855 ( .A(n_686), .B(n_775), .Y(n_855) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2x1_ASAP7_75t_SL g808 ( .A(n_688), .B(n_720), .Y(n_808) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g728 ( .A(n_689), .B(n_729), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_690), .B(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_690), .B(n_799), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_690), .B(n_799), .Y(n_872) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g775 ( .A(n_692), .B(n_748), .Y(n_775) );
AND2x2_ASAP7_75t_L g695 ( .A(n_693), .B(n_696), .Y(n_695) );
AOI221x1_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_697), .B1(n_704), .B2(n_713), .C(n_717), .Y(n_694) );
AOI32xp33_ASAP7_75t_L g876 ( .A1(n_696), .A2(n_877), .A3(n_882), .B1(n_883), .B2(n_885), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_701), .B(n_855), .Y(n_854) );
BUFx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g715 ( .A(n_703), .B(n_716), .Y(n_715) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_703), .Y(n_719) );
OR2x2_ASAP7_75t_L g832 ( .A(n_703), .B(n_833), .Y(n_832) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_710), .C(n_712), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g754 ( .A(n_707), .B(n_755), .Y(n_754) );
AND2x4_ASAP7_75t_L g771 ( .A(n_707), .B(n_772), .Y(n_771) );
AND2x4_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_710), .A2(n_807), .B1(n_809), .B2(n_810), .Y(n_806) );
INVx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g884 ( .A(n_714), .Y(n_884) );
INVx2_ASAP7_75t_L g729 ( .A(n_716), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_721), .B(n_725), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g853 ( .A(n_722), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_723), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_730), .B2(n_732), .Y(n_725) );
AND2x4_ASAP7_75t_L g822 ( .A(n_728), .B(n_737), .Y(n_822) );
INVx1_ASAP7_75t_L g881 ( .A(n_729), .Y(n_881) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g760 ( .A(n_733), .B(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_733), .B(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_733), .B(n_761), .Y(n_852) );
AOI211x1_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_741), .B(n_743), .C(n_769), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OR3x2_ASAP7_75t_L g844 ( .A(n_737), .B(n_739), .C(n_740), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_738), .A2(n_760), .B1(n_762), .B2(n_765), .Y(n_759) );
NOR2x1p5_ASAP7_75t_SL g738 ( .A(n_739), .B(n_740), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_739), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_877) );
INVx2_ASAP7_75t_L g761 ( .A(n_742), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_749), .B(n_753), .C(n_759), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_751), .B(n_755), .Y(n_766) );
INVx1_ASAP7_75t_L g793 ( .A(n_751), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_751), .B(n_858), .Y(n_866) );
OAI32xp33_ASAP7_75t_L g841 ( .A1(n_752), .A2(n_797), .A3(n_842), .B1(n_844), .B2(n_845), .Y(n_841) );
INVx1_ASAP7_75t_L g858 ( .A(n_752), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_752), .B(n_772), .Y(n_862) );
NAND2xp5_ASAP7_75t_SL g824 ( .A(n_755), .B(n_789), .Y(n_824) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g802 ( .A(n_761), .B(n_787), .Y(n_802) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g811 ( .A(n_764), .B(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g779 ( .A(n_767), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_773), .B1(n_778), .B2(n_780), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g817 ( .A(n_774), .Y(n_817) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AND2x2_ASAP7_75t_L g798 ( .A(n_775), .B(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_775), .B(n_782), .Y(n_886) );
INVx1_ASAP7_75t_SL g812 ( .A(n_776), .Y(n_812) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NOR3xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_806), .C(n_813), .Y(n_783) );
OAI21xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_797), .B(n_801), .Y(n_784) );
NOR2xp33_ASAP7_75t_SL g785 ( .A(n_786), .B(n_790), .Y(n_785) );
INVxp67_ASAP7_75t_L g818 ( .A(n_786), .Y(n_818) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g843 ( .A(n_788), .Y(n_843) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .C(n_794), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g805 ( .A(n_799), .Y(n_805) );
OAI21xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .B(n_804), .Y(n_801) );
INVx1_ASAP7_75t_L g814 ( .A(n_802), .Y(n_814) );
OAI221xp5_ASAP7_75t_L g857 ( .A1(n_807), .A2(n_858), .B1(n_859), .B2(n_862), .C(n_863), .Y(n_857) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI32xp33_ASAP7_75t_L g813 ( .A1(n_810), .A2(n_814), .A3(n_815), .B1(n_816), .B2(n_818), .Y(n_813) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI221xp5_ASAP7_75t_L g825 ( .A1(n_816), .A2(n_826), .B1(n_827), .B2(n_828), .C(n_834), .Y(n_825) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_838), .C(n_856), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B(n_825), .Y(n_820) );
AOI211x1_ASAP7_75t_L g838 ( .A1(n_821), .A2(n_839), .B(n_841), .C(n_848), .Y(n_838) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVxp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2x1_ASAP7_75t_SL g829 ( .A(n_830), .B(n_832), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g840 ( .A(n_831), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_837), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
AO21x1_ASAP7_75t_L g848 ( .A1(n_837), .A2(n_849), .B(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g882 ( .A(n_853), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_869), .Y(n_856) );
INVx3_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OAI21xp33_ASAP7_75t_SL g863 ( .A1(n_864), .A2(n_865), .B(n_867), .Y(n_863) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_876), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B(n_873), .Y(n_870) );
NOR2xp67_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g879 ( .A(n_878), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
BUFx12f_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B1(n_897), .B2(n_898), .Y(n_890) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
AOI21xp33_ASAP7_75t_SL g905 ( .A1(n_893), .A2(n_906), .B(n_909), .Y(n_905) );
NOR2x1_ASAP7_75t_R g893 ( .A(n_894), .B(n_895), .Y(n_893) );
BUFx12f_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
BUFx10_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
OR2x6_ASAP7_75t_L g912 ( .A(n_913), .B(n_918), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
OR2x4_ASAP7_75t_L g921 ( .A(n_916), .B(n_922), .Y(n_921) );
BUFx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx4_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
BUFx3_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
endmodule