module fake_aes_6244_n_346 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_346);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_346;
wire n_117;
wire n_185;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_252;
wire n_152;
wire n_113;
wire n_206;
wire n_288;
wire n_296;
wire n_157;
wire n_202;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_163;
wire n_105;
wire n_227;
wire n_231;
wire n_298;
wire n_144;
wire n_183;
wire n_199;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_236;
wire n_340;
wire n_150;
wire n_301;
wire n_222;
wire n_234;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_247;
wire n_304;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_235;
wire n_243;
wire n_331;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_88;
wire n_107;
wire n_254;
wire n_262;
wire n_239;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_342;
wire n_217;
wire n_139;
wire n_193;
wire n_273;
wire n_120;
wire n_245;
wire n_90;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_179;
wire n_315;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_344;
wire n_136;
wire n_283;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_168;
wire n_134;
wire n_233;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_225;
wire n_220;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_103;
wire n_180;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_188;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_138;
wire n_323;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_226;
wire n_159;
wire n_337;
wire n_176;
wire n_123;
wire n_223;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_164;
wire n_175;
wire n_145;
wire n_290;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_151;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g88 ( .A(n_52), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_23), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_8), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_50), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_56), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_46), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_72), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_71), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_73), .Y(n_97) );
INVx2_ASAP7_75t_SL g98 ( .A(n_77), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_45), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_76), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_75), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_58), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_59), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_80), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_81), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_78), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_68), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_30), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_44), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_16), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_82), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_36), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_55), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_57), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_27), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_53), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_32), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_28), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_35), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_63), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_54), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_65), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_29), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_26), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_70), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_69), .Y(n_132) );
INVxp33_ASAP7_75t_SL g133 ( .A(n_15), .Y(n_133) );
INVx4_ASAP7_75t_R g134 ( .A(n_85), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_37), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_20), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_34), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_41), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_40), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_60), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_21), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_7), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_22), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_12), .Y(n_144) );
CKINVDCx14_ASAP7_75t_R g145 ( .A(n_67), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_87), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_14), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_79), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_43), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_61), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_30), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_27), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_86), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_133), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_102), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_108), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_98), .B(n_0), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_112), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_90), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_113), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_130), .B(n_2), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_90), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_114), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_113), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_102), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_153), .B(n_3), .Y(n_168) );
BUFx8_ASAP7_75t_L g169 ( .A(n_102), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_119), .B(n_3), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_119), .B(n_4), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_93), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_91), .B(n_4), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_95), .B(n_5), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_102), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_117), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_169), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_170), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_169), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_160), .B(n_95), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_166), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_166), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_164), .B(n_145), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_164), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_170), .B(n_93), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
NAND2xp33_ASAP7_75t_L g195 ( .A(n_161), .B(n_117), .Y(n_195) );
INVxp67_ASAP7_75t_SL g196 ( .A(n_171), .Y(n_196) );
INVxp33_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_163), .B(n_96), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_172), .B(n_122), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_172), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_169), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_167), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_162), .B(n_115), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_172), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_173), .B(n_96), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_167), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_197), .B(n_175), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_192), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_197), .B(n_168), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_208), .B(n_157), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_182), .B(n_174), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_196), .B(n_89), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_185), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_186), .B(n_154), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_208), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_185), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_179), .B(n_146), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_198), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_180), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_198), .Y(n_225) );
INVx4_ASAP7_75t_SL g226 ( .A(n_181), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_188), .B(n_92), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_188), .B(n_126), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_188), .B(n_92), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_200), .Y(n_232) );
AND2x6_ASAP7_75t_L g233 ( .A(n_206), .B(n_88), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_204), .B(n_105), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_209), .A2(n_158), .B1(n_159), .B2(n_156), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_203), .A2(n_158), .B1(n_159), .B2(n_156), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_220), .B(n_203), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_213), .B(n_203), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_228), .A2(n_193), .B(n_187), .Y(n_239) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_230), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g241 ( .A1(n_215), .A2(n_203), .B(n_201), .C(n_210), .Y(n_241) );
OAI21xp33_ASAP7_75t_L g242 ( .A1(n_216), .A2(n_201), .B(n_187), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_214), .B(n_184), .Y(n_243) );
NAND2xp33_ASAP7_75t_L g244 ( .A(n_233), .B(n_184), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_216), .B(n_136), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_219), .A2(n_142), .B1(n_143), .B2(n_141), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_217), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_231), .A2(n_195), .B(n_211), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_235), .A2(n_151), .B1(n_152), .B2(n_147), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_229), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_232), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_212), .B(n_148), .Y(n_252) );
OAI22xp33_ASAP7_75t_L g253 ( .A1(n_234), .A2(n_150), .B1(n_127), .B2(n_177), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_234), .A2(n_127), .B1(n_94), .B2(n_97), .Y(n_254) );
CKINVDCx6p67_ASAP7_75t_R g255 ( .A(n_233), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_236), .B(n_118), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_224), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_222), .B(n_121), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_226), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_223), .A2(n_99), .B(n_101), .C(n_100), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_225), .B(n_103), .Y(n_261) );
AOI22x1_ASAP7_75t_L g262 ( .A1(n_218), .A2(n_178), .B1(n_176), .B2(n_124), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_235), .B(n_104), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_221), .A2(n_107), .B(n_106), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_227), .A2(n_110), .B(n_109), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_250), .B(n_111), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_238), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_251), .B(n_116), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_248), .A2(n_140), .B(n_120), .Y(n_269) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_239), .A2(n_128), .B(n_125), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g271 ( .A1(n_246), .A2(n_149), .B1(n_131), .B2(n_132), .C(n_137), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_241), .A2(n_139), .B(n_138), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_262), .A2(n_190), .B(n_189), .Y(n_273) );
OAI21x1_ASAP7_75t_SL g274 ( .A1(n_237), .A2(n_134), .B(n_176), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_237), .A2(n_207), .B(n_191), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_259), .B(n_117), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_247), .B(n_6), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_261), .A2(n_191), .B(n_189), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_264), .A2(n_202), .B(n_178), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_243), .A2(n_176), .B(n_123), .Y(n_280) );
AND2x6_ASAP7_75t_L g281 ( .A(n_259), .B(n_135), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_240), .A2(n_205), .B1(n_194), .B2(n_183), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_255), .A2(n_205), .B1(n_194), .B2(n_183), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_265), .A2(n_33), .B(n_31), .Y(n_284) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_244), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_263), .A2(n_205), .B1(n_194), .B2(n_183), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_245), .A2(n_205), .B1(n_194), .B2(n_183), .C(n_10), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_242), .A2(n_205), .B(n_194), .C(n_183), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_242), .A2(n_205), .B(n_194), .C(n_183), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_253), .A2(n_205), .B(n_194), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_263), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_260), .A2(n_252), .B(n_249), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_254), .A2(n_42), .B(n_39), .Y(n_293) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_257), .A2(n_17), .B(n_19), .Y(n_294) );
AOI21xp33_ASAP7_75t_L g295 ( .A1(n_292), .A2(n_258), .B(n_256), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_271), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_296) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_289), .A2(n_47), .B(n_48), .Y(n_297) );
AOI21xp33_ASAP7_75t_L g298 ( .A1(n_270), .A2(n_49), .B(n_51), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_285), .A2(n_64), .B(n_66), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_291), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_291), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_287), .A2(n_267), .B1(n_266), .B2(n_268), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_290), .A2(n_269), .B(n_286), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_294), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_276), .A2(n_286), .B1(n_280), .B2(n_283), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_290), .A2(n_278), .B(n_275), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_282), .A2(n_272), .B1(n_274), .B2(n_281), .Y(n_308) );
AOI21xp33_ASAP7_75t_L g309 ( .A1(n_293), .A2(n_284), .B(n_279), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_273), .A2(n_289), .B(n_288), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_304), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_301), .B(n_302), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_296), .B(n_295), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_295), .B(n_300), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_297), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_310), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_310), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_299), .B(n_308), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_306), .B(n_298), .Y(n_320) );
AO31x2_ASAP7_75t_L g321 ( .A1(n_309), .A2(n_307), .A3(n_305), .B(n_303), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_312), .B(n_314), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_312), .B(n_314), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_319), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_311), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_313), .B(n_320), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_316), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_321), .B(n_318), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_326), .B(n_317), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_322), .B(n_315), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_323), .B(n_315), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_329), .B(n_328), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_330), .B(n_324), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_332), .B(n_331), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_333), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_334), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_336), .B(n_335), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_337), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_338), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_339), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_340), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_341), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_342), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_343), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_344), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_345), .A2(n_325), .B(n_327), .Y(n_346) );
endmodule