module fake_jpeg_13715_n_475 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_475);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_475;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_73),
.Y(n_118)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g173 ( 
.A(n_65),
.Y(n_173)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_72),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_76),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_80),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_90),
.Y(n_193)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_50),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_92),
.B(n_114),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

NAND2x1_ASAP7_75t_SL g104 ( 
.A(n_20),
.B(n_1),
.Y(n_104)
);

OR2x2_ASAP7_75t_SL g142 ( 
.A(n_104),
.B(n_44),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_111),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_25),
.B(n_17),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_48),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_55),
.B1(n_52),
.B2(n_43),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_120),
.A2(n_157),
.B1(n_169),
.B2(n_189),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_31),
.B(n_29),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_131),
.B(n_158),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_57),
.A2(n_52),
.B1(n_55),
.B2(n_29),
.Y(n_134)
);

OAI22x1_ASAP7_75t_L g213 ( 
.A1(n_134),
.A2(n_162),
.B1(n_178),
.B2(n_9),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_56),
.A2(n_52),
.B1(n_47),
.B2(n_31),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_137),
.A2(n_153),
.B1(n_86),
.B2(n_7),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_77),
.B(n_26),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_138),
.B(n_139),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_26),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_142),
.A2(n_3),
.B(n_4),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_47),
.C(n_49),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_9),
.C(n_10),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_65),
.B(n_25),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_161),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_83),
.A2(n_54),
.B1(n_53),
.B2(n_51),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_68),
.B(n_54),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_179),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_70),
.A2(n_49),
.B1(n_53),
.B2(n_51),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_87),
.A2(n_44),
.B1(n_46),
.B2(n_38),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_59),
.B(n_46),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_88),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_42),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_164),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_95),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_99),
.A2(n_35),
.B1(n_32),
.B2(n_48),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_102),
.B(n_32),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_1),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_180),
.B(n_125),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_105),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_191),
.A2(n_115),
.B1(n_113),
.B2(n_109),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_195),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_107),
.B1(n_62),
.B2(n_48),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_196),
.Y(n_261)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_197),
.B(n_203),
.Y(n_280)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_199),
.Y(n_292)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_200),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_201),
.B(n_212),
.Y(n_264)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_122),
.A2(n_30),
.B1(n_5),
.B2(n_6),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_204),
.A2(n_206),
.B1(n_210),
.B2(n_213),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_30),
.B1(n_5),
.B2(n_7),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_205),
.A2(n_216),
.B(n_236),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_30),
.B1(n_7),
.B2(n_8),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_209),
.A2(n_229),
.B1(n_195),
.B2(n_219),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_165),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_140),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_214),
.B(n_222),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_118),
.B(n_11),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_218),
.B(n_239),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_137),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_219),
.A2(n_245),
.B1(n_200),
.B2(n_220),
.Y(n_275)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_159),
.A2(n_194),
.B1(n_181),
.B2(n_130),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_133),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_149),
.B1(n_132),
.B2(n_152),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_150),
.B(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_120),
.A2(n_14),
.B1(n_15),
.B2(n_134),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_227),
.A2(n_241),
.B1(n_244),
.B2(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_185),
.A2(n_146),
.B1(n_188),
.B2(n_183),
.Y(n_229)
);

AO22x2_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_184),
.B1(n_167),
.B2(n_175),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_235),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_126),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_231),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_173),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_234),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_187),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_233),
.Y(n_266)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_136),
.A2(n_176),
.B1(n_192),
.B2(n_155),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_237),
.B(n_238),
.Y(n_298)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_171),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_246),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_178),
.A2(n_162),
.B1(n_125),
.B2(n_129),
.Y(n_241)
);

INVx4_ASAP7_75t_SL g242 ( 
.A(n_173),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_242),
.B(n_243),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_177),
.B(n_174),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_193),
.A2(n_167),
.B1(n_166),
.B2(n_174),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_193),
.A2(n_129),
.B1(n_124),
.B2(n_141),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_148),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_248),
.Y(n_279)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_251),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_124),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_141),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_253),
.Y(n_286)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_257),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_190),
.A2(n_120),
.B1(n_131),
.B2(n_149),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_143),
.Y(n_257)
);

AOI32xp33_ASAP7_75t_L g258 ( 
.A1(n_208),
.A2(n_235),
.A3(n_202),
.B1(n_211),
.B2(n_255),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_258),
.B(n_264),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_302),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_209),
.A2(n_150),
.B1(n_225),
.B2(n_256),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_265),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_212),
.B(n_255),
.CI(n_201),
.CON(n_268),
.SN(n_268)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_264),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_227),
.C(n_217),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_297),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_271),
.A2(n_299),
.B1(n_266),
.B2(n_285),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_213),
.A2(n_241),
.B1(n_196),
.B2(n_245),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_196),
.A2(n_244),
.B1(n_230),
.B2(n_248),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_196),
.A2(n_244),
.B1(n_230),
.B2(n_254),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_291),
.A2(n_295),
.B1(n_302),
.B2(n_274),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_198),
.B(n_224),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_285),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_244),
.A2(n_230),
.B1(n_234),
.B2(n_251),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_247),
.C(n_240),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_233),
.A2(n_242),
.B1(n_207),
.B2(n_231),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_231),
.A2(n_256),
.B1(n_227),
.B2(n_249),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_303),
.B1(n_284),
.B2(n_261),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_253),
.A2(n_235),
.B1(n_209),
.B2(n_225),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_249),
.B1(n_227),
.B2(n_241),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_307),
.Y(n_341)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_280),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_326),
.B1(n_333),
.B2(n_288),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_310),
.A2(n_311),
.B(n_339),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_267),
.B(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_313),
.B(n_331),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_318),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_258),
.B(n_264),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_329),
.C(n_296),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_262),
.B(n_259),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_316),
.A2(n_310),
.B(n_330),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_293),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_319),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_276),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_327),
.Y(n_354)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_336),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_323),
.B(n_337),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_324),
.A2(n_335),
.B1(n_338),
.B2(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_303),
.A2(n_284),
.B1(n_261),
.B2(n_287),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_286),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_328),
.B(n_330),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_268),
.B(n_265),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_278),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_292),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_287),
.A2(n_269),
.B1(n_273),
.B2(n_294),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_295),
.B1(n_269),
.B2(n_275),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_298),
.B(n_283),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_268),
.B1(n_282),
.B2(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_340),
.A2(n_282),
.B1(n_292),
.B2(n_288),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_357),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_349),
.B(n_363),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_309),
.A2(n_297),
.B1(n_272),
.B2(n_300),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_352),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_316),
.A2(n_292),
.B(n_283),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_333),
.B1(n_310),
.B2(n_319),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_322),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_366),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_356),
.A2(n_359),
.B1(n_365),
.B2(n_344),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g357 ( 
.A1(n_319),
.A2(n_281),
.B(n_260),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_358),
.A2(n_314),
.B(n_312),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_317),
.A2(n_260),
.B1(n_296),
.B2(n_335),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_323),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_312),
.A2(n_339),
.B(n_329),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_317),
.A2(n_324),
.B1(n_338),
.B2(n_332),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_325),
.B1(n_321),
.B2(n_318),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_346),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_373),
.Y(n_392)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_370),
.A2(n_387),
.B(n_351),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_360),
.C(n_367),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_346),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_364),
.Y(n_374)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_305),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_380),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_359),
.A2(n_365),
.B1(n_356),
.B2(n_353),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_378),
.A2(n_384),
.B1(n_385),
.B2(n_343),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_362),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_358),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_381),
.B(n_382),
.Y(n_398)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_383),
.B(n_386),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_353),
.A2(n_328),
.B1(n_307),
.B2(n_315),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_363),
.A2(n_308),
.B(n_336),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_306),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_388),
.Y(n_401)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_389),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_334),
.B(n_352),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_391),
.A2(n_347),
.B(n_349),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_393),
.A2(n_403),
.B1(n_348),
.B2(n_385),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_360),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_397),
.C(n_400),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_367),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_402),
.A2(n_371),
.B1(n_379),
.B2(n_399),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_344),
.B1(n_351),
.B2(n_357),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_367),
.C(n_344),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_387),
.C(n_388),
.Y(n_415)
);

NOR2x1_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_361),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_406),
.B(n_408),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_390),
.A2(n_341),
.B(n_345),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_377),
.Y(n_425)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_379),
.A2(n_341),
.B(n_366),
.C(n_354),
.Y(n_411)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_411),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_370),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_417),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_414),
.A2(n_423),
.B1(n_408),
.B2(n_398),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_419),
.Y(n_435)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_416),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_384),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_387),
.C(n_391),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_422),
.C(n_397),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_390),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_393),
.A2(n_385),
.B1(n_378),
.B2(n_380),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_421),
.A2(n_424),
.B1(n_426),
.B2(n_408),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_379),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_402),
.A2(n_368),
.B1(n_373),
.B2(n_376),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_411),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_403),
.B1(n_399),
.B2(n_396),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_428),
.A2(n_436),
.B1(n_438),
.B2(n_414),
.Y(n_449)
);

OAI21xp33_ASAP7_75t_L g429 ( 
.A1(n_427),
.A2(n_392),
.B(n_395),
.Y(n_429)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_429),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_345),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_430),
.B(n_354),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_433),
.A2(n_418),
.B1(n_419),
.B2(n_401),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_401),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_439),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_424),
.B1(n_420),
.B2(n_410),
.Y(n_436)
);

XNOR2x1_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_413),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_420),
.A2(n_410),
.B1(n_396),
.B2(n_392),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_446),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_445),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_437),
.B(n_383),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_444),
.B(n_415),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_435),
.B(n_412),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_417),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_438),
.A2(n_427),
.B(n_411),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_447),
.A2(n_434),
.B(n_436),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_449),
.C(n_431),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_413),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_452),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_454),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_441),
.B(n_389),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_456),
.B(n_457),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_446),
.B(n_409),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_442),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_428),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_448),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_462),
.B(n_463),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_451),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_459),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_464),
.B(n_465),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_461),
.B(n_407),
.Y(n_467)
);

NAND4xp25_ASAP7_75t_SL g469 ( 
.A(n_467),
.B(n_376),
.C(n_406),
.D(n_407),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_432),
.C(n_447),
.Y(n_470)
);

NOR3xp33_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_468),
.C(n_466),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_471),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_472),
.A2(n_458),
.B(n_416),
.Y(n_473)
);

AOI321xp33_ASAP7_75t_SL g474 ( 
.A1(n_473),
.A2(n_458),
.A3(n_460),
.B1(n_433),
.B2(n_445),
.C(n_409),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_474),
.A2(n_398),
.B(n_431),
.Y(n_475)
);


endmodule