module fake_ariane_110_n_1878 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1878);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1878;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1608;
wire n_1304;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1806;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_3),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_40),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_2),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_42),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_63),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_67),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_16),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_9),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_100),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_43),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_28),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_24),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_81),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_8),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_43),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_142),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_104),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_131),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_44),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_135),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_99),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_72),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_77),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_157),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_49),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_82),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_74),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_103),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_79),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_50),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_95),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_123),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_28),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_31),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_36),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_22),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_97),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_86),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_35),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_154),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_96),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_92),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_122),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_1),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_32),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_137),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_47),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_130),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_75),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_119),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_69),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_114),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_83),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_23),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_61),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_153),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_132),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_71),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_7),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_84),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_57),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_115),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_105),
.Y(n_265)
);

INVx4_ASAP7_75t_R g266 ( 
.A(n_13),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_116),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_5),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_88),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_25),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_10),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_125),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_70),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_20),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_59),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_37),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_41),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_10),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_102),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_136),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_62),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_162),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_15),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_63),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_61),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_144),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_29),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_12),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_9),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_107),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_89),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_163),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_168),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_118),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_7),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_56),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_27),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_27),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_160),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_167),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_78),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_57),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_76),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_165),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_110),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_38),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_117),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_152),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_51),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_36),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_49),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_101),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_133),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_26),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_22),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_150),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_170),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_0),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_55),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_94),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_141),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_121),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_145),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_139),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_50),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_171),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_4),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_172),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_149),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_35),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_0),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_120),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_169),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_66),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_65),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_5),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_134),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_12),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_140),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_21),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_158),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_98),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_87),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_109),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_85),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_33),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_93),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_146),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_108),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_23),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_38),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_40),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_45),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_106),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_25),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_111),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_14),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_31),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_44),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_205),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_207),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_245),
.B(n_6),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_296),
.B(n_6),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_358),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_296),
.B(n_8),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_251),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_205),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_273),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_358),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_251),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_358),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_358),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_208),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_264),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_265),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_210),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_210),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_212),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_309),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_185),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_176),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_178),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_212),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_325),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_214),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_214),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_218),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_353),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_218),
.B(n_11),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_220),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_254),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_312),
.B(n_11),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_179),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_220),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_224),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_245),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_224),
.Y(n_405)
);

BUFx6f_ASAP7_75t_SL g406 ( 
.A(n_208),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_237),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_182),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_237),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_186),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_292),
.B(n_13),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_239),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_239),
.B(n_14),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_247),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_247),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_189),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_177),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_176),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_192),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_204),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_253),
.B(n_15),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_358),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_193),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_253),
.Y(n_424)
);

BUFx2_ASAP7_75t_SL g425 ( 
.A(n_254),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_290),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_259),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_259),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_190),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_248),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_194),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_292),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_303),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_197),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_352),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_201),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_290),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_297),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_217),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_297),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_226),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_298),
.B(n_17),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_229),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_232),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_L g445 ( 
.A(n_303),
.B(n_18),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_363),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_238),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_208),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_256),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_254),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_298),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_261),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_246),
.B(n_18),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_328),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_263),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_268),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_328),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_190),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_275),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_254),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_354),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_331),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_278),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_R g464 ( 
.A(n_187),
.B(n_73),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_331),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_366),
.B(n_246),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_387),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_399),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_378),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_R g473 ( 
.A(n_380),
.B(n_188),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_371),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_422),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_183),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_367),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_377),
.B(n_359),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_366),
.B(n_181),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_417),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_368),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g489 ( 
.A(n_399),
.B(n_181),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_450),
.A2(n_257),
.B1(n_271),
.B2(n_316),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_373),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_374),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_373),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_374),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_383),
.B(n_384),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_382),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_450),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_384),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_373),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_420),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_385),
.B(n_334),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_391),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_430),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_427),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_427),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_460),
.A2(n_365),
.B1(n_364),
.B2(n_314),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_385),
.B(n_359),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_370),
.A2(n_215),
.B1(n_233),
.B2(n_234),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

AND2x2_ASAP7_75t_SL g515 ( 
.A(n_460),
.B(n_196),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_390),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_390),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_392),
.B(n_393),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_393),
.B(n_394),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_395),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_397),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_381),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_394),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_398),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_435),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_386),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_398),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_402),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_434),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_402),
.B(n_354),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_403),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_403),
.B(n_334),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_436),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_405),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_439),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_446),
.B(n_281),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_405),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_407),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_375),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_407),
.Y(n_542)
);

CKINVDCx8_ASAP7_75t_R g543 ( 
.A(n_441),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_443),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_444),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_489),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_470),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_467),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_481),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_531),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_489),
.A2(n_515),
.B1(n_513),
.B2(n_532),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_467),
.Y(n_552)
);

INVxp33_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_458),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_545),
.B(n_372),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_377),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_482),
.B(n_466),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_489),
.A2(n_400),
.B1(n_413),
.B2(n_396),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_495),
.B(n_338),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_466),
.B(n_428),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_486),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_521),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_406),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_492),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_479),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_406),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_492),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_535),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_521),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_515),
.A2(n_421),
.B1(n_432),
.B2(n_404),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_471),
.B(n_428),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_495),
.B(n_338),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_469),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_494),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_479),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_481),
.B(n_447),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_498),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_529),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_516),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_516),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_498),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_473),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_472),
.B(n_409),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_516),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_R g589 ( 
.A(n_537),
.B(n_544),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_483),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_495),
.B(n_518),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_406),
.Y(n_593)
);

INVx4_ASAP7_75t_SL g594 ( 
.A(n_485),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_510),
.B(n_452),
.C(n_449),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_488),
.B(n_455),
.Y(n_596)
);

CKINVDCx6p67_ASAP7_75t_R g597 ( 
.A(n_470),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_508),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_518),
.B(n_388),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_516),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_488),
.B(n_512),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_515),
.B(n_456),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_499),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_475),
.B(n_412),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_518),
.B(n_418),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_516),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_410),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_529),
.B(n_412),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_517),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_484),
.B(n_429),
.Y(n_610)
);

AND2x2_ASAP7_75t_SL g611 ( 
.A(n_497),
.B(n_442),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_516),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_512),
.B(n_459),
.Y(n_613)
);

BUFx4f_ASAP7_75t_L g614 ( 
.A(n_485),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_517),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_504),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_529),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_529),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_525),
.B(n_414),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_510),
.B(n_525),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_480),
.B(n_463),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_536),
.B(n_414),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_477),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_536),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_539),
.B(n_415),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_487),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_496),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_539),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_506),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_513),
.B(n_369),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_522),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_503),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_480),
.B(n_389),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_540),
.B(n_341),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_484),
.A2(n_404),
.B1(n_432),
.B2(n_433),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_508),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_504),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_477),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_540),
.B(n_341),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_542),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_519),
.B(n_415),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_519),
.B(n_424),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_476),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_508),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_519),
.B(n_424),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_543),
.B(n_345),
.Y(n_649)
);

AND3x1_ASAP7_75t_L g650 ( 
.A(n_490),
.B(n_199),
.C(n_191),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_508),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_526),
.B(n_426),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_526),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_526),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_497),
.B(n_543),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_484),
.A2(n_433),
.B1(n_445),
.B2(n_411),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_543),
.B(n_431),
.C(n_419),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_476),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_490),
.A2(n_453),
.B1(n_320),
.B2(n_288),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_523),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_476),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_502),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_502),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_502),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_468),
.B(n_448),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_530),
.B(n_347),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_530),
.B(n_347),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_524),
.B(n_426),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_533),
.B(n_437),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_533),
.B(n_195),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_484),
.B(n_437),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_476),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_478),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_476),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_478),
.Y(n_677)
);

AND3x2_ASAP7_75t_L g678 ( 
.A(n_468),
.B(n_199),
.C(n_191),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_468),
.B(n_440),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_511),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_511),
.B(n_196),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_509),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_507),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_528),
.B(n_440),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_527),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_505),
.B(n_451),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_541),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_538),
.B(n_451),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_485),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_511),
.B(n_454),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_485),
.B(n_195),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_505),
.B(n_213),
.Y(n_692)
);

AND2x6_ASAP7_75t_L g693 ( 
.A(n_534),
.B(n_228),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_534),
.B(n_454),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_562),
.A2(n_307),
.B(n_336),
.C(n_270),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_602),
.B(n_461),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_602),
.B(n_509),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_569),
.B(n_457),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_686),
.B(n_457),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_686),
.B(n_462),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_549),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_SL g702 ( 
.A1(n_546),
.A2(n_284),
.B1(n_361),
.B2(n_180),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_621),
.B(n_538),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_546),
.B(n_509),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_575),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_557),
.B(n_462),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_554),
.B(n_465),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_649),
.B(n_500),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_592),
.B(n_485),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_554),
.B(n_465),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_554),
.B(n_500),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_551),
.A2(n_324),
.B(n_280),
.C(n_276),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_649),
.B(n_500),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_592),
.B(n_500),
.Y(n_714)
);

NAND2x1_ASAP7_75t_L g715 ( 
.A(n_592),
.B(n_501),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_579),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_618),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_617),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_559),
.A2(n_485),
.B1(n_215),
.B2(n_233),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_607),
.B(n_501),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_549),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_592),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_592),
.B(n_501),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_596),
.B(n_284),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_563),
.B(n_501),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_565),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_563),
.B(n_485),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_613),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_635),
.B(n_284),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_566),
.B(n_485),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_673),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_566),
.B(n_491),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_617),
.B(n_213),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_694),
.B(n_491),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_556),
.B(n_491),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_680),
.A2(n_302),
.B(n_234),
.C(n_241),
.Y(n_736)
);

BUFx6f_ASAP7_75t_SL g737 ( 
.A(n_568),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_670),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_623),
.B(n_581),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_601),
.B(n_241),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_617),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_623),
.B(n_493),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_684),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_586),
.B(n_493),
.Y(n_744)
);

NOR2x1_ASAP7_75t_L g745 ( 
.A(n_595),
.B(n_240),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_618),
.B(n_322),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_514),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_601),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_616),
.B(n_361),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_593),
.B(n_514),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_620),
.B(n_618),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_564),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_611),
.B(n_322),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_601),
.B(n_249),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_559),
.A2(n_343),
.B1(n_362),
.B2(n_289),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_567),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_620),
.B(n_514),
.Y(n_757)
);

INVxp33_ASAP7_75t_L g758 ( 
.A(n_688),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_679),
.B(n_249),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_673),
.B(n_286),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_690),
.B(n_270),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_560),
.B(n_287),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_559),
.B(n_276),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_559),
.B(n_279),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_599),
.B(n_279),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_561),
.B(n_280),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_666),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_571),
.B(n_293),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_611),
.B(n_228),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_599),
.B(n_299),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_548),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_574),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_573),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_653),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_572),
.B(n_291),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_576),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_574),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_578),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_608),
.A2(n_626),
.B(n_619),
.C(n_580),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_583),
.B(n_231),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_568),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_568),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_599),
.B(n_300),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_644),
.A2(n_324),
.B(n_307),
.C(n_319),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_585),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_683),
.B(n_547),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_578),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_572),
.A2(n_336),
.B1(n_319),
.B2(n_302),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_572),
.A2(n_294),
.B1(n_269),
.B2(n_274),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_630),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_590),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_572),
.B(n_301),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_603),
.B(n_609),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_553),
.B(n_361),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_583),
.B(n_231),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_632),
.A2(n_346),
.B1(n_357),
.B2(n_356),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_552),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_615),
.B(n_311),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_627),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_625),
.B(n_315),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_605),
.B(n_323),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_629),
.Y(n_802)
);

BUFx5_ASAP7_75t_L g803 ( 
.A(n_681),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_583),
.B(n_243),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_642),
.Y(n_805)
);

AND2x6_ASAP7_75t_SL g806 ( 
.A(n_601),
.B(n_180),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_636),
.A2(n_180),
.B1(n_235),
.B2(n_330),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_643),
.B(n_332),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_SL g809 ( 
.A(n_550),
.B(n_335),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_645),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_648),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_605),
.B(n_337),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_652),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_605),
.B(n_342),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_628),
.B(n_243),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_644),
.A2(n_344),
.B(n_340),
.C(n_306),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_587),
.B(n_198),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_654),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_SL g819 ( 
.A(n_591),
.B(n_354),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_661),
.B(n_267),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_654),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_SL g822 ( 
.A(n_597),
.B(n_180),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_631),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_654),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_604),
.B(n_200),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_555),
.B(n_235),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_655),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_636),
.A2(n_632),
.B1(n_681),
.B2(n_693),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_671),
.B(n_202),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_552),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_671),
.B(n_203),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_669),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_610),
.B(n_206),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_610),
.B(n_209),
.Y(n_834)
);

BUFx12f_ASAP7_75t_SL g835 ( 
.A(n_632),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_584),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_553),
.B(n_235),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_610),
.B(n_211),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_582),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_634),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_675),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_600),
.B(n_285),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_677),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_636),
.B(n_464),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_692),
.B(n_216),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_653),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_600),
.B(n_285),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_681),
.B(n_219),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_631),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_582),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_584),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_699),
.A2(n_639),
.B1(n_632),
.B2(n_570),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_716),
.B(n_656),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_722),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_706),
.B(n_681),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_826),
.A2(n_589),
.B1(n_555),
.B2(n_681),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_700),
.B(n_657),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_739),
.A2(n_606),
.B(n_588),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_840),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_751),
.A2(n_641),
.B(n_658),
.C(n_614),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_707),
.B(n_710),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_788),
.A2(n_636),
.B1(n_660),
.B2(n_693),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_826),
.A2(n_589),
.B1(n_636),
.B2(n_597),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_728),
.A2(n_641),
.B(n_668),
.C(n_667),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_722),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_696),
.B(n_631),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_720),
.B(n_637),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_725),
.A2(n_606),
.B(n_588),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_720),
.B(n_693),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_732),
.A2(n_606),
.B(n_588),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_786),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_737),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_698),
.B(n_693),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_742),
.A2(n_612),
.B(n_584),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_835),
.B(n_633),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_810),
.B(n_693),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_722),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_722),
.B(n_633),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_751),
.A2(n_614),
.B(n_612),
.C(n_668),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_729),
.B(n_633),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_712),
.A2(n_667),
.B(n_672),
.C(n_612),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_774),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_717),
.A2(n_779),
.B(n_730),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_727),
.A2(n_651),
.B(n_647),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_711),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_811),
.B(n_624),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_715),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_696),
.B(n_663),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_813),
.B(n_624),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_733),
.A2(n_647),
.B(n_663),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_737),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_762),
.B(n_640),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_762),
.B(n_640),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_752),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_793),
.A2(n_665),
.B1(n_663),
.B2(n_682),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_734),
.A2(n_665),
.B(n_622),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_718),
.A2(n_741),
.B(n_735),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_718),
.A2(n_665),
.B(n_622),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_803),
.B(n_653),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_701),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_741),
.A2(n_638),
.B(n_622),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_768),
.B(n_724),
.Y(n_902)
);

BUFx4f_ASAP7_75t_L g903 ( 
.A(n_721),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_836),
.A2(n_638),
.B(n_662),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_836),
.A2(n_638),
.B(n_662),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_738),
.B(n_687),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_757),
.A2(n_795),
.B(n_780),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_731),
.B(n_664),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_726),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_726),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_818),
.A2(n_674),
.B(n_646),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_756),
.B(n_682),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_767),
.B(n_653),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_753),
.B(n_685),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_712),
.A2(n_691),
.B(n_646),
.C(n_676),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_743),
.B(n_577),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_794),
.B(n_650),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_851),
.A2(n_676),
.B(n_674),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_819),
.B(n_577),
.Y(n_919)
);

OAI321xp33_ASAP7_75t_L g920 ( 
.A1(n_807),
.A2(n_340),
.A3(n_306),
.B1(n_476),
.B2(n_330),
.C(n_235),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_773),
.B(n_678),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_776),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_828),
.A2(n_659),
.B1(n_598),
.B2(n_577),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_799),
.B(n_577),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_785),
.B(n_791),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_705),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_781),
.B(n_598),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_772),
.Y(n_928)
);

OR2x6_ASAP7_75t_SL g929 ( 
.A(n_796),
.B(n_634),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_802),
.B(n_598),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_753),
.B(n_330),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_772),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_709),
.A2(n_689),
.B(n_221),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_788),
.A2(n_330),
.B1(n_689),
.B2(n_594),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_740),
.B(n_754),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_705),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_714),
.A2(n_295),
.B(n_355),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_805),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_723),
.A2(n_283),
.B(n_351),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_748),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_782),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_740),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_747),
.A2(n_282),
.B(n_350),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_750),
.A2(n_277),
.B(n_349),
.Y(n_944)
);

OAI21xp33_ASAP7_75t_L g945 ( 
.A1(n_770),
.A2(n_326),
.B(n_252),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_760),
.A2(n_272),
.B(n_348),
.C(n_339),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_777),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_777),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_770),
.B(n_783),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_760),
.B(n_841),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_821),
.A2(n_262),
.B(n_333),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_824),
.A2(n_260),
.B(n_329),
.Y(n_952)
);

BUFx8_ASAP7_75t_L g953 ( 
.A(n_782),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_766),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_827),
.A2(n_258),
.B(n_327),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_778),
.A2(n_790),
.B(n_787),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_843),
.B(n_594),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_740),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_823),
.B(n_222),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_817),
.A2(n_321),
.B(n_318),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_778),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_825),
.A2(n_317),
.B(n_313),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_812),
.A2(n_266),
.B(n_21),
.C(n_24),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_829),
.A2(n_310),
.B(n_308),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_837),
.B(n_20),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_827),
.A2(n_305),
.B(n_304),
.Y(n_966)
);

O2A1O1Ixp5_ASAP7_75t_L g967 ( 
.A1(n_746),
.A2(n_26),
.B(n_30),
.C(n_33),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_807),
.A2(n_255),
.B1(n_250),
.B2(n_244),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_783),
.B(n_801),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_787),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_801),
.B(n_30),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_795),
.A2(n_804),
.B(n_847),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_831),
.A2(n_242),
.B(n_236),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_749),
.B(n_230),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_844),
.A2(n_227),
.B(n_225),
.Y(n_975)
);

NAND2x1_ASAP7_75t_L g976 ( 
.A(n_771),
.B(n_80),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_790),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_759),
.B(n_223),
.Y(n_978)
);

NOR2x1_ASAP7_75t_R g979 ( 
.A(n_849),
.B(n_34),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_754),
.B(n_34),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_814),
.A2(n_37),
.B(n_39),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_755),
.B(n_816),
.C(n_703),
.Y(n_982)
);

AO22x1_ASAP7_75t_L g983 ( 
.A1(n_758),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_761),
.B(n_46),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_774),
.Y(n_985)
);

AO22x1_ASAP7_75t_L g986 ( 
.A1(n_748),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_746),
.A2(n_91),
.B(n_161),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_832),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_754),
.B(n_48),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_763),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_765),
.B(n_53),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_765),
.B(n_53),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_784),
.A2(n_54),
.B(n_58),
.C(n_59),
.Y(n_993)
);

OAI21xp33_ASAP7_75t_L g994 ( 
.A1(n_798),
.A2(n_60),
.B(n_62),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_769),
.B(n_60),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_L g996 ( 
.A(n_695),
.B(n_64),
.C(n_113),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_842),
.A2(n_164),
.B(n_64),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_769),
.B(n_775),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_774),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_847),
.A2(n_808),
.B(n_800),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_833),
.B(n_834),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_816),
.A2(n_708),
.B(n_713),
.C(n_764),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_838),
.B(n_830),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_719),
.A2(n_789),
.B1(n_792),
.B2(n_797),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_708),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_697),
.A2(n_713),
.B(n_784),
.C(n_771),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_839),
.A2(n_697),
.B(n_704),
.Y(n_1007)
);

AO22x1_ASAP7_75t_L g1008 ( 
.A1(n_745),
.A2(n_822),
.B1(n_806),
.B2(n_850),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_704),
.A2(n_848),
.B(n_845),
.Y(n_1009)
);

AO21x1_ASAP7_75t_L g1010 ( 
.A1(n_736),
.A2(n_803),
.B(n_719),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_744),
.A2(n_809),
.B(n_702),
.C(n_846),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_815),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_815),
.A2(n_820),
.B(n_803),
.C(n_846),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_846),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_815),
.B(n_820),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_820),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_803),
.A2(n_739),
.B(n_725),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_716),
.A2(n_728),
.B(n_700),
.C(n_699),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_699),
.A2(n_700),
.B1(n_739),
.B2(n_722),
.Y(n_1019)
);

BUFx8_ASAP7_75t_L g1020 ( 
.A(n_859),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_867),
.B(n_949),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_935),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_949),
.B(n_902),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_971),
.A2(n_969),
.B(n_1018),
.C(n_852),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_953),
.Y(n_1025)
);

AOI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_931),
.A2(n_1001),
.B(n_954),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_931),
.A2(n_1001),
.B(n_954),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_897),
.A2(n_893),
.B(n_892),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_894),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_950),
.B(n_866),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_884),
.A2(n_972),
.B(n_918),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_856),
.A2(n_1005),
.B1(n_888),
.B2(n_925),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_SL g1033 ( 
.A1(n_984),
.A2(n_873),
.B(n_995),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_883),
.A2(n_868),
.B(n_870),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1005),
.A2(n_1006),
.B(n_855),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_866),
.B(n_857),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_L g1037 ( 
.A(n_878),
.B(n_941),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_896),
.A2(n_858),
.B(n_874),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_1009),
.A2(n_905),
.B(n_904),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_936),
.B(n_917),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_926),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_935),
.B(n_942),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_901),
.A2(n_888),
.B(n_898),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_936),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_853),
.A2(n_880),
.B1(n_914),
.B2(n_863),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_1006),
.A2(n_994),
.B(n_981),
.C(n_993),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_861),
.B(n_965),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_853),
.B(n_885),
.Y(n_1048)
);

OA22x2_ASAP7_75t_L g1049 ( 
.A1(n_935),
.A2(n_1016),
.B1(n_1015),
.B2(n_940),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_922),
.B(n_938),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_940),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_862),
.A2(n_978),
.B1(n_934),
.B2(n_982),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_899),
.A2(n_879),
.B(n_890),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_990),
.B(n_1003),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_862),
.A2(n_934),
.B1(n_912),
.B2(n_889),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_990),
.B(n_1003),
.Y(n_1057)
);

NOR2x1_ASAP7_75t_SL g1058 ( 
.A(n_865),
.B(n_882),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_923),
.A2(n_876),
.B(n_976),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_909),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_910),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_865),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_958),
.B(n_913),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_913),
.B(n_974),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1012),
.B(n_871),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_886),
.A2(n_930),
.B1(n_860),
.B2(n_946),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_988),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_881),
.A2(n_1004),
.B(n_864),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1012),
.B(n_980),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_906),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_953),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1008),
.B(n_914),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_895),
.A2(n_998),
.B(n_939),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_928),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_937),
.A2(n_966),
.B(n_955),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_903),
.A2(n_887),
.B1(n_968),
.B2(n_908),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_943),
.A2(n_944),
.B(n_964),
.Y(n_1077)
);

AOI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_921),
.B(n_1013),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_932),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_973),
.A2(n_960),
.B(n_962),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_952),
.A2(n_957),
.B(n_1014),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_924),
.A2(n_927),
.B(n_887),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_947),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_991),
.B(n_992),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_872),
.B(n_875),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_996),
.A2(n_980),
.B(n_989),
.C(n_967),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_989),
.A2(n_1016),
.B1(n_919),
.B2(n_903),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1010),
.A2(n_997),
.B(n_933),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_948),
.Y(n_1089)
);

OA22x2_ASAP7_75t_L g1090 ( 
.A1(n_929),
.A2(n_900),
.B1(n_959),
.B2(n_916),
.Y(n_1090)
);

AOI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_920),
.A2(n_963),
.B(n_977),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_865),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_882),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_891),
.B(n_986),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_961),
.A2(n_970),
.B(n_985),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_891),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1011),
.B(n_877),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_877),
.B(n_985),
.Y(n_1098)
);

AO21x1_ASAP7_75t_L g1099 ( 
.A1(n_987),
.A2(n_975),
.B(n_951),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_983),
.B(n_967),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_882),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_854),
.A2(n_882),
.B(n_999),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_999),
.Y(n_1103)
);

AO21x2_ASAP7_75t_L g1104 ( 
.A1(n_999),
.A2(n_1009),
.B(n_1002),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_979),
.B(n_867),
.Y(n_1105)
);

AND2x6_ASAP7_75t_L g1106 ( 
.A(n_865),
.B(n_854),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1005),
.A2(n_751),
.B(n_1006),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_867),
.B(n_949),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_935),
.B(n_722),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_867),
.B(n_949),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1019),
.A2(n_1007),
.B(n_1017),
.Y(n_1113)
);

O2A1O1Ixp5_ASAP7_75t_L g1114 ( 
.A1(n_1019),
.A2(n_869),
.B(n_971),
.C(n_1017),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1005),
.A2(n_751),
.B(n_1006),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_954),
.B(n_729),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_872),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_865),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_SL g1122 ( 
.A1(n_971),
.A2(n_1018),
.B1(n_728),
.B2(n_716),
.C(n_558),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_971),
.A2(n_949),
.B(n_751),
.C(n_856),
.Y(n_1123)
);

CKINVDCx14_ASAP7_75t_R g1124 ( 
.A(n_872),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_971),
.A2(n_949),
.B(n_751),
.C(n_856),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_935),
.B(n_722),
.Y(n_1126)
);

BUFx2_ASAP7_75t_SL g1127 ( 
.A(n_941),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_956),
.A2(n_907),
.B(n_911),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_971),
.A2(n_949),
.B(n_751),
.C(n_856),
.Y(n_1130)
);

AO21x2_ASAP7_75t_L g1131 ( 
.A1(n_1009),
.A2(n_1002),
.B(n_1000),
.Y(n_1131)
);

O2A1O1Ixp5_ASAP7_75t_L g1132 ( 
.A1(n_1019),
.A2(n_869),
.B(n_971),
.C(n_1017),
.Y(n_1132)
);

AOI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_949),
.A2(n_589),
.B(n_826),
.Y(n_1133)
);

AOI221xp5_ASAP7_75t_SL g1134 ( 
.A1(n_971),
.A2(n_1018),
.B1(n_728),
.B2(n_716),
.C(n_558),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_953),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1019),
.A2(n_1013),
.B(n_865),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_867),
.B(n_949),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_872),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_865),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_L g1146 ( 
.A(n_865),
.B(n_592),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_872),
.Y(n_1147)
);

AOI221x1_ASAP7_75t_L g1148 ( 
.A1(n_996),
.A2(n_971),
.B1(n_994),
.B2(n_1019),
.C(n_981),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_926),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_865),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_956),
.A2(n_907),
.B(n_911),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_956),
.A2(n_907),
.B(n_911),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1002),
.A2(n_1019),
.A3(n_1010),
.B(n_915),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1017),
.A2(n_897),
.B(n_1019),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_867),
.B(n_949),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_956),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_SL g1157 ( 
.A1(n_1010),
.A2(n_950),
.B(n_883),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_1080),
.A2(n_1077),
.B(n_1075),
.C(n_1024),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1029),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1021),
.B(n_1110),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1112),
.A2(n_1139),
.B1(n_1155),
.B2(n_1053),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1041),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1023),
.B(n_1030),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1040),
.B(n_1116),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1036),
.B(n_1123),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1133),
.A2(n_1090),
.B1(n_1026),
.B2(n_1027),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1123),
.A2(n_1125),
.B1(n_1130),
.B2(n_1086),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_SL g1168 ( 
.A(n_1071),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1105),
.B(n_1045),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_SL g1170 ( 
.A(n_1120),
.B(n_1141),
.Y(n_1170)
);

AO21x1_ASAP7_75t_L g1171 ( 
.A1(n_1032),
.A2(n_1066),
.B(n_1097),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1050),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1125),
.A2(n_1130),
.B(n_1043),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1044),
.B(n_1069),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1086),
.A2(n_1047),
.B1(n_1046),
.B2(n_1109),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1028),
.A2(n_1108),
.B(n_1107),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1117),
.A2(n_1143),
.B(n_1140),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1044),
.B(n_1051),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1148),
.B(n_1046),
.C(n_1068),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1020),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1048),
.B(n_1149),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1118),
.A2(n_1142),
.B(n_1138),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1111),
.B(n_1126),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1119),
.A2(n_1144),
.B(n_1136),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1020),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1111),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1111),
.B(n_1126),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1067),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1020),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1072),
.B(n_1051),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1128),
.A2(n_1154),
.B(n_1034),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1055),
.B(n_1057),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1087),
.B(n_1084),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1074),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1126),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1096),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1085),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1065),
.B(n_1022),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1085),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1122),
.B(n_1134),
.C(n_1115),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1070),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1127),
.Y(n_1202)
);

OR2x6_ASAP7_75t_L g1203 ( 
.A(n_1042),
.B(n_1090),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1114),
.A2(n_1132),
.B(n_1038),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1042),
.B(n_1037),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1042),
.Y(n_1206)
);

OAI21xp33_ASAP7_75t_L g1207 ( 
.A1(n_1100),
.A2(n_1064),
.B(n_1035),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1120),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1056),
.A2(n_1146),
.B1(n_1070),
.B2(n_1094),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1141),
.B(n_1147),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1025),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1058),
.B(n_1052),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1063),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1079),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1071),
.B(n_1049),
.Y(n_1215)
);

CKINVDCx6p67_ASAP7_75t_R g1216 ( 
.A(n_1025),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1096),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1083),
.Y(n_1218)
);

OR2x6_ASAP7_75t_L g1219 ( 
.A(n_1049),
.B(n_1135),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_1106),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1039),
.A2(n_1054),
.B(n_1146),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1060),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1103),
.Y(n_1223)
);

BUFx8_ASAP7_75t_SL g1224 ( 
.A(n_1147),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1060),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1106),
.Y(n_1226)
);

NOR2xp67_ASAP7_75t_SL g1227 ( 
.A(n_1093),
.B(n_1150),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1076),
.A2(n_1098),
.B1(n_1073),
.B2(n_1137),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1061),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1124),
.B(n_1103),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1089),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1089),
.B(n_1157),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1093),
.Y(n_1233)
);

INVx5_ASAP7_75t_L g1234 ( 
.A(n_1106),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1078),
.A2(n_1081),
.B1(n_1082),
.B2(n_1091),
.Y(n_1235)
);

NAND2xp33_ASAP7_75t_L g1236 ( 
.A(n_1106),
.B(n_1093),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1124),
.A2(n_1131),
.B(n_1099),
.C(n_1101),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1052),
.B(n_1121),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1062),
.B(n_1092),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1095),
.Y(n_1240)
);

INVxp67_ASAP7_75t_L g1241 ( 
.A(n_1121),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1121),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1106),
.B(n_1150),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1145),
.B(n_1153),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1145),
.B(n_1102),
.Y(n_1245)
);

CKINVDCx8_ASAP7_75t_R g1246 ( 
.A(n_1145),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1104),
.B(n_1153),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1104),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1153),
.B(n_1131),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1153),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1156),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1059),
.B(n_1031),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1129),
.A2(n_1152),
.B(n_1151),
.Y(n_1253)
);

INVx5_ASAP7_75t_L g1254 ( 
.A(n_1033),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1088),
.B(n_1113),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1021),
.A2(n_1110),
.B1(n_1139),
.B2(n_1112),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1111),
.B(n_1126),
.Y(n_1257)
);

AOI211xp5_ASAP7_75t_L g1258 ( 
.A1(n_1133),
.A2(n_949),
.B(n_971),
.C(n_866),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_1020),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1041),
.B(n_1149),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1123),
.A2(n_1130),
.B(n_1125),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1021),
.B(n_1110),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1021),
.B(n_1110),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1021),
.B(n_1110),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1041),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1029),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1020),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1111),
.B(n_1126),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1111),
.B(n_1126),
.Y(n_1269)
);

INVx5_ASAP7_75t_L g1270 ( 
.A(n_1096),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1041),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1020),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1041),
.Y(n_1273)
);

BUFx8_ASAP7_75t_SL g1274 ( 
.A(n_1025),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1123),
.A2(n_1130),
.B(n_1125),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1123),
.A2(n_1130),
.B(n_1125),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1020),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1029),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1085),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1107),
.A2(n_1117),
.B(n_1108),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1020),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1096),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1021),
.B(n_1110),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1029),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1111),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1029),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_1120),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1107),
.A2(n_1117),
.B(n_1108),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1020),
.Y(n_1289)
);

INVx5_ASAP7_75t_L g1290 ( 
.A(n_1096),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1020),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1052),
.B(n_1062),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1111),
.B(n_1126),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1021),
.B(n_1110),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1123),
.A2(n_1130),
.B(n_1125),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1021),
.B(n_1110),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1220),
.B(n_1226),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1226),
.B(n_1234),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1199),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1203),
.B(n_1215),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1258),
.A2(n_1256),
.B(n_1161),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1178),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1244),
.B(n_1250),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1274),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1224),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1191),
.A2(n_1182),
.B(n_1177),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1255),
.A2(n_1235),
.B(n_1221),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_SL g1308 ( 
.A(n_1197),
.B(n_1279),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1266),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1260),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1278),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1183),
.B(n_1187),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1284),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1169),
.A2(n_1167),
.B1(n_1193),
.B2(n_1203),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1286),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1203),
.A2(n_1166),
.B1(n_1215),
.B2(n_1167),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1249),
.B(n_1174),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1188),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1164),
.B(n_1261),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1179),
.A2(n_1256),
.B1(n_1175),
.B2(n_1215),
.Y(n_1320)
);

AO21x1_ASAP7_75t_L g1321 ( 
.A1(n_1258),
.A2(n_1175),
.B(n_1295),
.Y(n_1321)
);

OAI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1161),
.A2(n_1209),
.B1(n_1163),
.B2(n_1262),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1179),
.A2(n_1165),
.B1(n_1276),
.B2(n_1275),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1194),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1257),
.B(n_1293),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1251),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1214),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1218),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1222),
.Y(n_1329)
);

BUFx10_ASAP7_75t_L g1330 ( 
.A(n_1210),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1219),
.A2(n_1171),
.B1(n_1181),
.B2(n_1209),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1225),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1184),
.A2(n_1176),
.B(n_1204),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1229),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1165),
.B(n_1190),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1231),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1172),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1219),
.A2(n_1296),
.B1(n_1160),
.B2(n_1283),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1219),
.A2(n_1296),
.B1(n_1160),
.B2(n_1283),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1247),
.B(n_1207),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1264),
.B(n_1263),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1246),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1263),
.A2(n_1294),
.B1(n_1173),
.B2(n_1192),
.Y(n_1343)
);

AO21x1_ASAP7_75t_L g1344 ( 
.A1(n_1235),
.A2(n_1228),
.B(n_1237),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1213),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1216),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1247),
.B(n_1223),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1230),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1201),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1294),
.B(n_1208),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1234),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1232),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1206),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1238),
.Y(n_1354)
);

INVx8_ASAP7_75t_L g1355 ( 
.A(n_1168),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1271),
.A2(n_1273),
.B1(n_1200),
.B2(n_1162),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1252),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1211),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1198),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1205),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1248),
.A2(n_1158),
.B(n_1240),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1162),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1238),
.Y(n_1363)
);

AOI222xp33_ASAP7_75t_L g1364 ( 
.A1(n_1200),
.A2(n_1265),
.B1(n_1205),
.B2(n_1168),
.C1(n_1228),
.C2(n_1202),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1252),
.A2(n_1253),
.B(n_1227),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1253),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1202),
.B(n_1257),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1292),
.A2(n_1241),
.B(n_1254),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1245),
.B(n_1242),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1254),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1293),
.B(n_1285),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1233),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1242),
.Y(n_1373)
);

BUFx2_ASAP7_75t_R g1374 ( 
.A(n_1180),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1280),
.A2(n_1288),
.B(n_1243),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1233),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1239),
.Y(n_1377)
);

INVxp33_ASAP7_75t_L g1378 ( 
.A(n_1186),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1195),
.A2(n_1189),
.B1(n_1281),
.B2(n_1289),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1195),
.A2(n_1259),
.B1(n_1185),
.B2(n_1267),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1238),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1287),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1268),
.B(n_1269),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1212),
.B(n_1272),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1236),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1291),
.A2(n_1277),
.B1(n_1170),
.B2(n_1196),
.Y(n_1386)
);

AO21x1_ASAP7_75t_SL g1387 ( 
.A1(n_1212),
.A2(n_1270),
.B(n_1282),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1287),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1217),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1290),
.A2(n_1191),
.B(n_1182),
.Y(n_1390)
);

AO21x1_ASAP7_75t_L g1391 ( 
.A1(n_1196),
.A2(n_1167),
.B(n_1258),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1290),
.A2(n_1133),
.B1(n_703),
.B2(n_826),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1159),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1159),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1274),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1220),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1258),
.A2(n_949),
.B1(n_1110),
.B2(n_1021),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1178),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1274),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1159),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1250),
.B(n_1249),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1199),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1169),
.A2(n_1133),
.B1(n_703),
.B2(n_826),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1251),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1244),
.B(n_1178),
.Y(n_1405)
);

BUFx8_ASAP7_75t_SL g1406 ( 
.A(n_1274),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_SL g1407 ( 
.A1(n_1171),
.A2(n_1275),
.B(n_1261),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1250),
.B(n_1249),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1258),
.A2(n_1133),
.B(n_1125),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1251),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1159),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1159),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1159),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1244),
.B(n_1178),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1169),
.B(n_591),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1169),
.A2(n_1133),
.B1(n_703),
.B2(n_826),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1159),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1199),
.Y(n_1418)
);

BUFx8_ASAP7_75t_L g1419 ( 
.A(n_1168),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1159),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1349),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1405),
.B(n_1414),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1322),
.B(n_1314),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1366),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1302),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1357),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1307),
.A2(n_1344),
.B(n_1365),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1357),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1395),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1352),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1405),
.B(n_1414),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1329),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1335),
.B(n_1341),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1332),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1415),
.B(n_1350),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1344),
.A2(n_1390),
.B(n_1391),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1390),
.Y(n_1437)
);

AOI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1390),
.A2(n_1391),
.B(n_1333),
.Y(n_1438)
);

CKINVDCx6p67_ASAP7_75t_R g1439 ( 
.A(n_1395),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1334),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1317),
.B(n_1319),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1336),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1299),
.B(n_1402),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1317),
.B(n_1319),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1403),
.A2(n_1416),
.B1(n_1316),
.B2(n_1301),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1401),
.B(n_1408),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1340),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1340),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1303),
.B(n_1335),
.Y(n_1449)
);

OAI21xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1409),
.A2(n_1331),
.B(n_1364),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1407),
.A2(n_1321),
.B(n_1375),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1303),
.B(n_1398),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1347),
.B(n_1369),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1420),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1347),
.B(n_1401),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1362),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1361),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1408),
.B(n_1309),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1361),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1361),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1333),
.A2(n_1306),
.B(n_1370),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1343),
.B(n_1359),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1311),
.B(n_1313),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1315),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1318),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1397),
.B(n_1320),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1393),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1394),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1400),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1411),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1321),
.A2(n_1306),
.B(n_1323),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1345),
.B(n_1337),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1412),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1413),
.B(n_1417),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1324),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1327),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1372),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1328),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1376),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1299),
.B(n_1402),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1353),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1418),
.B(n_1308),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1348),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1418),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1392),
.A2(n_1356),
.B(n_1368),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1373),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1381),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1360),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1300),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1385),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1377),
.A2(n_1367),
.B(n_1371),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1355),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1300),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1326),
.B(n_1404),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1354),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1326),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1363),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1410),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1351),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1351),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1351),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1396),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1396),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1410),
.B(n_1339),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1338),
.A2(n_1297),
.B(n_1298),
.Y(n_1505)
);

INVxp33_ASAP7_75t_L g1506 ( 
.A(n_1312),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1310),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1441),
.B(n_1330),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1432),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1477),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1435),
.B(n_1330),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1432),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1446),
.B(n_1355),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1434),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1433),
.B(n_1330),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1424),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1434),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1449),
.B(n_1355),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1444),
.B(n_1384),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1422),
.B(n_1325),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1440),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1449),
.B(n_1389),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1425),
.B(n_1389),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1422),
.B(n_1325),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_SL g1526 ( 
.A(n_1466),
.B(n_1383),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1447),
.B(n_1386),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1431),
.B(n_1453),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1431),
.B(n_1325),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1453),
.B(n_1312),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1448),
.B(n_1342),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1458),
.B(n_1382),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1450),
.A2(n_1445),
.B1(n_1471),
.B2(n_1462),
.C(n_1504),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1458),
.B(n_1382),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1452),
.B(n_1387),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1452),
.B(n_1387),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1440),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_1380),
.B2(n_1379),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1484),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1455),
.B(n_1448),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1442),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1421),
.B(n_1419),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1426),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1430),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1430),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1481),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1456),
.B(n_1419),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1483),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1496),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1426),
.B(n_1358),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1498),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1428),
.B(n_1358),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1428),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1463),
.B(n_1474),
.Y(n_1555)
);

CKINVDCx16_ASAP7_75t_R g1556 ( 
.A(n_1429),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1498),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1454),
.B(n_1378),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1464),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1534),
.B(n_1450),
.C(n_1490),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1511),
.A2(n_1485),
.B1(n_1482),
.B2(n_1480),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1552),
.B(n_1490),
.C(n_1504),
.Y(n_1562)
);

OAI21xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1517),
.A2(n_1443),
.B(n_1494),
.Y(n_1563)
);

NAND4xp25_ASAP7_75t_L g1564 ( 
.A(n_1515),
.B(n_1494),
.C(n_1486),
.D(n_1478),
.Y(n_1564)
);

OAI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1539),
.A2(n_1436),
.B1(n_1506),
.B2(n_1505),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1526),
.A2(n_1472),
.B1(n_1478),
.B2(n_1468),
.C(n_1464),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1540),
.B(n_1436),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1539),
.A2(n_1438),
.B(n_1427),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_L g1569 ( 
.A(n_1557),
.B(n_1495),
.C(n_1497),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_L g1570 ( 
.A(n_1547),
.B(n_1495),
.C(n_1497),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_SL g1571 ( 
.A(n_1524),
.B(n_1346),
.C(n_1399),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1510),
.B(n_1465),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1550),
.B(n_1486),
.C(n_1467),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1532),
.B(n_1465),
.Y(n_1574)
);

NOR3xp33_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1427),
.C(n_1460),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1526),
.A2(n_1505),
.B1(n_1437),
.B2(n_1493),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1508),
.B(n_1468),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1555),
.B(n_1451),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1526),
.A2(n_1437),
.B1(n_1493),
.B2(n_1489),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1451),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1508),
.B(n_1469),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1451),
.Y(n_1582)
);

AND4x1_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1406),
.C(n_1439),
.D(n_1374),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1541),
.B(n_1451),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1549),
.B(n_1470),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1558),
.B(n_1473),
.C(n_1475),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1545),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1536),
.A2(n_1492),
.B(n_1499),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1545),
.B(n_1546),
.Y(n_1589)
);

OAI21xp33_ASAP7_75t_L g1590 ( 
.A1(n_1527),
.A2(n_1438),
.B(n_1460),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1546),
.B(n_1475),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1509),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1521),
.B(n_1476),
.Y(n_1593)
);

NAND3xp33_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1487),
.C(n_1457),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1516),
.A2(n_1461),
.B(n_1459),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1521),
.B(n_1507),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1520),
.B(n_1500),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1520),
.B(n_1500),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1525),
.B(n_1491),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1525),
.B(n_1491),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1519),
.A2(n_1439),
.B1(n_1492),
.B2(n_1346),
.Y(n_1601)
);

OAI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1509),
.A2(n_1457),
.B(n_1503),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1531),
.B(n_1487),
.C(n_1502),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1529),
.B(n_1491),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1529),
.B(n_1491),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1512),
.B(n_1488),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1512),
.B(n_1488),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1514),
.B(n_1501),
.Y(n_1608)
);

OAI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1514),
.A2(n_1559),
.B(n_1522),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1599),
.B(n_1544),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1578),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1530),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1578),
.B(n_1518),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1582),
.B(n_1530),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1600),
.B(n_1544),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1570),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1592),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1582),
.B(n_1554),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1595),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1609),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1608),
.Y(n_1622)
);

CKINVDCx14_ASAP7_75t_R g1623 ( 
.A(n_1571),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1584),
.B(n_1518),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1591),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1606),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1607),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1587),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1595),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1586),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1572),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1595),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1574),
.Y(n_1633)
);

NOR2xp67_ASAP7_75t_L g1634 ( 
.A(n_1588),
.B(n_1437),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1604),
.B(n_1522),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1585),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1605),
.B(n_1538),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1573),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1567),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1575),
.B(n_1538),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1567),
.Y(n_1641)
);

INVx4_ASAP7_75t_R g1642 ( 
.A(n_1597),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1596),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1594),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1597),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1602),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1617),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1619),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1634),
.B(n_1569),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1617),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1646),
.B(n_1577),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1612),
.B(n_1563),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1622),
.Y(n_1654)
);

NOR2xp67_ASAP7_75t_L g1655 ( 
.A(n_1634),
.B(n_1562),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1643),
.Y(n_1656)
);

NOR2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1560),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1612),
.B(n_1598),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1622),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1619),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1612),
.B(n_1598),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1625),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1625),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1626),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1626),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1616),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1614),
.B(n_1577),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1619),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1614),
.B(n_1536),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1638),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1630),
.B(n_1593),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1616),
.B(n_1561),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1630),
.B(n_1581),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1627),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1621),
.Y(n_1676)
);

BUFx3_ASAP7_75t_L g1677 ( 
.A(n_1639),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1646),
.B(n_1564),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1638),
.B(n_1566),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1629),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1614),
.B(n_1537),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1621),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1629),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_L g1684 ( 
.A(n_1640),
.B(n_1551),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1624),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1645),
.B(n_1537),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1636),
.B(n_1542),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1624),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1645),
.B(n_1551),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1648),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1648),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1666),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1651),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1651),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1672),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1672),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1674),
.Y(n_1697)
);

OAI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1679),
.A2(n_1620),
.B(n_1641),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1657),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1674),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1657),
.A2(n_1644),
.B1(n_1565),
.B2(n_1647),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1653),
.B(n_1641),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1653),
.B(n_1645),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1687),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1655),
.B(n_1639),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1620),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1673),
.B(n_1655),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1678),
.B(n_1647),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1678),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1662),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1650),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1667),
.B(n_1645),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1649),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1650),
.A2(n_1623),
.B(n_1644),
.C(n_1576),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.B(n_1640),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1662),
.Y(n_1716)
);

NOR3xp33_ASAP7_75t_SL g1717 ( 
.A(n_1652),
.B(n_1556),
.C(n_1399),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1663),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1663),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1656),
.B(n_1635),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1664),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1667),
.B(n_1636),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1664),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1650),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1684),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1665),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1665),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1685),
.B(n_1635),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1684),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1685),
.B(n_1643),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1671),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1671),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1677),
.B(n_1623),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1708),
.B(n_1688),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1692),
.B(n_1675),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1699),
.B(n_1675),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1708),
.B(n_1688),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1701),
.A2(n_1568),
.B1(n_1590),
.B2(n_1683),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1721),
.Y(n_1740)
);

NOR2x1_ASAP7_75t_L g1741 ( 
.A(n_1707),
.B(n_1677),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1709),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1701),
.A2(n_1660),
.B1(n_1680),
.B2(n_1683),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1690),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1698),
.A2(n_1677),
.B1(n_1639),
.B2(n_1683),
.C(n_1668),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1720),
.B(n_1676),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1713),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1691),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1713),
.Y(n_1749)
);

CKINVDCx16_ASAP7_75t_R g1750 ( 
.A(n_1699),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1706),
.B(n_1676),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1693),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1720),
.B(n_1682),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1703),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1734),
.A2(n_1660),
.B1(n_1649),
.B2(n_1668),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1715),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1715),
.B(n_1406),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1705),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1703),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1705),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1694),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1702),
.B(n_1669),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1729),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1710),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1714),
.A2(n_1682),
.B(n_1659),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1712),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1734),
.A2(n_1611),
.B1(n_1649),
.B2(n_1660),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1714),
.B(n_1659),
.C(n_1654),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1705),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1712),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1711),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1695),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1739),
.A2(n_1724),
.B1(n_1711),
.B2(n_1704),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1750),
.B(n_1556),
.Y(n_1774)
);

AOI21xp33_ASAP7_75t_L g1775 ( 
.A1(n_1768),
.A2(n_1724),
.B(n_1725),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1742),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1744),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1763),
.B(n_1696),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_SL g1779 ( 
.A(n_1768),
.B(n_1743),
.C(n_1765),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1771),
.B(n_1760),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1771),
.B(n_1697),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1750),
.B(n_1304),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1741),
.A2(n_1700),
.B1(n_1702),
.B2(n_1730),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1755),
.A2(n_1680),
.B1(n_1668),
.B2(n_1731),
.C(n_1732),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1744),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1762),
.B(n_1717),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1760),
.B(n_1722),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1736),
.B(n_1728),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1748),
.Y(n_1789)
);

NAND3xp33_ASAP7_75t_SL g1790 ( 
.A(n_1745),
.B(n_1304),
.C(n_1733),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1748),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1752),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1752),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1741),
.A2(n_1733),
.B(n_1583),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1758),
.Y(n_1795)
);

NOR3xp33_ASAP7_75t_L g1796 ( 
.A(n_1758),
.B(n_1718),
.C(n_1716),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1761),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1761),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1795),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1777),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1776),
.B(n_1760),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1779),
.B(n_1757),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1785),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1789),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1779),
.B(n_1758),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1782),
.B(n_1762),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1773),
.A2(n_1769),
.B1(n_1767),
.B2(n_1749),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1780),
.B(n_1769),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1774),
.B(n_1758),
.Y(n_1809)
);

NAND2x1_ASAP7_75t_L g1810 ( 
.A(n_1786),
.B(n_1759),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1791),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1778),
.Y(n_1812)
);

NAND2x1_ASAP7_75t_L g1813 ( 
.A(n_1783),
.B(n_1759),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1794),
.B(n_1769),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1788),
.B(n_1759),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1772),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1796),
.B(n_1740),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1792),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1805),
.A2(n_1775),
.B(n_1793),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1802),
.A2(n_1790),
.B1(n_1787),
.B2(n_1784),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1805),
.A2(n_1796),
.B1(n_1790),
.B2(n_1798),
.C(n_1797),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1812),
.B(n_1781),
.Y(n_1822)
);

O2A1O1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1817),
.A2(n_1740),
.B(n_1737),
.C(n_1738),
.Y(n_1823)
);

NAND4xp75_ASAP7_75t_L g1824 ( 
.A(n_1814),
.B(n_1747),
.C(n_1749),
.D(n_1754),
.Y(n_1824)
);

OAI211xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1802),
.A2(n_1754),
.B(n_1766),
.C(n_1770),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1816),
.B(n_1766),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_R g1827 ( 
.A(n_1809),
.B(n_1305),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1807),
.A2(n_1751),
.B1(n_1764),
.B2(n_1749),
.C(n_1747),
.Y(n_1828)
);

OAI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1807),
.A2(n_1735),
.B1(n_1738),
.B2(n_1753),
.C(n_1746),
.Y(n_1829)
);

OAI211xp5_ASAP7_75t_L g1830 ( 
.A1(n_1813),
.A2(n_1770),
.B(n_1388),
.C(n_1764),
.Y(n_1830)
);

AO22x2_ASAP7_75t_L g1831 ( 
.A1(n_1824),
.A2(n_1799),
.B1(n_1810),
.B2(n_1811),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1822),
.B(n_1800),
.Y(n_1832)
);

NAND4xp75_ASAP7_75t_L g1833 ( 
.A(n_1819),
.B(n_1809),
.C(n_1801),
.D(n_1808),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_L g1834 ( 
.A(n_1825),
.B(n_1803),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1826),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1828),
.B(n_1815),
.Y(n_1836)
);

NOR2xp67_ASAP7_75t_L g1837 ( 
.A(n_1830),
.B(n_1806),
.Y(n_1837)
);

OA22x2_ASAP7_75t_L g1838 ( 
.A1(n_1820),
.A2(n_1804),
.B1(n_1818),
.B2(n_1827),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_L g1839 ( 
.A(n_1821),
.B(n_1829),
.C(n_1823),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1824),
.Y(n_1840)
);

AOI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1819),
.A2(n_1747),
.B(n_1735),
.Y(n_1841)
);

INVx1_ASAP7_75t_SL g1842 ( 
.A(n_1827),
.Y(n_1842)
);

OAI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1839),
.A2(n_1388),
.B(n_1305),
.C(n_1753),
.Y(n_1843)
);

NAND4xp25_ASAP7_75t_L g1844 ( 
.A(n_1837),
.B(n_1746),
.C(n_1727),
.D(n_1719),
.Y(n_1844)
);

NOR3xp33_ASAP7_75t_L g1845 ( 
.A(n_1840),
.B(n_1680),
.C(n_1723),
.Y(n_1845)
);

AOI21xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1831),
.A2(n_1726),
.B(n_1728),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1835),
.B(n_1658),
.Y(n_1847)
);

NOR3x1_ASAP7_75t_L g1848 ( 
.A(n_1833),
.B(n_1553),
.C(n_1601),
.Y(n_1848)
);

NOR3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1841),
.B(n_1836),
.C(n_1838),
.Y(n_1849)
);

INVx2_ASAP7_75t_SL g1850 ( 
.A(n_1847),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1834),
.B1(n_1832),
.B2(n_1842),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1848),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1846),
.B(n_1654),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1843),
.A2(n_1611),
.B1(n_1632),
.B2(n_1629),
.Y(n_1854)
);

BUFx6f_ASAP7_75t_L g1855 ( 
.A(n_1844),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1845),
.B(n_1628),
.Y(n_1856)
);

NOR2x1_ASAP7_75t_L g1857 ( 
.A(n_1852),
.B(n_1553),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1850),
.Y(n_1858)
);

AND2x4_ASAP7_75t_SL g1859 ( 
.A(n_1851),
.B(n_1689),
.Y(n_1859)
);

OAI311xp33_ASAP7_75t_L g1860 ( 
.A1(n_1854),
.A2(n_1856),
.A3(n_1855),
.B1(n_1853),
.C1(n_1535),
.Y(n_1860)
);

NAND4xp25_ASAP7_75t_L g1861 ( 
.A(n_1855),
.B(n_1689),
.C(n_1533),
.D(n_1686),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1851),
.A2(n_1628),
.B1(n_1633),
.B2(n_1631),
.Y(n_1862)
);

NOR3xp33_ASAP7_75t_L g1863 ( 
.A(n_1858),
.B(n_1632),
.C(n_1637),
.Y(n_1863)
);

NOR3xp33_ASAP7_75t_L g1864 ( 
.A(n_1857),
.B(n_1632),
.C(n_1637),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1859),
.A2(n_1633),
.B1(n_1631),
.B2(n_1669),
.Y(n_1865)
);

AND2x2_ASAP7_75t_SL g1866 ( 
.A(n_1860),
.B(n_1686),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1866),
.A2(n_1862),
.B1(n_1861),
.B2(n_1686),
.Y(n_1867)
);

NOR3xp33_ASAP7_75t_L g1868 ( 
.A(n_1867),
.B(n_1864),
.C(n_1865),
.Y(n_1868)
);

AO22x2_ASAP7_75t_L g1869 ( 
.A1(n_1868),
.A2(n_1863),
.B1(n_1681),
.B2(n_1611),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1868),
.A2(n_1681),
.B(n_1661),
.Y(n_1870)
);

OA21x2_ASAP7_75t_L g1871 ( 
.A1(n_1870),
.A2(n_1661),
.B(n_1658),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1869),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1872),
.A2(n_1613),
.B(n_1610),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1871),
.B(n_1613),
.Y(n_1874)
);

AO21x2_ASAP7_75t_L g1875 ( 
.A1(n_1873),
.A2(n_1871),
.B(n_1523),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1874),
.B1(n_1610),
.B2(n_1615),
.Y(n_1876)
);

OAI221xp5_ASAP7_75t_R g1877 ( 
.A1(n_1876),
.A2(n_1579),
.B1(n_1642),
.B2(n_1686),
.C(n_1618),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1615),
.B(n_1610),
.C(n_1513),
.Y(n_1878)
);


endmodule