module fake_jpeg_7181_n_249 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_18),
.B1(n_26),
.B2(n_20),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_40),
.B1(n_20),
.B2(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_18),
.B1(n_26),
.B2(n_20),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

OR2x4_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_14),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_20),
.Y(n_48)
);

FAx1_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_20),
.CI(n_14),
.CON(n_58),
.SN(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_63),
.CI(n_67),
.CON(n_85),
.SN(n_85)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_56),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_33),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_73),
.B1(n_18),
.B2(n_26),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_23),
.B(n_16),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_48),
.C(n_17),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_35),
.B1(n_51),
.B2(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_59),
.B1(n_76),
.B2(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_58),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_92),
.B1(n_23),
.B2(n_15),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_49),
.B1(n_47),
.B2(n_52),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_84),
.B1(n_91),
.B2(n_94),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_90),
.B1(n_58),
.B2(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_47),
.B1(n_55),
.B2(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_45),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_43),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_32),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_41),
.B1(n_35),
.B2(n_45),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_26),
.B1(n_38),
.B2(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_43),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_19),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_33),
.B1(n_17),
.B2(n_24),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_104),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_85),
.B(n_78),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_61),
.B1(n_76),
.B2(n_58),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_101),
.B1(n_81),
.B2(n_84),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_69),
.B1(n_66),
.B2(n_61),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_68),
.B1(n_17),
.B2(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_68),
.B1(n_31),
.B2(n_32),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_79),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_0),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_116),
.B(n_94),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_95),
.B(n_19),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_15),
.B1(n_16),
.B2(n_23),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_113),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_78),
.B1(n_89),
.B2(n_87),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_16),
.B1(n_11),
.B2(n_12),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_79),
.B(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_77),
.Y(n_122)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_121),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_112),
.B1(n_107),
.B2(n_103),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_128),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_129),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_109),
.B(n_21),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_92),
.B1(n_85),
.B2(n_91),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_110),
.B1(n_115),
.B2(n_106),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_85),
.C(n_92),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_109),
.C(n_21),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_135),
.B(n_137),
.Y(n_157)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_136),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_85),
.B(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_25),
.B(n_22),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_136),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_143),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_156),
.B1(n_159),
.B2(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_123),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_107),
.B1(n_106),
.B2(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_137),
.C(n_131),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_158),
.B(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_121),
.B1(n_120),
.B2(n_21),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_109),
.B1(n_19),
.B2(n_24),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_173),
.B1(n_178),
.B2(n_24),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_140),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_124),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_165),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_125),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_126),
.C(n_123),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_120),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_120),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_152),
.C(n_153),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_143),
.Y(n_181)
);

AOI22x1_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_141),
.B1(n_150),
.B2(n_158),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_134),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_146),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_185),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_142),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_187),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_159),
.B1(n_161),
.B2(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_190),
.B1(n_188),
.B2(n_187),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_167),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_145),
.B(n_151),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_191),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_156),
.B1(n_155),
.B2(n_139),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_174),
.B1(n_176),
.B2(n_169),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_108),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_194),
.C(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_57),
.C(n_70),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_173),
.CI(n_177),
.CON(n_196),
.SN(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_178),
.C(n_70),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_70),
.C(n_57),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_24),
.C(n_22),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_193),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_8),
.B1(n_7),
.B2(n_13),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_195),
.B1(n_200),
.B2(n_12),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_8),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_207),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_8),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_196),
.B1(n_205),
.B2(n_199),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_203),
.A2(n_180),
.B(n_7),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_204),
.C(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_225),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_3),
.B(n_4),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_206),
.C(n_22),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_226),
.C(n_2),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_22),
.C(n_34),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_228),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_231),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_226),
.Y(n_238)
);

AOI31xp33_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_212),
.A3(n_4),
.B(n_5),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_224),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_3),
.B(n_4),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_231),
.B(n_6),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_240),
.B(n_232),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_5),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_233),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_243),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_5),
.A3(n_6),
.B1(n_34),
.B2(n_244),
.C(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_247),
.B(n_6),
.Y(n_248)
);

XNOR2x2_ASAP7_75t_SL g249 ( 
.A(n_248),
.B(n_34),
.Y(n_249)
);


endmodule