module fake_jpeg_23891_n_272 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_46),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_23),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_0),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_50),
.B1(n_22),
.B2(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_36),
.B1(n_24),
.B2(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_17),
.B1(n_23),
.B2(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_71),
.B1(n_24),
.B2(n_19),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_22),
.Y(n_56)
);

FAx1_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_66),
.CI(n_72),
.CON(n_88),
.SN(n_88)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_30),
.B1(n_26),
.B2(n_22),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_63),
.B1(n_67),
.B2(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_69),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_33),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_26),
.B1(n_18),
.B2(n_33),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_19),
.B1(n_13),
.B2(n_21),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_33),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_49),
.C(n_44),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_78),
.Y(n_99)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_70),
.B1(n_65),
.B2(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_90),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_92),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_54),
.B1(n_40),
.B2(n_46),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_110),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_61),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_111),
.C(n_87),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_73),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_112),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_116),
.B1(n_82),
.B2(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_74),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_56),
.C(n_49),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_56),
.B(n_66),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_43),
.B(n_39),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_44),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_44),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_62),
.B1(n_51),
.B2(n_13),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_125),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_85),
.B1(n_81),
.B2(n_84),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_129),
.B1(n_132),
.B2(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_123),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_91),
.C(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_88),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_111),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_100),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_88),
.B1(n_78),
.B2(n_93),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_137),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_77),
.B1(n_62),
.B2(n_76),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_77),
.B1(n_76),
.B2(n_75),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_147),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_143),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_104),
.A3(n_113),
.B1(n_98),
.B2(n_106),
.C1(n_107),
.C2(n_112),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_158),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_112),
.B(n_107),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_159),
.B1(n_131),
.B2(n_119),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_150),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_12),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_122),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_96),
.B1(n_109),
.B2(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_98),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_130),
.B1(n_128),
.B2(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_98),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_116),
.B1(n_100),
.B2(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_104),
.B(n_100),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_124),
.B(n_104),
.Y(n_162)
);

XNOR2x2_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_18),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_170),
.B1(n_174),
.B2(n_176),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_168),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_131),
.B1(n_123),
.B2(n_117),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_120),
.B1(n_77),
.B2(n_64),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_64),
.B1(n_58),
.B2(n_21),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_140),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_184),
.B(n_159),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_153),
.C(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_194),
.C(n_197),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_139),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_153),
.C(n_162),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_150),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_147),
.B1(n_146),
.B2(n_64),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_201),
.B1(n_169),
.B2(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_51),
.C(n_25),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_51),
.C(n_25),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_174),
.C(n_175),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_173),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_25),
.B1(n_16),
.B2(n_14),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_173),
.B1(n_163),
.B2(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_211),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.C(n_220),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_167),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_218),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_193),
.B1(n_188),
.B2(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_178),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_215),
.B(n_216),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_18),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_12),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_0),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_25),
.C(n_16),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_229),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_200),
.B(n_197),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_1),
.B(n_2),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_191),
.B1(n_186),
.B2(n_185),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_213),
.B1(n_208),
.B2(n_12),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_218),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_234),
.C(n_220),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_201),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_242),
.B1(n_245),
.B2(n_3),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_16),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_243),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_16),
.C(n_14),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_241),
.B(n_246),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_1),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_1),
.C(n_3),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_222),
.B1(n_221),
.B2(n_230),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_228),
.B(n_226),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_254),
.B(n_251),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_227),
.B1(n_4),
.B2(n_5),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_6),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_246),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_249),
.B(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_262),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_250),
.B(n_8),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_6),
.B(n_7),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_261),
.A2(n_252),
.B(n_8),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_7),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_266),
.A2(n_260),
.B(n_8),
.Y(n_268)
);

AOI221xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_268),
.B1(n_265),
.B2(n_264),
.C(n_10),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_7),
.B(n_9),
.Y(n_270)
);

AOI221xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_9),
.B1(n_10),
.B2(n_257),
.C(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_9),
.Y(n_272)
);


endmodule