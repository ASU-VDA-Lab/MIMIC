module fake_jpeg_25479_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_22),
.Y(n_32)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_2),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_25),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_19),
.A2(n_13),
.B1(n_18),
.B2(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_31),
.B1(n_20),
.B2(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_18),
.B1(n_14),
.B2(n_9),
.Y(n_31)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_24),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_10),
.B(n_17),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_26),
.B(n_20),
.C(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_26),
.C(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_22),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_41),
.B(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_21),
.B1(n_33),
.B2(n_10),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_26),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_51),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_27),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_44),
.CI(n_42),
.CON(n_55),
.SN(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_65),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_39),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_23),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_59),
.B1(n_21),
.B2(n_52),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_39),
.B1(n_40),
.B2(n_33),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_63),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_55),
.Y(n_67)
);

NOR4xp25_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_17),
.C(n_9),
.D(n_14),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_8),
.C(n_3),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_59),
.B1(n_55),
.B2(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_25),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_86),
.B1(n_73),
.B2(n_71),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_35),
.B1(n_29),
.B2(n_25),
.Y(n_86)
);

AO21x2_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_88),
.B(n_78),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_70),
.B1(n_74),
.B2(n_76),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.C(n_79),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_81),
.B(n_86),
.C(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_97),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_89),
.B1(n_92),
.B2(n_29),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.C(n_23),
.Y(n_100)
);

NOR2xp67_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_85),
.Y(n_96)
);

AOI321xp33_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_81),
.A3(n_23),
.B1(n_29),
.B2(n_25),
.C(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_101),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_0),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_3),
.C(n_4),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_25),
.C(n_3),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_103),
.B(n_4),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_SL g107 ( 
.A1(n_105),
.A2(n_106),
.A3(n_7),
.B1(n_8),
.B2(n_25),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_104),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_8),
.Y(n_108)
);


endmodule