module fake_netlist_1_6954_n_1385 (n_303, n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_304, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_305, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_301, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_302, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1385);
input n_303;
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_304;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_305;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_301;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_302;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1385;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVxp67_ASAP7_75t_SL g306 ( .A(n_29), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_136), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_79), .Y(n_309) );
CKINVDCx14_ASAP7_75t_R g310 ( .A(n_285), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_17), .Y(n_311) );
CKINVDCx16_ASAP7_75t_R g312 ( .A(n_194), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_178), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_11), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_155), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_14), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_181), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_42), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_143), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_6), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_82), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_26), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_179), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_232), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_229), .Y(n_326) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_201), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_174), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_75), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_82), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_119), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_103), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_207), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_278), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_247), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_59), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_26), .Y(n_337) );
CKINVDCx14_ASAP7_75t_R g338 ( .A(n_273), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_123), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_131), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_124), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_164), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_80), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_38), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_46), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_112), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_270), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_72), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_225), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_76), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_296), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_172), .Y(n_352) );
INVxp33_ASAP7_75t_SL g353 ( .A(n_305), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_81), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_196), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_149), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_150), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_25), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_235), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_288), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_35), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_193), .Y(n_362) );
CKINVDCx14_ASAP7_75t_R g363 ( .A(n_254), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_22), .B(n_111), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_190), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_182), .Y(n_366) );
INVxp33_ASAP7_75t_L g367 ( .A(n_269), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_45), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_217), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_197), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_85), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_126), .Y(n_372) );
CKINVDCx14_ASAP7_75t_R g373 ( .A(n_203), .Y(n_373) );
CKINVDCx14_ASAP7_75t_R g374 ( .A(n_161), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_55), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_12), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_233), .Y(n_377) );
INVxp33_ASAP7_75t_L g378 ( .A(n_56), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_28), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_55), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_57), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_299), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_261), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_183), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_47), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_39), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_18), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_222), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_221), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_160), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_304), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_20), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_231), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_95), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_110), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_170), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_199), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_294), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_267), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_206), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_89), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_275), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_100), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_98), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_227), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_171), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_198), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_84), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_147), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_117), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_157), .Y(n_411) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_263), .B(n_209), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_250), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_17), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_104), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_195), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_302), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_152), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_173), .Y(n_419) );
INVxp33_ASAP7_75t_L g420 ( .A(n_29), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_78), .Y(n_421) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_62), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_52), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_137), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_158), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_271), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_7), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_292), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_265), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_100), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_107), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_12), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_118), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_266), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_88), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_276), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_191), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_138), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_87), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_303), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_109), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_219), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_242), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_91), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_259), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_301), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_165), .Y(n_447) );
INVxp33_ASAP7_75t_SL g448 ( .A(n_106), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_56), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_1), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_253), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_83), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_102), .Y(n_453) );
INVxp33_ASAP7_75t_SL g454 ( .A(n_268), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_255), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_142), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_168), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_332), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_332), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_332), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_383), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_317), .Y(n_462) );
INVx4_ASAP7_75t_L g463 ( .A(n_324), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_325), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_325), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_334), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_324), .B(n_0), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_383), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_334), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_317), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_383), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_383), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_339), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_430), .B(n_0), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_403), .B(n_322), .Y(n_475) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_383), .Y(n_476) );
AND2x6_ASAP7_75t_L g477 ( .A(n_342), .B(n_105), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_339), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_331), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_430), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_378), .B(n_1), .Y(n_481) );
AND3x1_ASAP7_75t_L g482 ( .A(n_403), .B(n_2), .C(n_3), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_331), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_341), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_340), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_341), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_420), .B(n_2), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_340), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_360), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_360), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_342), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_463), .B(n_312), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_463), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_480), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_460), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_460), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_460), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_463), .B(n_419), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_488), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_463), .B(n_326), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_474), .B(n_364), .Y(n_502) );
BUFx4f_ASAP7_75t_L g503 ( .A(n_477), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_474), .A2(n_463), .B1(n_487), .B2(n_481), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_488), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_488), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_463), .B(n_391), .Y(n_507) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_467), .A2(n_347), .B(n_346), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_474), .B(n_376), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_467), .B(n_439), .C(n_404), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_460), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_480), .Y(n_512) );
OA22x2_ASAP7_75t_L g513 ( .A1(n_474), .A2(n_323), .B1(n_329), .B2(n_322), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_460), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_477), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_485), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_481), .A2(n_336), .B1(n_386), .B2(n_368), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_464), .B(n_437), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_481), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_488), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_485), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_481), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_464), .B(n_437), .Y(n_525) );
INVx4_ASAP7_75t_L g526 ( .A(n_477), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_471), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_487), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_471), .Y(n_529) );
BUFx3_ASAP7_75t_L g530 ( .A(n_492), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_487), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_471), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_464), .B(n_307), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_487), .B(n_376), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_467), .B(n_336), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_465), .B(n_328), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_485), .Y(n_537) );
AO22x2_ASAP7_75t_L g538 ( .A1(n_465), .A2(n_364), .B1(n_347), .B2(n_351), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_494), .B(n_465), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_531), .B(n_475), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_503), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_495), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_495), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_512), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_517), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_494), .Y(n_546) );
INVx4_ASAP7_75t_L g547 ( .A(n_515), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_520), .B(n_466), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_517), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_521), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_521), .Y(n_551) );
INVxp33_ASAP7_75t_L g552 ( .A(n_535), .Y(n_552) );
CKINVDCx11_ASAP7_75t_R g553 ( .A(n_528), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_538), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_502), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_523), .Y(n_556) );
BUFx8_ASAP7_75t_L g557 ( .A(n_535), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_509), .B(n_482), .Y(n_558) );
INVx5_ASAP7_75t_L g559 ( .A(n_515), .Y(n_559) );
OR2x6_ASAP7_75t_L g560 ( .A(n_502), .B(n_475), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_523), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_537), .Y(n_562) );
BUFx3_ASAP7_75t_L g563 ( .A(n_530), .Y(n_563) );
BUFx3_ASAP7_75t_L g564 ( .A(n_530), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_520), .B(n_466), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_510), .A2(n_482), .B1(n_386), .B2(n_401), .Y(n_567) );
AND2x6_ASAP7_75t_L g568 ( .A(n_509), .B(n_466), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_537), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_496), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_504), .B(n_328), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_497), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_497), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_498), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_524), .B(n_475), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_498), .Y(n_577) );
BUFx12f_ASAP7_75t_L g578 ( .A(n_502), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_513), .A2(n_473), .B1(n_478), .B2(n_469), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_509), .B(n_469), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_511), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_514), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_509), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_534), .B(n_469), .Y(n_585) );
BUFx3_ASAP7_75t_L g586 ( .A(n_530), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_514), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_516), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_518), .A2(n_482), .B1(n_401), .B2(n_414), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_534), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_500), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_538), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_519), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_519), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_525), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_493), .B(n_473), .Y(n_599) );
BUFx4f_ASAP7_75t_L g600 ( .A(n_503), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_525), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_499), .B(n_473), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_499), .B(n_536), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_538), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_501), .B(n_478), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_500), .Y(n_606) );
AND3x1_ASAP7_75t_SL g607 ( .A(n_518), .B(n_311), .C(n_309), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_507), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_538), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_508), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_508), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_515), .B(n_333), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_508), .B(n_478), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_500), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_508), .Y(n_615) );
OR2x6_ASAP7_75t_L g616 ( .A(n_513), .B(n_323), .Y(n_616) );
NAND3xp33_ASAP7_75t_SL g617 ( .A(n_533), .B(n_440), .C(n_411), .Y(n_617) );
INVx4_ASAP7_75t_L g618 ( .A(n_515), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_505), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_533), .A2(n_486), .B(n_484), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_513), .B(n_484), .Y(n_621) );
BUFx4f_ASAP7_75t_L g622 ( .A(n_526), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_526), .B(n_484), .Y(n_623) );
BUFx4f_ASAP7_75t_L g624 ( .A(n_526), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_526), .B(n_367), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_505), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_596), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_596), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_555), .B(n_458), .Y(n_629) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_595), .B(n_354), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_597), .B(n_486), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_545), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_604), .A2(n_486), .B1(n_477), .B2(n_459), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_545), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_560), .A2(n_414), .B1(n_421), .B2(n_368), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_549), .Y(n_636) );
AND2x2_ASAP7_75t_SL g637 ( .A(n_595), .B(n_458), .Y(n_637) );
BUFx5_ASAP7_75t_L g638 ( .A(n_568), .Y(n_638) );
BUFx3_ASAP7_75t_L g639 ( .A(n_578), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_552), .B(n_421), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_604), .A2(n_477), .B1(n_459), .B2(n_458), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_578), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_597), .B(n_459), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_568), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_598), .Y(n_645) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_568), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_560), .A2(n_315), .B1(n_448), .B2(n_353), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_598), .B(n_492), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_568), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_601), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_560), .B(n_306), .Y(n_651) );
INVx3_ASAP7_75t_L g652 ( .A(n_549), .Y(n_652) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_568), .Y(n_653) );
BUFx4_ASAP7_75t_SL g654 ( .A(n_560), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_551), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_601), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_551), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_561), .Y(n_658) );
OR2x2_ASAP7_75t_SL g659 ( .A(n_617), .B(n_329), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_567), .B(n_335), .C(n_333), .Y(n_660) );
OR2x6_ASAP7_75t_L g661 ( .A(n_555), .B(n_337), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_609), .A2(n_477), .B1(n_470), .B2(n_462), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_620), .A2(n_485), .B(n_483), .C(n_479), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_554), .A2(n_609), .B1(n_593), .B2(n_579), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_554), .A2(n_477), .B1(n_470), .B2(n_462), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_590), .B(n_343), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_548), .A2(n_483), .B1(n_491), .B2(n_479), .Y(n_667) );
BUFx12f_ASAP7_75t_L g668 ( .A(n_553), .Y(n_668) );
BUFx3_ASAP7_75t_L g669 ( .A(n_557), .Y(n_669) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_616), .B(n_314), .Y(n_670) );
AND2x4_ASAP7_75t_SL g671 ( .A(n_542), .B(n_337), .Y(n_671) );
INVx8_ASAP7_75t_L g672 ( .A(n_568), .Y(n_672) );
INVx4_ASAP7_75t_L g673 ( .A(n_561), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_546), .B(n_335), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_543), .B(n_380), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_SL g676 ( .A1(n_625), .A2(n_310), .B(n_363), .C(n_338), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_613), .B(n_492), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_576), .A2(n_353), .B1(n_448), .B2(n_315), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_613), .B(n_492), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_540), .A2(n_454), .B1(n_422), .B2(n_372), .Y(n_680) );
INVx2_ASAP7_75t_SL g681 ( .A(n_557), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_608), .B(n_454), .Y(n_682) );
INVx3_ASAP7_75t_L g683 ( .A(n_569), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_569), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_584), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_599), .B(n_316), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_557), .Y(n_687) );
OR2x6_ASAP7_75t_L g688 ( .A(n_544), .B(n_345), .Y(n_688) );
OAI21x1_ASAP7_75t_SL g689 ( .A1(n_621), .A2(n_351), .B(n_346), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_607), .Y(n_690) );
BUFx3_ASAP7_75t_L g691 ( .A(n_550), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_613), .B(n_492), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g693 ( .A(n_608), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_610), .B(n_462), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_546), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_550), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_558), .A2(n_372), .B1(n_377), .B2(n_349), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_558), .A2(n_377), .B1(n_384), .B2(n_349), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_610), .B(n_462), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_585), .B(n_345), .Y(n_700) );
INVx4_ASAP7_75t_L g701 ( .A(n_563), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_623), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_556), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_589), .B(n_348), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_556), .Y(n_705) );
CKINVDCx8_ASAP7_75t_R g706 ( .A(n_558), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_572), .B(n_318), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_599), .B(n_321), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_562), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_581), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_616), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_570), .Y(n_712) );
AND2x6_ASAP7_75t_L g713 ( .A(n_611), .B(n_615), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_570), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_611), .A2(n_483), .B(n_491), .C(n_479), .Y(n_715) );
INVx3_ASAP7_75t_L g716 ( .A(n_563), .Y(n_716) );
INVx3_ASAP7_75t_L g717 ( .A(n_564), .Y(n_717) );
O2A1O1Ixp33_ASAP7_75t_L g718 ( .A1(n_565), .A2(n_348), .B(n_358), .C(n_350), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_599), .B(n_330), .Y(n_719) );
INVx5_ASAP7_75t_L g720 ( .A(n_616), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_571), .Y(n_721) );
OR2x6_ASAP7_75t_L g722 ( .A(n_616), .B(n_350), .Y(n_722) );
BUFx4f_ASAP7_75t_L g723 ( .A(n_615), .Y(n_723) );
INVx4_ASAP7_75t_L g724 ( .A(n_564), .Y(n_724) );
INVx5_ASAP7_75t_L g725 ( .A(n_541), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_605), .B(n_371), .Y(n_726) );
INVx2_ASAP7_75t_SL g727 ( .A(n_602), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_539), .A2(n_375), .B1(n_387), .B2(n_385), .C(n_379), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_603), .A2(n_358), .B1(n_444), .B2(n_361), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_577), .Y(n_730) );
BUFx2_ASAP7_75t_SL g731 ( .A(n_623), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_571), .A2(n_483), .B1(n_491), .B2(n_479), .Y(n_732) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_586), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_623), .A2(n_477), .B1(n_470), .B2(n_462), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_574), .A2(n_477), .B1(n_470), .B2(n_462), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_577), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_574), .Y(n_737) );
BUFx12f_ASAP7_75t_L g738 ( .A(n_541), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_575), .B(n_470), .Y(n_739) );
BUFx12f_ASAP7_75t_L g740 ( .A(n_541), .Y(n_740) );
BUFx12f_ASAP7_75t_L g741 ( .A(n_541), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_586), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g743 ( .A(n_575), .Y(n_743) );
OR2x2_ASAP7_75t_SL g744 ( .A(n_582), .B(n_361), .Y(n_744) );
BUFx2_ASAP7_75t_L g745 ( .A(n_582), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_580), .A2(n_477), .B1(n_489), .B2(n_470), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_580), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g748 ( .A1(n_626), .A2(n_327), .B(n_320), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_583), .Y(n_749) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_583), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_612), .B(n_393), .C(n_384), .Y(n_751) );
BUFx4_ASAP7_75t_SL g752 ( .A(n_587), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_631), .A2(n_624), .B(n_622), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_718), .A2(n_587), .B(n_591), .C(n_573), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_723), .A2(n_626), .B1(n_588), .B2(n_374), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_723), .A2(n_588), .B1(n_373), .B2(n_600), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_631), .A2(n_600), .B1(n_395), .B2(n_402), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_643), .A2(n_624), .B(n_622), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_677), .A2(n_622), .B(n_624), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g760 ( .A1(n_627), .A2(n_491), .B(n_489), .C(n_600), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_743), .A2(n_393), .B1(n_402), .B2(n_395), .Y(n_761) );
BUFx2_ASAP7_75t_L g762 ( .A(n_639), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_720), .B(n_559), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_727), .B(n_547), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_642), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_682), .B(n_547), .Y(n_766) );
NAND2x1p5_ASAP7_75t_L g767 ( .A(n_720), .B(n_547), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_654), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_628), .B(n_392), .Y(n_769) );
INVx3_ASAP7_75t_SL g770 ( .A(n_687), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_711), .A2(n_405), .B1(n_455), .B2(n_413), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_673), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_668), .Y(n_773) );
INVx8_ASAP7_75t_L g774 ( .A(n_672), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_645), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_650), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_661), .A2(n_450), .B1(n_452), .B2(n_449), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_673), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_656), .Y(n_779) );
INVxp67_ASAP7_75t_L g780 ( .A(n_731), .Y(n_780) );
AOI221xp5_ASAP7_75t_L g781 ( .A1(n_728), .A2(n_394), .B1(n_423), .B2(n_415), .C(n_408), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_682), .B(n_618), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_722), .A2(n_413), .B1(n_455), .B2(n_405), .Y(n_783) );
INVx3_ASAP7_75t_L g784 ( .A(n_738), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_752), .Y(n_785) );
INVxp67_ASAP7_75t_L g786 ( .A(n_695), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_722), .A2(n_566), .B1(n_594), .B2(n_541), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_661), .B(n_449), .Y(n_788) );
AND2x4_ASAP7_75t_L g789 ( .A(n_722), .B(n_618), .Y(n_789) );
INVx6_ASAP7_75t_SL g790 ( .A(n_688), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_750), .A2(n_594), .B1(n_566), .B2(n_416), .Y(n_791) );
INVx1_ASAP7_75t_SL g792 ( .A(n_752), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_720), .B(n_618), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_704), .A2(n_477), .B1(n_489), .B2(n_432), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_643), .Y(n_795) );
INVx4_ASAP7_75t_L g796 ( .A(n_672), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g797 ( .A1(n_630), .A2(n_452), .B1(n_453), .B2(n_450), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_744), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_637), .A2(n_477), .B1(n_489), .B2(n_435), .Y(n_799) );
INVx2_ASAP7_75t_SL g800 ( .A(n_654), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_718), .A2(n_489), .B(n_355), .C(n_356), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_691), .Y(n_802) );
INVx2_ASAP7_75t_SL g803 ( .A(n_669), .Y(n_803) );
INVx1_ASAP7_75t_SL g804 ( .A(n_671), .Y(n_804) );
INVx3_ASAP7_75t_L g805 ( .A(n_740), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_685), .Y(n_806) );
OAI221xp5_ASAP7_75t_L g807 ( .A1(n_688), .A2(n_427), .B1(n_453), .B2(n_381), .C(n_344), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_750), .A2(n_702), .B1(n_720), .B2(n_745), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_696), .Y(n_809) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_629), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_688), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_702), .A2(n_566), .B1(n_594), .B2(n_406), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_644), .A2(n_566), .B1(n_594), .B2(n_489), .Y(n_813) );
INVx2_ASAP7_75t_SL g814 ( .A(n_681), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_700), .Y(n_815) );
OAI22xp33_ASAP7_75t_L g816 ( .A1(n_706), .A2(n_381), .B1(n_344), .B2(n_355), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_635), .A2(n_566), .B1(n_594), .B2(n_477), .Y(n_817) );
A2O1A1Ixp33_ASAP7_75t_L g818 ( .A1(n_707), .A2(n_356), .B(n_357), .C(n_352), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_686), .A2(n_490), .B1(n_488), .B2(n_357), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_703), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_629), .Y(n_821) );
AOI21xp33_ASAP7_75t_L g822 ( .A1(n_660), .A2(n_559), .B(n_382), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_644), .A2(n_359), .B1(n_362), .B2(n_352), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_686), .A2(n_490), .B1(n_488), .B2(n_362), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_690), .A2(n_365), .B1(n_446), .B2(n_434), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_708), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_651), .A2(n_313), .B1(n_319), .B2(n_308), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_651), .A2(n_366), .B1(n_441), .B2(n_359), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_705), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_675), .A2(n_366), .B1(n_442), .B2(n_441), .Y(n_830) );
INVxp67_ASAP7_75t_L g831 ( .A(n_713), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_675), .A2(n_443), .B1(n_445), .B2(n_442), .Y(n_832) );
AOI222xp33_ASAP7_75t_L g833 ( .A1(n_728), .A2(n_457), .B1(n_443), .B2(n_445), .C1(n_447), .C2(n_451), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_708), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_649), .A2(n_451), .B1(n_457), .B2(n_447), .Y(n_835) );
O2A1O1Ixp33_ASAP7_75t_L g836 ( .A1(n_748), .A2(n_707), .B(n_664), .C(n_726), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_719), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_649), .A2(n_369), .B1(n_388), .B2(n_370), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_646), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_709), .Y(n_840) );
AO31x2_ASAP7_75t_L g841 ( .A1(n_715), .A2(n_472), .A3(n_468), .B(n_461), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_719), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_739), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_640), .A2(n_389), .B1(n_396), .B2(n_390), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_693), .A2(n_397), .B1(n_399), .B2(n_398), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g846 ( .A1(n_678), .A2(n_438), .B1(n_400), .B2(n_407), .C(n_409), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_664), .A2(n_490), .B1(n_488), .B2(n_410), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_739), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_710), .B(n_559), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_721), .A2(n_490), .B1(n_488), .B2(n_417), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_694), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_677), .A2(n_606), .B(n_592), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_684), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_672), .A2(n_418), .B1(n_425), .B2(n_424), .Y(n_854) );
AOI21xp33_ASAP7_75t_L g855 ( .A1(n_676), .A2(n_559), .B(n_428), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_697), .Y(n_856) );
NOR2xp33_ASAP7_75t_SL g857 ( .A(n_646), .B(n_559), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_666), .A2(n_426), .B1(n_431), .B2(n_429), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_666), .A2(n_433), .B1(n_456), .B2(n_436), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_748), .A2(n_434), .B1(n_446), .B2(n_365), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_713), .A2(n_488), .B1(n_490), .B2(n_472), .Y(n_861) );
BUFx2_ASAP7_75t_L g862 ( .A(n_713), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g863 ( .A1(n_726), .A2(n_488), .B1(n_490), .B2(n_606), .C(n_592), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_694), .Y(n_864) );
O2A1O1Ixp33_ASAP7_75t_L g865 ( .A1(n_689), .A2(n_505), .B(n_522), .C(n_506), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_699), .Y(n_866) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_713), .A2(n_490), .B1(n_472), .B2(n_5), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_670), .A2(n_490), .B1(n_619), .B2(n_614), .Y(n_868) );
BUFx3_ASAP7_75t_L g869 ( .A(n_741), .Y(n_869) );
CKINVDCx8_ASAP7_75t_R g870 ( .A(n_646), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_713), .A2(n_490), .B1(n_619), .B2(n_614), .Y(n_871) );
AND2x4_ASAP7_75t_L g872 ( .A(n_653), .B(n_412), .Y(n_872) );
CKINVDCx6p67_ASAP7_75t_R g873 ( .A(n_653), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_638), .A2(n_490), .B1(n_472), .B2(n_5), .Y(n_874) );
INVx3_ASAP7_75t_L g875 ( .A(n_653), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_737), .A2(n_472), .B1(n_468), .B2(n_461), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_638), .A2(n_6), .B1(n_3), .B2(n_4), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_684), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_679), .A2(n_468), .B1(n_461), .B2(n_506), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_729), .B(n_4), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_679), .A2(n_468), .B1(n_461), .B2(n_506), .Y(n_881) );
O2A1O1Ixp33_ASAP7_75t_L g882 ( .A1(n_667), .A2(n_522), .B(n_9), .C(n_7), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_684), .Y(n_883) );
AND2x4_ASAP7_75t_L g884 ( .A(n_747), .B(n_8), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_701), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_647), .A2(n_522), .B1(n_476), .B2(n_471), .Y(n_886) );
AOI22xp33_ASAP7_75t_SL g887 ( .A1(n_638), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_729), .A2(n_476), .B1(n_471), .B2(n_527), .Y(n_888) );
INVx2_ASAP7_75t_L g889 ( .A(n_636), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_692), .A2(n_476), .B1(n_471), .B2(n_13), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_788), .B(n_680), .Y(n_891) );
AOI222xp33_ASAP7_75t_L g892 ( .A1(n_815), .A2(n_674), .B1(n_699), .B2(n_667), .C1(n_732), .C2(n_734), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_795), .A2(n_692), .B1(n_749), .B2(n_730), .Y(n_893) );
OAI221xp5_ASAP7_75t_SL g894 ( .A1(n_797), .A2(n_698), .B1(n_734), .B2(n_662), .C(n_735), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_777), .A2(n_652), .B1(n_683), .B2(n_636), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_809), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_820), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_797), .B(n_632), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_836), .A2(n_665), .B(n_662), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_811), .A2(n_638), .B1(n_683), .B2(n_652), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_829), .Y(n_901) );
AOI221xp5_ASAP7_75t_L g902 ( .A1(n_781), .A2(n_732), .B1(n_663), .B2(n_648), .C(n_735), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_798), .A2(n_714), .B1(n_736), .B2(n_712), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_806), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_810), .B(n_634), .Y(n_905) );
CKINVDCx11_ASAP7_75t_R g906 ( .A(n_770), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_880), .A2(n_655), .B1(n_658), .B2(n_657), .Y(n_907) );
A2O1A1Ixp33_ASAP7_75t_L g908 ( .A1(n_754), .A2(n_648), .B(n_746), .C(n_633), .Y(n_908) );
AOI22xp33_ASAP7_75t_SL g909 ( .A1(n_768), .A2(n_638), .B1(n_659), .B2(n_701), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_777), .A2(n_665), .B1(n_633), .B2(n_641), .Y(n_910) );
BUFx12f_ASAP7_75t_L g911 ( .A(n_773), .Y(n_911) );
AOI31xp33_ASAP7_75t_L g912 ( .A1(n_792), .A2(n_746), .A3(n_641), .B(n_751), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_884), .A2(n_638), .B1(n_724), .B2(n_717), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_810), .B(n_724), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_884), .A2(n_717), .B1(n_742), .B2(n_716), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_821), .B(n_716), .Y(n_916) );
BUFx3_ASAP7_75t_L g917 ( .A(n_869), .Y(n_917) );
BUFx12f_ASAP7_75t_L g918 ( .A(n_785), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_807), .A2(n_742), .B1(n_733), .B2(n_725), .Y(n_919) );
AND2x4_ASAP7_75t_L g920 ( .A(n_789), .B(n_725), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_851), .A2(n_733), .B1(n_725), .B2(n_476), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_846), .A2(n_733), .B1(n_725), .B2(n_476), .C(n_471), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_790), .A2(n_476), .B1(n_471), .B2(n_13), .Y(n_923) );
BUFx3_ASAP7_75t_L g924 ( .A(n_762), .Y(n_924) );
AOI22xp33_ASAP7_75t_SL g925 ( .A1(n_768), .A2(n_476), .B1(n_471), .B2(n_15), .Y(n_925) );
A2O1A1Ixp33_ASAP7_75t_L g926 ( .A1(n_882), .A2(n_476), .B(n_471), .C(n_527), .Y(n_926) );
OAI21x1_ASAP7_75t_L g927 ( .A1(n_865), .A2(n_476), .B(n_527), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_786), .B(n_11), .Y(n_928) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_790), .A2(n_476), .B1(n_15), .B2(n_16), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_804), .A2(n_532), .B1(n_529), .B2(n_527), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_864), .A2(n_532), .B1(n_529), .B2(n_527), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_786), .B(n_14), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_775), .B(n_16), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_776), .Y(n_934) );
INVx3_ASAP7_75t_L g935 ( .A(n_870), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_866), .A2(n_532), .B1(n_529), .B2(n_527), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_799), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_843), .A2(n_532), .B1(n_529), .B2(n_22), .Y(n_938) );
INVx2_ASAP7_75t_SL g939 ( .A(n_784), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_856), .A2(n_532), .B1(n_529), .B2(n_23), .Y(n_940) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_808), .Y(n_941) );
OAI221xp5_ASAP7_75t_L g942 ( .A1(n_844), .A2(n_532), .B1(n_529), .B2(n_23), .C(n_24), .Y(n_942) );
AOI31xp33_ASAP7_75t_L g943 ( .A1(n_800), .A2(n_19), .A3(n_21), .B(n_24), .Y(n_943) );
AOI222xp33_ASAP7_75t_L g944 ( .A1(n_826), .A2(n_21), .B1(n_25), .B2(n_27), .C1(n_28), .C2(n_30), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_848), .A2(n_27), .B1(n_30), .B2(n_31), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_771), .B(n_31), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_799), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_947) );
INVx2_ASAP7_75t_SL g948 ( .A(n_784), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_779), .Y(n_949) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_845), .A2(n_32), .B1(n_33), .B2(n_34), .C(n_35), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g951 ( .A1(n_783), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_840), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_761), .B(n_36), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g954 ( .A(n_874), .B(n_37), .C(n_39), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_765), .Y(n_955) );
AOI22xp5_ASAP7_75t_L g956 ( .A1(n_766), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_956) );
BUFx3_ASAP7_75t_L g957 ( .A(n_805), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_841), .Y(n_958) );
AO21x2_ASAP7_75t_L g959 ( .A1(n_760), .A2(n_113), .B(n_108), .Y(n_959) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_782), .A2(n_40), .B1(n_41), .B2(n_43), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_780), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_961) );
OAI221xp5_ASAP7_75t_L g962 ( .A1(n_830), .A2(n_44), .B1(n_46), .B2(n_47), .C(n_48), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_833), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_816), .A2(n_49), .B1(n_50), .B2(n_51), .C(n_52), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_834), .B(n_51), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_837), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_842), .A2(n_816), .B1(n_825), .B2(n_858), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_878), .Y(n_968) );
OAI21x1_ASAP7_75t_L g969 ( .A1(n_852), .A2(n_115), .B(n_114), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_859), .B(n_53), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_841), .Y(n_971) );
AOI222xp33_ASAP7_75t_L g972 ( .A1(n_832), .A2(n_53), .B1(n_54), .B2(n_57), .C1(n_58), .C2(n_59), .Y(n_972) );
AND2x6_ASAP7_75t_L g973 ( .A(n_789), .B(n_116), .Y(n_973) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_878), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_841), .Y(n_975) );
INVx5_ASAP7_75t_L g976 ( .A(n_774), .Y(n_976) );
OAI33xp33_ASAP7_75t_L g977 ( .A1(n_854), .A2(n_54), .A3(n_58), .B1(n_60), .B2(n_61), .B3(n_62), .Y(n_977) );
BUFx6f_ASAP7_75t_L g978 ( .A(n_767), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_805), .B(n_60), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_818), .A2(n_61), .B1(n_63), .B2(n_64), .C(n_65), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_825), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_981) );
AOI33xp33_ASAP7_75t_L g982 ( .A1(n_828), .A2(n_66), .A3(n_67), .B1(n_68), .B2(n_69), .B3(n_70), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_780), .B(n_66), .Y(n_983) );
OAI322xp33_ASAP7_75t_L g984 ( .A1(n_827), .A2(n_67), .A3(n_68), .B1(n_69), .B2(n_70), .C1(n_71), .C2(n_72), .Y(n_984) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_767), .Y(n_985) );
XNOR2xp5_ASAP7_75t_L g986 ( .A(n_803), .B(n_71), .Y(n_986) );
NOR2xp67_ASAP7_75t_SL g987 ( .A(n_796), .B(n_73), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_847), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_769), .B(n_74), .Y(n_989) );
OAI22x1_ASAP7_75t_L g990 ( .A1(n_770), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_802), .B(n_77), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_801), .A2(n_79), .B1(n_80), .B2(n_81), .C(n_83), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_841), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_867), .A2(n_84), .B1(n_85), .B2(n_86), .Y(n_994) );
AOI22xp33_ASAP7_75t_SL g995 ( .A1(n_755), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_814), .B(n_89), .Y(n_996) );
OA21x2_ASAP7_75t_L g997 ( .A1(n_847), .A2(n_300), .B(n_202), .Y(n_997) );
OA21x2_ASAP7_75t_L g998 ( .A1(n_863), .A2(n_298), .B(n_200), .Y(n_998) );
CKINVDCx5p33_ASAP7_75t_R g999 ( .A(n_774), .Y(n_999) );
OAI21xp33_ASAP7_75t_L g1000 ( .A1(n_794), .A2(n_90), .B(n_91), .Y(n_1000) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_890), .A2(n_90), .B1(n_92), .B2(n_93), .C(n_94), .Y(n_1001) );
AOI21xp5_ASAP7_75t_SL g1002 ( .A1(n_831), .A2(n_204), .B(n_295), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_867), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_1003) );
OAI221xp5_ASAP7_75t_L g1004 ( .A1(n_794), .A2(n_95), .B1(n_96), .B2(n_97), .C(n_98), .Y(n_1004) );
AO31x2_ASAP7_75t_L g1005 ( .A1(n_787), .A2(n_96), .A3(n_97), .B(n_99), .Y(n_1005) );
OAI22xp5_ASAP7_75t_SL g1006 ( .A1(n_877), .A2(n_99), .B1(n_101), .B2(n_102), .Y(n_1006) );
O2A1O1Ixp33_ASAP7_75t_L g1007 ( .A1(n_838), .A2(n_101), .B(n_103), .C(n_104), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_772), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_764), .B(n_120), .Y(n_1009) );
OAI21x1_ASAP7_75t_L g1010 ( .A1(n_871), .A2(n_121), .B(n_122), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_877), .A2(n_125), .B1(n_127), .B2(n_128), .Y(n_1011) );
NOR2xp33_ASAP7_75t_R g1012 ( .A(n_774), .B(n_297), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1013 ( .A(n_793), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_778), .Y(n_1014) );
OAI21xp33_ASAP7_75t_SL g1015 ( .A1(n_831), .A2(n_129), .B(n_130), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1016 ( .A(n_796), .B(n_132), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_889), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_887), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_968), .Y(n_1019) );
INVx1_ASAP7_75t_SL g1020 ( .A(n_917), .Y(n_1020) );
INVx1_ASAP7_75t_SL g1021 ( .A(n_917), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_967), .A2(n_887), .B1(n_874), .B2(n_872), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_904), .Y(n_1023) );
INVx3_ASAP7_75t_L g1024 ( .A(n_978), .Y(n_1024) );
AOI21xp5_ASAP7_75t_L g1025 ( .A1(n_893), .A2(n_862), .B(n_753), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_891), .B(n_764), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_967), .A2(n_861), .B1(n_888), .B2(n_756), .Y(n_1027) );
NAND3xp33_ASAP7_75t_L g1028 ( .A(n_982), .B(n_860), .C(n_872), .Y(n_1028) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_963), .A2(n_886), .B1(n_817), .B2(n_819), .C(n_824), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g1030 ( .A(n_968), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_974), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_924), .B(n_885), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_958), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_958), .Y(n_1034) );
AOI221xp5_ASAP7_75t_L g1035 ( .A1(n_984), .A2(n_835), .B1(n_823), .B2(n_822), .C(n_824), .Y(n_1035) );
BUFx6f_ASAP7_75t_L g1036 ( .A(n_978), .Y(n_1036) );
INVx2_ASAP7_75t_L g1037 ( .A(n_975), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_924), .B(n_885), .Y(n_1038) );
CKINVDCx8_ASAP7_75t_R g1039 ( .A(n_955), .Y(n_1039) );
OAI211xp5_ASAP7_75t_L g1040 ( .A1(n_944), .A2(n_819), .B(n_855), .C(n_861), .Y(n_1040) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_963), .A2(n_757), .B1(n_881), .B2(n_879), .C(n_850), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_898), .A2(n_791), .B1(n_849), .B2(n_812), .Y(n_1042) );
AOI222xp33_ASAP7_75t_L g1043 ( .A1(n_1006), .A2(n_850), .B1(n_793), .B2(n_759), .C1(n_763), .C2(n_876), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_905), .B(n_839), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_934), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1046 ( .A(n_1012), .Y(n_1046) );
NAND4xp25_ASAP7_75t_L g1047 ( .A(n_981), .B(n_876), .C(n_868), .D(n_758), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_943), .A2(n_857), .B1(n_873), .B2(n_875), .Y(n_1048) );
AOI22xp33_ASAP7_75t_SL g1049 ( .A1(n_1012), .A2(n_875), .B1(n_883), .B2(n_853), .Y(n_1049) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_973), .A2(n_813), .B1(n_140), .B2(n_141), .Y(n_1050) );
OA21x2_ASAP7_75t_L g1051 ( .A1(n_975), .A2(n_139), .B(n_144), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_949), .Y(n_1052) );
INVx2_ASAP7_75t_L g1053 ( .A(n_993), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_952), .B(n_145), .Y(n_1054) );
INVxp67_ASAP7_75t_SL g1055 ( .A(n_978), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_974), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_928), .B(n_146), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_993), .Y(n_1058) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_973), .A2(n_946), .B1(n_954), .B2(n_1013), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_978), .Y(n_1060) );
INVx4_ASAP7_75t_L g1061 ( .A(n_976), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_914), .B(n_148), .Y(n_1062) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_932), .B(n_293), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g1064 ( .A1(n_973), .A2(n_151), .B1(n_153), .B2(n_154), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_966), .Y(n_1065) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_985), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_896), .B(n_291), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_977), .A2(n_156), .B1(n_159), .B2(n_162), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_979), .B(n_163), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_897), .Y(n_1070) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_973), .A2(n_166), .B1(n_167), .B2(n_169), .Y(n_1071) );
OAI321xp33_ASAP7_75t_L g1072 ( .A1(n_929), .A2(n_175), .A3(n_176), .B1(n_177), .B2(n_180), .C(n_184), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_971), .Y(n_1073) );
AOI21xp5_ASAP7_75t_L g1074 ( .A1(n_895), .A2(n_185), .B(n_186), .Y(n_1074) );
OAI21xp33_ASAP7_75t_L g1075 ( .A1(n_982), .A2(n_187), .B(n_188), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_985), .B(n_189), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_915), .A2(n_192), .B1(n_205), .B2(n_208), .Y(n_1077) );
NAND2xp5_ASAP7_75t_SL g1078 ( .A(n_929), .B(n_210), .Y(n_1078) );
OAI22xp5_ASAP7_75t_SL g1079 ( .A1(n_986), .A2(n_211), .B1(n_212), .B2(n_213), .Y(n_1079) );
AOI211xp5_ASAP7_75t_L g1080 ( .A1(n_950), .A2(n_214), .B(n_215), .C(n_216), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_996), .B(n_218), .Y(n_1081) );
NAND4xp25_ASAP7_75t_L g1082 ( .A(n_981), .B(n_220), .C(n_223), .D(n_224), .Y(n_1082) );
OAI22xp5_ASAP7_75t_SL g1083 ( .A1(n_990), .A2(n_226), .B1(n_228), .B2(n_230), .Y(n_1083) );
OAI31xp33_ASAP7_75t_SL g1084 ( .A1(n_961), .A2(n_234), .A3(n_236), .B(n_237), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_989), .B(n_290), .Y(n_1085) );
NOR2x1_ASAP7_75t_L g1086 ( .A(n_957), .B(n_238), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_915), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_1087) );
OAI321xp33_ASAP7_75t_L g1088 ( .A1(n_994), .A2(n_243), .A3(n_244), .B1(n_245), .B2(n_246), .C(n_248), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_901), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1017), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1017), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_913), .A2(n_249), .B1(n_251), .B2(n_256), .Y(n_1092) );
OAI22xp5_ASAP7_75t_SL g1093 ( .A1(n_999), .A2(n_257), .B1(n_258), .B2(n_260), .Y(n_1093) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_910), .A2(n_262), .B1(n_264), .B2(n_272), .Y(n_1094) );
AO21x2_ASAP7_75t_L g1095 ( .A1(n_926), .A2(n_274), .B(n_277), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_957), .B(n_279), .Y(n_1096) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_976), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_991), .Y(n_1098) );
OAI33xp33_ASAP7_75t_L g1099 ( .A1(n_937), .A2(n_280), .A3(n_281), .B1(n_283), .B2(n_284), .B3(n_286), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_933), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_953), .B(n_287), .Y(n_1101) );
NAND3xp33_ASAP7_75t_L g1102 ( .A(n_972), .B(n_289), .C(n_964), .Y(n_1102) );
INVx1_ASAP7_75t_SL g1103 ( .A(n_906), .Y(n_1103) );
AND2x2_ASAP7_75t_SL g1104 ( .A(n_997), .B(n_1016), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_965), .B(n_920), .Y(n_1105) );
AOI22xp33_ASAP7_75t_SL g1106 ( .A1(n_973), .A2(n_997), .B1(n_985), .B2(n_1016), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_920), .B(n_939), .Y(n_1107) );
BUFx8_ASAP7_75t_SL g1108 ( .A(n_911), .Y(n_1108) );
AND2x4_ASAP7_75t_L g1109 ( .A(n_976), .B(n_1009), .Y(n_1109) );
OAI21x1_ASAP7_75t_L g1110 ( .A1(n_927), .A2(n_969), .B(n_1010), .Y(n_1110) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_997), .A2(n_998), .B1(n_976), .B2(n_1004), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_918), .Y(n_1112) );
OAI322xp33_ASAP7_75t_L g1113 ( .A1(n_956), .A2(n_960), .A3(n_951), .B1(n_962), .B2(n_970), .C1(n_983), .C2(n_992), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_892), .A2(n_1001), .B1(n_1000), .B2(n_995), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1115 ( .A1(n_940), .A2(n_942), .B1(n_988), .B2(n_947), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_980), .A2(n_994), .B1(n_1003), .B2(n_899), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1008), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1014), .Y(n_1118) );
OR2x2_ASAP7_75t_L g1119 ( .A(n_948), .B(n_916), .Y(n_1119) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_941), .A2(n_998), .B1(n_923), .B2(n_912), .Y(n_1120) );
AO21x2_ASAP7_75t_L g1121 ( .A1(n_926), .A2(n_941), .B(n_908), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1033), .Y(n_1122) );
BUFx3_ASAP7_75t_L g1123 ( .A(n_1097), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1090), .B(n_1005), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1033), .Y(n_1125) );
AOI222xp33_ASAP7_75t_SL g1126 ( .A1(n_1103), .A2(n_894), .B1(n_935), .B2(n_1005), .C1(n_987), .C2(n_945), .Y(n_1126) );
NAND3xp33_ASAP7_75t_L g1127 ( .A(n_1059), .B(n_945), .C(n_1003), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1023), .B(n_1005), .Y(n_1128) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1034), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_1043), .A2(n_909), .B1(n_925), .B2(n_919), .Y(n_1130) );
OAI211xp5_ASAP7_75t_SL g1131 ( .A1(n_1020), .A2(n_1007), .B(n_919), .C(n_913), .Y(n_1131) );
OAI33xp33_ASAP7_75t_L g1132 ( .A1(n_1048), .A2(n_1005), .A3(n_903), .B1(n_938), .B2(n_1018), .B3(n_1011), .Y(n_1132) );
NAND3xp33_ASAP7_75t_L g1133 ( .A(n_1114), .B(n_1018), .C(n_1011), .Y(n_1133) );
AOI21xp5_ASAP7_75t_L g1134 ( .A1(n_1104), .A2(n_998), .B(n_931), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1034), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1045), .B(n_903), .Y(n_1136) );
NOR2xp33_ASAP7_75t_L g1137 ( .A(n_1021), .B(n_935), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_1046), .A2(n_1027), .B1(n_1114), .B2(n_1022), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1037), .Y(n_1139) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_1104), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1037), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1053), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1090), .B(n_907), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_1022), .A2(n_938), .B1(n_907), .B2(n_922), .C(n_1015), .Y(n_1144) );
NAND4xp25_ASAP7_75t_L g1145 ( .A(n_1116), .B(n_902), .C(n_921), .D(n_908), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_1097), .Y(n_1146) );
INVx3_ASAP7_75t_L g1147 ( .A(n_1036), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1091), .B(n_959), .Y(n_1148) );
AO22x1_ASAP7_75t_L g1149 ( .A1(n_1061), .A2(n_1002), .B1(n_959), .B2(n_921), .Y(n_1149) );
NOR3xp33_ASAP7_75t_SL g1150 ( .A(n_1048), .B(n_900), .C(n_930), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1053), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1091), .B(n_931), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1058), .B(n_936), .Y(n_1153) );
OAI21xp5_ASAP7_75t_L g1154 ( .A1(n_1028), .A2(n_936), .B(n_1075), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1058), .Y(n_1155) );
INVxp67_ASAP7_75t_SL g1156 ( .A(n_1019), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1052), .Y(n_1157) );
INVx2_ASAP7_75t_SL g1158 ( .A(n_1036), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1026), .B(n_1065), .Y(n_1159) );
AO31x2_ASAP7_75t_L g1160 ( .A1(n_1073), .A2(n_1025), .A3(n_1100), .B(n_1092), .Y(n_1160) );
INVx1_ASAP7_75t_SL g1161 ( .A(n_1032), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1073), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1117), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1121), .B(n_1019), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1121), .B(n_1030), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1098), .B(n_1118), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1030), .B(n_1031), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1070), .B(n_1089), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1169 ( .A1(n_1106), .A2(n_1049), .B1(n_1116), .B2(n_1078), .Y(n_1169) );
INVx2_ASAP7_75t_SL g1170 ( .A(n_1036), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1031), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1056), .B(n_1060), .Y(n_1172) );
INVxp67_ASAP7_75t_L g1173 ( .A(n_1038), .Y(n_1173) );
BUFx3_ASAP7_75t_L g1174 ( .A(n_1061), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1056), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1060), .B(n_1066), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_1066), .Y(n_1177) );
INVx1_ASAP7_75t_SL g1178 ( .A(n_1107), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1051), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1044), .B(n_1055), .Y(n_1180) );
NAND3xp33_ASAP7_75t_L g1181 ( .A(n_1080), .B(n_1084), .C(n_1078), .Y(n_1181) );
OAI31xp33_ASAP7_75t_L g1182 ( .A1(n_1079), .A2(n_1083), .A3(n_1115), .B(n_1082), .Y(n_1182) );
INVx2_ASAP7_75t_L g1183 ( .A(n_1036), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1105), .B(n_1119), .Y(n_1184) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_1102), .A2(n_1115), .B1(n_1109), .B2(n_1040), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1051), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1024), .B(n_1061), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1076), .B(n_1095), .Y(n_1188) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_1113), .A2(n_1120), .B1(n_1101), .B2(n_1029), .C(n_1068), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1054), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1051), .Y(n_1191) );
BUFx3_ASAP7_75t_L g1192 ( .A(n_1109), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1067), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1063), .B(n_1109), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1076), .B(n_1095), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_1047), .A2(n_1120), .B1(n_1111), .B2(n_1041), .Y(n_1196) );
OAI31xp33_ASAP7_75t_L g1197 ( .A1(n_1093), .A2(n_1057), .A3(n_1069), .B(n_1087), .Y(n_1197) );
AO21x2_ASAP7_75t_L g1198 ( .A1(n_1110), .A2(n_1074), .B(n_1072), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1081), .B(n_1042), .Y(n_1199) );
BUFx2_ASAP7_75t_L g1200 ( .A(n_1076), .Y(n_1200) );
AOI33xp33_ASAP7_75t_L g1201 ( .A1(n_1112), .A2(n_1042), .A3(n_1068), .B1(n_1071), .B2(n_1064), .B3(n_1050), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1062), .Y(n_1202) );
AOI21xp33_ASAP7_75t_SL g1203 ( .A1(n_1108), .A2(n_1039), .B(n_1096), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1086), .B(n_1094), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1035), .B(n_1085), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1110), .Y(n_1206) );
INVx1_ASAP7_75t_SL g1207 ( .A(n_1161), .Y(n_1207) );
OAI211xp5_ASAP7_75t_L g1208 ( .A1(n_1138), .A2(n_1077), .B(n_1108), .C(n_1088), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1124), .B(n_1099), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1171), .B(n_1175), .Y(n_1210) );
NAND4xp25_ASAP7_75t_L g1211 ( .A(n_1182), .B(n_1196), .C(n_1185), .D(n_1197), .Y(n_1211) );
AOI321xp33_ASAP7_75t_L g1212 ( .A1(n_1169), .A2(n_1189), .A3(n_1199), .B1(n_1205), .B2(n_1130), .C(n_1165), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1124), .B(n_1164), .Y(n_1213) );
OAI21xp33_ASAP7_75t_L g1214 ( .A1(n_1201), .A2(n_1133), .B(n_1127), .Y(n_1214) );
INVx2_ASAP7_75t_SL g1215 ( .A(n_1174), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1171), .B(n_1175), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1125), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1164), .B(n_1165), .Y(n_1218) );
INVxp67_ASAP7_75t_L g1219 ( .A(n_1137), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1157), .Y(n_1220) );
OR2x6_ASAP7_75t_L g1221 ( .A(n_1200), .B(n_1140), .Y(n_1221) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1122), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1140), .B(n_1125), .Y(n_1223) );
HB1xp67_ASAP7_75t_L g1224 ( .A(n_1167), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1141), .B(n_1155), .Y(n_1225) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1129), .Y(n_1226) );
OAI211xp5_ASAP7_75t_L g1227 ( .A1(n_1203), .A2(n_1181), .B(n_1173), .C(n_1145), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1163), .B(n_1166), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1141), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1142), .B(n_1151), .Y(n_1230) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_1174), .Y(n_1231) );
CKINVDCx16_ASAP7_75t_R g1232 ( .A(n_1123), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1142), .B(n_1151), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1155), .B(n_1162), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1128), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1162), .B(n_1135), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1129), .B(n_1135), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1139), .Y(n_1238) );
INVx2_ASAP7_75t_L g1239 ( .A(n_1139), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_1172), .B(n_1156), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1172), .B(n_1180), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1143), .B(n_1176), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1159), .B(n_1168), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1143), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1202), .B(n_1190), .Y(n_1245) );
INVxp67_ASAP7_75t_SL g1246 ( .A(n_1177), .Y(n_1246) );
NAND4xp25_ASAP7_75t_L g1247 ( .A(n_1184), .B(n_1178), .C(n_1131), .D(n_1144), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1180), .B(n_1176), .Y(n_1248) );
NAND4xp25_ASAP7_75t_L g1249 ( .A(n_1134), .B(n_1136), .C(n_1193), .D(n_1154), .Y(n_1249) );
NAND2x1p5_ASAP7_75t_L g1250 ( .A(n_1200), .B(n_1123), .Y(n_1250) );
AND4x1_ASAP7_75t_L g1251 ( .A(n_1150), .B(n_1132), .C(n_1204), .D(n_1195), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1146), .B(n_1194), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1146), .B(n_1194), .Y(n_1253) );
NAND4xp75_ASAP7_75t_L g1254 ( .A(n_1204), .B(n_1195), .C(n_1188), .D(n_1126), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1148), .B(n_1153), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1192), .B(n_1187), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1179), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1148), .B(n_1153), .Y(n_1258) );
AND2x4_ASAP7_75t_L g1259 ( .A(n_1188), .B(n_1192), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1152), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1152), .B(n_1183), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1183), .B(n_1206), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1206), .B(n_1191), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1158), .Y(n_1264) );
INVx1_ASAP7_75t_SL g1265 ( .A(n_1158), .Y(n_1265) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_1160), .B(n_1170), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1179), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1186), .Y(n_1268) );
NAND2xp67_ASAP7_75t_SL g1269 ( .A(n_1149), .B(n_1198), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1241), .B(n_1160), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1213), .B(n_1186), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1213), .B(n_1191), .Y(n_1272) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1257), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1255), .B(n_1160), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_1231), .Y(n_1275) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1241), .B(n_1160), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1257), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1214), .B(n_1170), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1242), .B(n_1160), .Y(n_1279) );
INVx1_ASAP7_75t_SL g1280 ( .A(n_1231), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1242), .B(n_1147), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1255), .B(n_1147), .Y(n_1282) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1267), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1258), .B(n_1147), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1248), .B(n_1149), .Y(n_1285) );
NOR3xp33_ASAP7_75t_L g1286 ( .A(n_1211), .B(n_1198), .C(n_1227), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1287 ( .A(n_1215), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1267), .Y(n_1288) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1263), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1268), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1248), .B(n_1224), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1268), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1258), .B(n_1218), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1244), .B(n_1245), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1218), .B(n_1261), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1260), .B(n_1207), .Y(n_1296) );
CKINVDCx16_ASAP7_75t_R g1297 ( .A(n_1232), .Y(n_1297) );
INVxp67_ASAP7_75t_L g1298 ( .A(n_1246), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1219), .B(n_1243), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1228), .B(n_1220), .Y(n_1300) );
AOI22xp5_ASAP7_75t_L g1301 ( .A1(n_1247), .A2(n_1208), .B1(n_1254), .B2(n_1249), .Y(n_1301) );
NOR3xp33_ASAP7_75t_L g1302 ( .A(n_1254), .B(n_1264), .C(n_1252), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1261), .B(n_1263), .Y(n_1303) );
AO21x1_ASAP7_75t_L g1304 ( .A1(n_1210), .A2(n_1216), .B(n_1240), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1210), .B(n_1216), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1251), .B(n_1233), .Y(n_1306) );
OR2x6_ASAP7_75t_L g1307 ( .A(n_1221), .B(n_1259), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1235), .B(n_1259), .Y(n_1308) );
XNOR2x1_ASAP7_75t_L g1309 ( .A(n_1256), .B(n_1253), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1293), .B(n_1209), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1293), .B(n_1209), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1291), .B(n_1256), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1291), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1295), .B(n_1259), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1271), .B(n_1233), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1295), .B(n_1223), .Y(n_1316) );
A2O1A1Ixp33_ASAP7_75t_SL g1317 ( .A1(n_1286), .A2(n_1301), .B(n_1278), .C(n_1302), .Y(n_1317) );
NAND2xp5_ASAP7_75t_SL g1318 ( .A(n_1297), .B(n_1212), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1297), .B(n_1265), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1273), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1272), .B(n_1225), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1299), .B(n_1309), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1273), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1303), .B(n_1225), .Y(n_1324) );
INVxp67_ASAP7_75t_L g1325 ( .A(n_1287), .Y(n_1325) );
BUFx2_ASAP7_75t_L g1326 ( .A(n_1307), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1274), .B(n_1223), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1273), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1283), .Y(n_1329) );
OAI32xp33_ASAP7_75t_L g1330 ( .A1(n_1306), .A2(n_1250), .A3(n_1266), .B1(n_1217), .B2(n_1229), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1283), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1283), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1305), .B(n_1289), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1289), .B(n_1230), .Y(n_1334) );
O2A1O1Ixp33_ASAP7_75t_L g1335 ( .A1(n_1298), .A2(n_1266), .B(n_1250), .C(n_1221), .Y(n_1335) );
OAI321xp33_ASAP7_75t_L g1336 ( .A1(n_1301), .A2(n_1221), .A3(n_1250), .B1(n_1262), .B2(n_1234), .C(n_1238), .Y(n_1336) );
NAND2x1_ASAP7_75t_L g1337 ( .A(n_1307), .B(n_1221), .Y(n_1337) );
INVxp67_ASAP7_75t_SL g1338 ( .A(n_1275), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1274), .B(n_1237), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1277), .Y(n_1340) );
INVx2_ASAP7_75t_SL g1341 ( .A(n_1287), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1282), .B(n_1237), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1277), .Y(n_1343) );
XNOR2xp5_ASAP7_75t_L g1344 ( .A(n_1309), .B(n_1234), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1345 ( .A(n_1294), .B(n_1236), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1300), .B(n_1236), .Y(n_1346) );
OAI21xp5_ASAP7_75t_SL g1347 ( .A1(n_1285), .A2(n_1269), .B(n_1226), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1296), .B(n_1222), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1304), .B(n_1239), .Y(n_1349) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1281), .B(n_1239), .Y(n_1350) );
OAI322xp33_ASAP7_75t_L g1351 ( .A1(n_1270), .A2(n_1269), .A3(n_1276), .B1(n_1279), .B2(n_1280), .C1(n_1290), .C2(n_1288), .Y(n_1351) );
AOI21xp5_ASAP7_75t_L g1352 ( .A1(n_1318), .A2(n_1337), .B(n_1335), .Y(n_1352) );
AOI211xp5_ASAP7_75t_L g1353 ( .A1(n_1317), .A2(n_1351), .B(n_1336), .C(n_1330), .Y(n_1353) );
OAI221xp5_ASAP7_75t_L g1354 ( .A1(n_1326), .A2(n_1337), .B1(n_1322), .B2(n_1347), .C(n_1344), .Y(n_1354) );
AO22x2_ASAP7_75t_L g1355 ( .A1(n_1341), .A2(n_1338), .B1(n_1313), .B2(n_1325), .Y(n_1355) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1312), .Y(n_1356) );
AOI21xp33_ASAP7_75t_SL g1357 ( .A1(n_1319), .A2(n_1344), .B(n_1341), .Y(n_1357) );
AOI21xp5_ASAP7_75t_L g1358 ( .A1(n_1304), .A2(n_1330), .B(n_1349), .Y(n_1358) );
BUFx2_ASAP7_75t_L g1359 ( .A(n_1307), .Y(n_1359) );
OAI21xp5_ASAP7_75t_L g1360 ( .A1(n_1280), .A2(n_1314), .B(n_1348), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1311), .B(n_1310), .Y(n_1361) );
AOI21xp5_ASAP7_75t_L g1362 ( .A1(n_1352), .A2(n_1307), .B(n_1346), .Y(n_1362) );
AOI221xp5_ASAP7_75t_L g1363 ( .A1(n_1357), .A2(n_1350), .B1(n_1333), .B2(n_1327), .C(n_1340), .Y(n_1363) );
AOI211xp5_ASAP7_75t_L g1364 ( .A1(n_1354), .A2(n_1308), .B(n_1314), .C(n_1284), .Y(n_1364) );
OR2x2_ASAP7_75t_L g1365 ( .A(n_1356), .B(n_1345), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_1359), .A2(n_1308), .B1(n_1282), .B2(n_1284), .Y(n_1366) );
NOR2x1_ASAP7_75t_L g1367 ( .A(n_1360), .B(n_1316), .Y(n_1367) );
AOI22xp5_ASAP7_75t_L g1368 ( .A1(n_1364), .A2(n_1353), .B1(n_1355), .B2(n_1358), .Y(n_1368) );
OAI211xp5_ASAP7_75t_SL g1369 ( .A1(n_1362), .A2(n_1361), .B(n_1324), .C(n_1321), .Y(n_1369) );
OAI21xp33_ASAP7_75t_L g1370 ( .A1(n_1367), .A2(n_1345), .B(n_1334), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1365), .Y(n_1371) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_1363), .A2(n_1343), .B1(n_1315), .B2(n_1323), .C(n_1328), .Y(n_1372) );
AOI22xp5_ASAP7_75t_L g1373 ( .A1(n_1368), .A2(n_1366), .B1(n_1339), .B2(n_1316), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g1374 ( .A1(n_1370), .A2(n_1339), .B1(n_1323), .B2(n_1332), .C(n_1331), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1371), .Y(n_1375) );
OAI222xp33_ASAP7_75t_L g1376 ( .A1(n_1372), .A2(n_1342), .B1(n_1320), .B2(n_1328), .C1(n_1332), .C2(n_1331), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1375), .Y(n_1377) );
NOR3xp33_ASAP7_75t_SL g1378 ( .A(n_1376), .B(n_1369), .C(n_1290), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1373), .Y(n_1379) );
AOI22xp5_ASAP7_75t_L g1380 ( .A1(n_1379), .A2(n_1374), .B1(n_1329), .B2(n_1292), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1377), .Y(n_1381) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1381), .Y(n_1382) );
OR3x1_ASAP7_75t_L g1383 ( .A(n_1380), .B(n_1378), .C(n_1292), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1382), .Y(n_1384) );
AOI21xp5_ASAP7_75t_L g1385 ( .A1(n_1384), .A2(n_1382), .B(n_1383), .Y(n_1385) );
endmodule