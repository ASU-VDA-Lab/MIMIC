module real_jpeg_23338_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_80),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_1),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_1),
.A2(n_42),
.B(n_88),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_100),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_1),
.A2(n_103),
.B1(n_200),
.B2(n_203),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_1),
.A2(n_37),
.B(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_27),
.B1(n_37),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_69),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_26),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_5),
.A2(n_27),
.B1(n_37),
.B2(n_73),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_73),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_73),
.Y(n_200)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_7),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_27),
.B1(n_37),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_8),
.A2(n_26),
.B1(n_66),
.B2(n_72),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_66),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_9),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_72),
.B1(n_78),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_27),
.B1(n_37),
.B2(n_83),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_83),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_83),
.Y(n_190)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_13),
.A2(n_27),
.B1(n_37),
.B2(n_95),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_15),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_19),
.B(n_114),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_84),
.C(n_101),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_20),
.A2(n_21),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_22),
.B(n_56),
.C(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_23),
.A2(n_38),
.B1(n_39),
.B2(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_23),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.A3(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_23)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_27),
.A2(n_37),
.B1(n_59),
.B2(n_63),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_27),
.B(n_35),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_30),
.A2(n_31),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_33),
.A2(n_35),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_35),
.A2(n_61),
.B(n_90),
.C(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_35),
.B(n_91),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_35),
.B(n_108),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_37),
.A2(n_59),
.A3(n_61),
.B1(n_216),
.B2(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_49),
.B2(n_53),
.Y(n_39)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_40),
.B(n_109),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_40),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_41),
.A2(n_42),
.B1(n_88),
.B2(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_41),
.B(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_47),
.A2(n_130),
.B(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_50),
.A2(n_103),
.B1(n_190),
.B2(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_52),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_70),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_65),
.B(n_67),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_65),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_57),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_57),
.A2(n_99),
.B1(n_100),
.B2(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_58),
.A2(n_124),
.B1(n_154),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_58)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_61),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_60),
.B(n_63),
.Y(n_223)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_68),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_74),
.B1(n_80),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_76),
.B1(n_82),
.B2(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_84),
.B(n_101),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_96),
.C(n_98),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_98),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B(n_93),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_86),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_86),
.A2(n_173),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_86),
.A2(n_181),
.B1(n_182),
.B2(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_111),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_91),
.A2(n_135),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_92),
.B(n_181),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_110),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_110),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_103),
.A2(n_131),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_103),
.A2(n_105),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_128),
.B2(n_137),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_127),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_128),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_135),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_163),
.B(n_251),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_160),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_145),
.B(n_160),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_148),
.Y(n_249)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_152),
.B(n_234),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_245),
.B(n_250),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_229),
.B(n_244),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_209),
.B(n_228),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_186),
.B(n_208),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_176),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_183),
.C(n_184),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_196),
.B(n_207),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_194),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_201),
.B(n_206),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_198),
.B(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_221),
.B1(n_226),
.B2(n_227),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_212)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_220),
.C(n_226),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_231),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_239),
.C(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);


endmodule