module fake_jpeg_4874_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx13_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_12),
.Y(n_36)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_21),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_21),
.B1(n_24),
.B2(n_18),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_46),
.B1(n_20),
.B2(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_21),
.B1(n_24),
.B2(n_13),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_17),
.B1(n_15),
.B2(n_19),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_54),
.B1(n_56),
.B2(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_15),
.B1(n_19),
.B2(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_70),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_40),
.B1(n_35),
.B2(n_46),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_53),
.B1(n_50),
.B2(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_71),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_43),
.B1(n_27),
.B2(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_27),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_79),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_78),
.B(n_65),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_33),
.B1(n_30),
.B2(n_41),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_58),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_64),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.C(n_88),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_90),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_69),
.C(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_37),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.C(n_85),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_37),
.C(n_60),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_22),
.C(n_37),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

OAI22x1_ASAP7_75t_R g95 ( 
.A1(n_78),
.A2(n_33),
.B1(n_30),
.B2(n_41),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_103),
.C(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_104),
.B(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_72),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_76),
.B1(n_83),
.B2(n_73),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_78),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_83),
.B1(n_95),
.B2(n_58),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_28),
.B1(n_22),
.B2(n_4),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_1),
.B(n_4),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_22),
.C(n_8),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_112),
.A2(n_11),
.B(n_7),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_7),
.B(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_119),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_6),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_108),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_107),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_118),
.B(n_109),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_111),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_121),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_8),
.C(n_10),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_129),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_1),
.B1(n_5),
.B2(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_5),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_133),
.B(n_128),
.CI(n_132),
.CON(n_135),
.SN(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);


endmodule