module fake_jpeg_6252_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_43),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_27),
.B(n_20),
.C(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_27),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_24),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_90),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_63),
.B1(n_74),
.B2(n_53),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_97),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_28),
.B1(n_18),
.B2(n_29),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_65),
.B1(n_70),
.B2(n_69),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_92),
.B1(n_49),
.B2(n_54),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_31),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_61),
.B1(n_60),
.B2(n_65),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_104),
.B(n_107),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_51),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_78),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_124),
.B1(n_128),
.B2(n_86),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_57),
.B(n_66),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_126),
.B(n_108),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_85),
.B1(n_79),
.B2(n_97),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_63),
.B1(n_55),
.B2(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_118),
.B1(n_127),
.B2(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_67),
.B1(n_40),
.B2(n_38),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_91),
.B1(n_75),
.B2(n_81),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_76),
.A2(n_67),
.B1(n_46),
.B2(n_40),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_91),
.B1(n_75),
.B2(n_87),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_133),
.B1(n_144),
.B2(n_154),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_102),
.B(n_1),
.Y(n_185)
);

AO21x2_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_67),
.B(n_21),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_145),
.B1(n_116),
.B2(n_21),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_141),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_99),
.B(n_96),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_34),
.B(n_26),
.Y(n_178)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_96),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_99),
.B1(n_76),
.B2(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_150),
.B1(n_125),
.B2(n_111),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_31),
.C(n_21),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_119),
.B(n_130),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_31),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_112),
.A2(n_34),
.B1(n_26),
.B2(n_23),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_17),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_34),
.B1(n_26),
.B2(n_23),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_178),
.B(n_182),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_114),
.B1(n_129),
.B2(n_107),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_164),
.B1(n_166),
.B2(n_171),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_128),
.C(n_104),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_173),
.Y(n_186)
);

AOI22x1_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_124),
.B1(n_86),
.B2(n_21),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_127),
.B1(n_117),
.B2(n_125),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_174),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_184),
.B1(n_135),
.B2(n_174),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_170),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_34),
.B1(n_23),
.B2(n_26),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_111),
.C(n_100),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_135),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_102),
.C(n_86),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_181),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_23),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_173),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_206),
.B1(n_161),
.B2(n_182),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_210),
.C(n_186),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_135),
.B1(n_155),
.B2(n_133),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_196),
.B1(n_202),
.B2(n_116),
.Y(n_227)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_199),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_157),
.B1(n_131),
.B2(n_138),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_138),
.B(n_137),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_198),
.B(n_177),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_140),
.B(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_148),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_201),
.B(n_182),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_154),
.B1(n_145),
.B2(n_150),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_164),
.B1(n_158),
.B2(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_186),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_151),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_162),
.CI(n_168),
.CON(n_213),
.SN(n_213)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_15),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_214),
.A2(n_222),
.B(n_193),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_195),
.B1(n_201),
.B2(n_199),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_215),
.A2(n_219),
.B1(n_223),
.B2(n_226),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_224),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_175),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_231),
.C(n_234),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_160),
.B(n_165),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_165),
.B1(n_163),
.B2(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_163),
.B1(n_151),
.B2(n_167),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

OAI22x1_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_142),
.B1(n_116),
.B2(n_3),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_232),
.B1(n_197),
.B2(n_194),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_187),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_229),
.A2(n_238),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_247),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_248),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_205),
.C(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_4),
.Y(n_250)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_252),
.B(n_260),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_16),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_254),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_15),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_229),
.C(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_213),
.B(n_216),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_224),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_276),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_241),
.B(n_256),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_235),
.B1(n_227),
.B2(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_259),
.C(n_253),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_280),
.C(n_254),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_219),
.B1(n_230),
.B2(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_274),
.B1(n_278),
.B2(n_257),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_261),
.A2(n_215),
.B1(n_213),
.B2(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_240),
.B(n_5),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_275),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_7),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_239),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_279),
.B(n_251),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_7),
.C(n_8),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_244),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_284),
.B(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_244),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_291),
.C(n_296),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_266),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_11),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_270),
.B1(n_278),
.B2(n_277),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_251),
.C(n_249),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_292),
.B(n_9),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_249),
.C(n_247),
.Y(n_296)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_243),
.C(n_10),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_265),
.C(n_264),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_305),
.C(n_307),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_274),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_311),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_306),
.B1(n_288),
.B2(n_284),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_268),
.C(n_269),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_262),
.C(n_10),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_309),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_9),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_10),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_11),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_285),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_287),
.B1(n_290),
.B2(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_320),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_295),
.B1(n_289),
.B2(n_13),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_300),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_11),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_12),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_12),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_299),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_331),
.B(n_14),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_299),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_330),
.A2(n_313),
.B(n_316),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_14),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_334),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_313),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_335),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_314),
.B(n_322),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_336),
.B(n_337),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_338),
.A2(n_328),
.B(n_327),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_340),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_325),
.Y(n_343)
);

AOI321xp33_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_339),
.C(n_335),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_12),
.B(n_13),
.Y(n_345)
);


endmodule