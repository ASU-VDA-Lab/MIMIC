module fake_jpeg_29113_n_45 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_13),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_7),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_8),
.B1(n_10),
.B2(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_22),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_4),
.B(n_5),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_25),
.B2(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_36),
.C(n_37),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_36),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_29),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_39),
.B(n_38),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_35),
.B(n_30),
.Y(n_45)
);


endmodule