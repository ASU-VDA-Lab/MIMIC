module fake_jpeg_15347_n_117 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_117);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_0),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_20),
.C(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_32),
.Y(n_37)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_24),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_25),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_15),
.B1(n_27),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_50),
.B1(n_51),
.B2(n_17),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_15),
.B1(n_28),
.B2(n_17),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_48),
.B1(n_58),
.B2(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_55),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_15),
.B1(n_18),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_17),
.B1(n_29),
.B2(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_32),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_13),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_66),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_31),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_73),
.C(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_70),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_35),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_74),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_35),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_80),
.C(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_38),
.C(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_46),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_12),
.C(n_44),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_65),
.C(n_72),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

AO221x1_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_57),
.B1(n_22),
.B2(n_4),
.C(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_12),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_20),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_85),
.B1(n_20),
.B2(n_12),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_57),
.C(n_12),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_101),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_4),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_100),
.B1(n_96),
.B2(n_99),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_105),
.B(n_106),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_11),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_109),
.A2(n_110),
.B(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_113),
.B(n_4),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_111),
.Y(n_117)
);


endmodule