module fake_jpeg_25123_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_SL g33 ( 
.A(n_17),
.Y(n_33)
);

OR2x4_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_17),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx9p33_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_16),
.B1(n_13),
.B2(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_54),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_60),
.B1(n_24),
.B2(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_58),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_37),
.B1(n_41),
.B2(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_20),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_38),
.C(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_73),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_37),
.B1(n_39),
.B2(n_29),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_31),
.B1(n_29),
.B2(n_18),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_13),
.B1(n_19),
.B2(n_24),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_31),
.B1(n_47),
.B2(n_38),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_79),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_47),
.B1(n_38),
.B2(n_44),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_86),
.B1(n_44),
.B2(n_63),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_44),
.B1(n_27),
.B2(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_58),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_27),
.C(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_59),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_1),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_1),
.B(n_2),
.Y(n_115)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_67),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_82),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_86),
.B(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_109),
.C(n_112),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_85),
.B(n_81),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_85),
.C(n_84),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_116),
.C(n_92),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_82),
.B(n_62),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_59),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_127),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_87),
.B1(n_93),
.B2(n_96),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_120),
.B1(n_106),
.B2(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_90),
.C(n_87),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_110),
.C(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_138),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_120),
.C(n_108),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_142),
.C(n_130),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_129),
.B1(n_132),
.B2(n_126),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_107),
.B(n_112),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_133),
.B(n_126),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_109),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_122),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_94),
.C(n_101),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_145),
.A2(n_143),
.B(n_140),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_99),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_149),
.C(n_135),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_57),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_124),
.C(n_133),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_115),
.B(n_98),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_152),
.B(n_18),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_115),
.B1(n_100),
.B2(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_153),
.B(n_154),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_138),
.C(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_152),
.B(n_18),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_64),
.A3(n_95),
.B1(n_63),
.B2(n_57),
.C1(n_61),
.C2(n_59),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_151),
.A3(n_49),
.B1(n_61),
.B2(n_27),
.C1(n_5),
.C2(n_7),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_1),
.B(n_2),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.C(n_3),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_151),
.A3(n_61),
.B1(n_3),
.B2(n_4),
.C1(n_8),
.C2(n_9),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_169),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.C(n_163),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_3),
.B(n_4),
.C(n_8),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_27),
.C2(n_171),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_11),
.B(n_27),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);


endmodule