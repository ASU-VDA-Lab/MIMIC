module fake_jpeg_1908_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_1),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_75),
.A2(n_52),
.B1(n_51),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_49),
.B1(n_53),
.B2(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_66),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_62),
.B1(n_59),
.B2(n_69),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_61),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_106),
.B1(n_8),
.B2(n_9),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_89),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_54),
.B(n_48),
.C(n_46),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_125)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_77),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_77),
.B1(n_69),
.B2(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_1),
.Y(n_117)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_53),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_98),
.C(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_53),
.B1(n_62),
.B2(n_59),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_84),
.B(n_82),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_82),
.A3(n_65),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_117),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_30),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_124),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_89),
.B1(n_81),
.B2(n_91),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_129),
.B1(n_24),
.B2(n_42),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_2),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_127),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_7),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_134),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_103),
.B(n_10),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_128),
.B(n_17),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_26),
.B1(n_31),
.B2(n_36),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_23),
.C(n_41),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_145),
.B1(n_149),
.B2(n_40),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_37),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_150),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_161),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_159),
.B(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_19),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_21),
.B(n_22),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_44),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_38),
.C(n_39),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_141),
.C(n_162),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_159),
.B1(n_158),
.B2(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_178),
.C(n_163),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_157),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_176),
.B1(n_154),
.B2(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_164),
.C(n_156),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_153),
.C(n_166),
.Y(n_188)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_181),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_187),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_185),
.C(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_182),
.C(n_176),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_186),
.C(n_165),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_171),
.Y(n_195)
);


endmodule