module fake_jpeg_14219_n_487 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_487);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_487;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_52),
.Y(n_114)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_70),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_61),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_28),
.B(n_17),
.C(n_16),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_47),
.C(n_43),
.Y(n_133)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_26),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_69),
.B(n_80),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_84),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_0),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_4),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_4),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_90),
.Y(n_111)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_94),
.Y(n_118)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_41),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_30),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_50),
.A2(n_49),
.B1(n_48),
.B2(n_37),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_100),
.A2(n_108),
.B1(n_116),
.B2(n_19),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_24),
.B(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_103),
.B(n_144),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_30),
.B1(n_25),
.B2(n_48),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_110),
.B(n_52),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_58),
.A2(n_49),
.B1(n_30),
.B2(n_43),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_113),
.A2(n_134),
.B1(n_139),
.B2(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_32),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_137),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_54),
.A2(n_47),
.B1(n_43),
.B2(n_32),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_133),
.B(n_19),
.C(n_41),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_53),
.A2(n_47),
.B1(n_32),
.B2(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_57),
.B(n_21),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_85),
.A2(n_23),
.B1(n_21),
.B2(n_31),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_52),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_71),
.B(n_21),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_36),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_23),
.B1(n_31),
.B2(n_33),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_89),
.Y(n_162)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_67),
.B1(n_62),
.B2(n_51),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_158),
.A2(n_120),
.B1(n_135),
.B2(n_72),
.Y(n_213)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_145),
.CON(n_159),
.SN(n_159)
);

NOR3xp33_ASAP7_75t_L g225 ( 
.A(n_159),
.B(n_188),
.C(n_192),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_111),
.A2(n_23),
.B(n_52),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_160),
.B(n_162),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_109),
.B(n_76),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_165),
.B(n_174),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_61),
.B1(n_93),
.B2(n_92),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_142),
.B(n_112),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_101),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_167),
.B(n_172),
.Y(n_251)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_169),
.B(n_177),
.Y(n_233)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_75),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_184),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_118),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_104),
.B(n_33),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_175),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_117),
.B(n_59),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_178),
.Y(n_220)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_128),
.B(n_59),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_181),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_182),
.B(n_185),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_89),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_183),
.B(n_190),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_110),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_146),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_186),
.Y(n_221)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_189),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_81),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_201),
.B1(n_203),
.B2(n_206),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_36),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_194),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_36),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_195),
.B(n_200),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_107),
.A2(n_87),
.B(n_18),
.C(n_41),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_199),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_155),
.C(n_163),
.Y(n_211)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_112),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_124),
.Y(n_203)
);

BUFx16f_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_204),
.B(n_88),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_27),
.B1(n_19),
.B2(n_18),
.Y(n_235)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_207),
.A2(n_114),
.B1(n_140),
.B2(n_136),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_131),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_211),
.C(n_189),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_213),
.A2(n_216),
.B1(n_218),
.B2(n_224),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_214),
.A2(n_14),
.B(n_15),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_155),
.A2(n_105),
.B1(n_83),
.B2(n_96),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_205),
.A2(n_105),
.B1(n_65),
.B2(n_63),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_102),
.B1(n_135),
.B2(n_120),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_219),
.A2(n_230),
.B1(n_244),
.B2(n_188),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_131),
.C(n_142),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_222),
.B(n_249),
.C(n_8),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_82),
.B1(n_122),
.B2(n_102),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_169),
.A2(n_122),
.B1(n_119),
.B2(n_132),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_235),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_159),
.A2(n_119),
.B1(n_132),
.B2(n_136),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_171),
.B1(n_177),
.B2(n_157),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_114),
.B1(n_140),
.B2(n_33),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_237),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_166),
.A2(n_27),
.B1(n_18),
.B2(n_56),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_240),
.A2(n_243),
.B1(n_252),
.B2(n_14),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_27),
.B1(n_56),
.B2(n_22),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_177),
.A2(n_74),
.B1(n_22),
.B2(n_6),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_22),
.C(n_5),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_197),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_185),
.B(n_206),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_255),
.A2(n_279),
.B(n_285),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_256),
.A2(n_227),
.B1(n_221),
.B2(n_238),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_208),
.B(n_201),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_257),
.B(n_262),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_164),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_186),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_271),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_234),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_260),
.B(n_275),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_168),
.B1(n_175),
.B2(n_173),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_266),
.B1(n_282),
.B2(n_243),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_199),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_264),
.B(n_274),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_272),
.C(n_284),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_230),
.A2(n_178),
.B1(n_187),
.B2(n_154),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_214),
.A2(n_182),
.B(n_191),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_288),
.B(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g271 ( 
.A1(n_218),
.A2(n_161),
.B(n_170),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_210),
.B(n_204),
.C(n_207),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_204),
.B(n_6),
.C(n_7),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_273),
.B(n_276),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_156),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_232),
.B(n_4),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_233),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_224),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_278),
.A2(n_298),
.B1(n_212),
.B2(n_226),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_8),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_290),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_215),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_245),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_211),
.B(n_9),
.C(n_10),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_9),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_232),
.B(n_215),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_286),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_222),
.B(n_9),
.C(n_11),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_292),
.C(n_281),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_223),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_251),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_289),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_233),
.B(n_223),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_249),
.B(n_14),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_295),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_219),
.B(n_231),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_235),
.B(n_15),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_253),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_296),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_253),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_297),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_216),
.A2(n_15),
.B1(n_228),
.B2(n_213),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_308),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_220),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_307),
.C(n_316),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_302),
.A2(n_304),
.B1(n_314),
.B2(n_322),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_252),
.B1(n_240),
.B2(n_235),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_220),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_235),
.B1(n_244),
.B2(n_225),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_333),
.Y(n_342)
);

OAI22x1_ASAP7_75t_SL g314 ( 
.A1(n_293),
.A2(n_235),
.B1(n_245),
.B2(n_248),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_237),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_284),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_237),
.C(n_248),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_323),
.C(n_269),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_259),
.B(n_237),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_267),
.A2(n_212),
.B(n_209),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_331),
.B(n_266),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_221),
.B1(n_238),
.B2(n_217),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_325),
.A2(n_327),
.B1(n_332),
.B2(n_336),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_271),
.A2(n_217),
.B1(n_246),
.B2(n_209),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_291),
.A2(n_241),
.B(n_246),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_271),
.A2(n_15),
.B1(n_242),
.B2(n_270),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_268),
.A2(n_298),
.B1(n_255),
.B2(n_260),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_271),
.A2(n_258),
.B1(n_263),
.B2(n_296),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_304),
.A2(n_268),
.B1(n_255),
.B2(n_294),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_341),
.A2(n_314),
.B1(n_299),
.B2(n_308),
.Y(n_374)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_257),
.A3(n_286),
.B1(n_280),
.B2(n_264),
.Y(n_343)
);

AOI221xp5_ASAP7_75t_L g373 ( 
.A1(n_343),
.A2(n_335),
.B1(n_301),
.B2(n_309),
.C(n_330),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_337),
.Y(n_344)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_281),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_347),
.C(n_352),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_349),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_297),
.Y(n_348)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_258),
.Y(n_349)
);

AO32x1_ASAP7_75t_L g350 ( 
.A1(n_319),
.A2(n_269),
.A3(n_273),
.B1(n_288),
.B2(n_258),
.Y(n_350)
);

AND2x4_ASAP7_75t_SL g394 ( 
.A(n_350),
.B(n_273),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_351),
.B(n_361),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_274),
.C(n_279),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_315),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_355),
.Y(n_389)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_354),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_320),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_289),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_356),
.B(n_359),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_287),
.C(n_283),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_363),
.C(n_312),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_328),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_368),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_303),
.B(n_285),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_319),
.A2(n_335),
.B(n_331),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_360),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_275),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_313),
.Y(n_362)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_283),
.C(n_261),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_307),
.B(n_282),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_365),
.Y(n_388)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_369),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_305),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_378),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_373),
.B(n_355),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_374),
.A2(n_380),
.B1(n_384),
.B2(n_332),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_367),
.A2(n_368),
.B1(n_342),
.B2(n_338),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_339),
.B1(n_369),
.B2(n_364),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_316),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_341),
.A2(n_299),
.B1(n_329),
.B2(n_301),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_329),
.B1(n_321),
.B2(n_318),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_340),
.B(n_323),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_390),
.B(n_396),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_393),
.C(n_363),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_312),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_349),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_357),
.B(n_302),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_398),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_402),
.B1(n_374),
.B2(n_384),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_352),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_405),
.Y(n_436)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_401),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_406),
.C(n_408),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_360),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_358),
.C(n_342),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_382),
.B(n_359),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_407),
.B(n_413),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_348),
.C(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_346),
.C(n_338),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_412),
.C(n_414),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_354),
.C(n_339),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_344),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_353),
.C(n_350),
.Y(n_414)
);

NOR3xp33_ASAP7_75t_SL g415 ( 
.A(n_372),
.B(n_350),
.C(n_343),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_415),
.B(n_417),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_416),
.A2(n_375),
.B1(n_392),
.B2(n_381),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_362),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_306),
.C(n_362),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_394),
.C(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_411),
.A2(n_377),
.B(n_380),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_421),
.A2(n_425),
.B(n_405),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_423),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_424),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_412),
.A2(n_377),
.B(n_395),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_433),
.Y(n_441)
);

AOI321xp33_ASAP7_75t_L g432 ( 
.A1(n_414),
.A2(n_395),
.A3(n_394),
.B1(n_388),
.B2(n_377),
.C(n_376),
.Y(n_432)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_437),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_383),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_406),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_439),
.B(n_451),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_404),
.C(n_403),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_450),
.C(n_437),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_408),
.B(n_418),
.Y(n_442)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_306),
.Y(n_444)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_423),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_428),
.A2(n_409),
.B1(n_400),
.B2(n_283),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_448),
.A2(n_421),
.B1(n_434),
.B2(n_424),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_409),
.C(n_261),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_438),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_278),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_452),
.B(n_426),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_456),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_445),
.A2(n_435),
.B(n_432),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_426),
.C(n_430),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_461),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_446),
.B(n_427),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_460),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_449),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_427),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_444),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_436),
.C(n_435),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_463),
.A2(n_447),
.B(n_450),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_466),
.A2(n_472),
.B1(n_464),
.B2(n_430),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_446),
.C(n_443),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_469),
.C(n_458),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_436),
.C(n_448),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_453),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_473),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_474),
.B(n_476),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_475),
.A2(n_477),
.B1(n_463),
.B2(n_467),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_478),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_479),
.B(n_481),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_480),
.A2(n_478),
.B(n_471),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_482),
.A2(n_454),
.B(n_470),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_483),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_456),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_486),
.Y(n_487)
);


endmodule