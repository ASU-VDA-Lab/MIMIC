module fake_jpeg_29765_n_95 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_7),
.B(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_30),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_30),
.B1(n_26),
.B2(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_26),
.B1(n_42),
.B2(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_59),
.B1(n_45),
.B2(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_31),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_33),
.C(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_66),
.B1(n_70),
.B2(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_52),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_46),
.B1(n_40),
.B2(n_49),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_37),
.C(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_39),
.B1(n_50),
.B2(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_75),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_56),
.C(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_79),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_76),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_77),
.B1(n_78),
.B2(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

AOI322xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_73),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_5),
.C2(n_8),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_83),
.B1(n_57),
.B2(n_8),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_9),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_5),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_89),
.B(n_10),
.Y(n_91)
);

OAI21x1_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_20),
.B(n_24),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_90),
.A2(n_19),
.B(n_23),
.C(n_12),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_10),
.B1(n_11),
.B2(n_15),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_93),
.B(n_22),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_94),
.Y(n_95)
);


endmodule