module fake_jpeg_21343_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_18),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_40),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_16),
.C(n_26),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_43),
.C(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_31),
.B1(n_22),
.B2(n_34),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_57),
.B1(n_58),
.B2(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_31),
.B1(n_22),
.B2(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_22),
.B1(n_32),
.B2(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_30),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_67),
.B(n_80),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_90),
.Y(n_110)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_86),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_29),
.B1(n_38),
.B2(n_23),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_38),
.B1(n_29),
.B2(n_27),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_29),
.B1(n_24),
.B2(n_30),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_79),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_29),
.B1(n_35),
.B2(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_54),
.B1(n_49),
.B2(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_23),
.B1(n_35),
.B2(n_27),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_93),
.B1(n_99),
.B2(n_101),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_33),
.B(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_33),
.B1(n_28),
.B2(n_21),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_20),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_25),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_28),
.B1(n_21),
.B2(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_103),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_43),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_43),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_108),
.B(n_115),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_40),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_123),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_131),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g123 ( 
.A1(n_79),
.A2(n_39),
.B1(n_43),
.B2(n_26),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_68),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_18),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_90),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_104),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_18),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_142),
.Y(n_175)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_167),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_66),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_141),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_66),
.C(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_147),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_73),
.B(n_106),
.C(n_74),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_154),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_148),
.B(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_74),
.B1(n_85),
.B2(n_73),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_126),
.B1(n_120),
.B2(n_128),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_70),
.B1(n_69),
.B2(n_65),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_161),
.B1(n_164),
.B2(n_129),
.Y(n_172)
);

AO21x2_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_101),
.B(n_103),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_123),
.B(n_126),
.C(n_115),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_104),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_153),
.B(n_11),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_91),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_160),
.Y(n_195)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_107),
.A2(n_86),
.B1(n_84),
.B2(n_20),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_20),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_25),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_123),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_118),
.A2(n_28),
.B1(n_26),
.B2(n_105),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_28),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_168),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_108),
.A2(n_26),
.B(n_1),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_120),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_187),
.B(n_190),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_132),
.B1(n_8),
.B2(n_3),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_129),
.B1(n_118),
.B2(n_131),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_186),
.B1(n_152),
.B2(n_139),
.Y(n_207)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_162),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_144),
.A2(n_128),
.B(n_114),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_114),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_152),
.B1(n_125),
.B2(n_94),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_121),
.B(n_113),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_196),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_146),
.A2(n_125),
.B(n_137),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_163),
.B(n_141),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_146),
.B(n_14),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_145),
.B(n_11),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_140),
.B(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_0),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_127),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_208),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_201),
.B(n_220),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_152),
.C(n_109),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_211),
.C(n_221),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_215),
.B1(n_176),
.B2(n_171),
.Y(n_235)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_198),
.C(n_170),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_212),
.B(n_223),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_132),
.B1(n_9),
.B2(n_4),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_9),
.C(n_14),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_7),
.B1(n_13),
.B2(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_15),
.C(n_7),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_9),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_225),
.A2(n_226),
.B1(n_196),
.B2(n_171),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_5),
.B(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_245),
.B1(n_218),
.B2(n_169),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_184),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_246),
.B(n_200),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_186),
.B1(n_172),
.B2(n_187),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_214),
.B(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_244),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_177),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_207),
.A2(n_186),
.B1(n_183),
.B2(n_169),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_211),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_265),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_219),
.B1(n_186),
.B2(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_253),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_259),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_186),
.B1(n_231),
.B2(n_227),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_255),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_201),
.C(n_203),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_261),
.C(n_262),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_192),
.C(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_220),
.C(n_209),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_221),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_266),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_274),
.B(n_279),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_247),
.C(n_229),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_277),
.C(n_278),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_246),
.C(n_239),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_185),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_233),
.C(n_217),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_265),
.C(n_252),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_210),
.B1(n_259),
.B2(n_260),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_285),
.B1(n_272),
.B2(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_250),
.C(n_251),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_229),
.B1(n_256),
.B2(n_241),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_264),
.B(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_191),
.B(n_213),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_263),
.B1(n_216),
.B2(n_195),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_289),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_216),
.B1(n_197),
.B2(n_213),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_173),
.C(n_179),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_269),
.C(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_299),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_272),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_295),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_224),
.B1(n_173),
.B2(n_234),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_230),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_298),
.A2(n_282),
.B(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_291),
.C(n_284),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_295),
.B(n_293),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_303),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_180),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_307),
.B(n_297),
.Y(n_309)
);

NAND4xp25_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_234),
.C(n_297),
.D(n_193),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_304),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_309),
.B(n_6),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_6),
.B(n_10),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_12),
.B(n_15),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_312),
.Y(n_313)
);


endmodule