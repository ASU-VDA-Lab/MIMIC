module fake_netlist_5_945_n_196 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_196);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_196;

wire n_137;
wire n_168;
wire n_164;
wire n_191;
wire n_91;
wire n_82;
wire n_122;
wire n_194;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_98;
wire n_66;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_195;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_193;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_192;
wire n_53;
wire n_160;
wire n_188;
wire n_190;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_64;
wire n_77;
wire n_102;
wire n_161;
wire n_106;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_141;
wire n_97;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_R g55 ( 
.A(n_41),
.B(n_35),
.Y(n_55)
);

INVxp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_R g66 ( 
.A(n_46),
.B(n_0),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_48),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_52),
.B1(n_51),
.B2(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_65),
.B(n_70),
.Y(n_91)
);

OAI21x1_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_73),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_67),
.Y(n_93)
);

NAND2x1p5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_72),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_76),
.B(n_51),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_68),
.B(n_60),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_73),
.B(n_49),
.C(n_45),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_86),
.B1(n_87),
.B2(n_82),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_78),
.B1(n_79),
.B2(n_84),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_45),
.B(n_43),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_R g114 ( 
.A(n_103),
.B(n_99),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_93),
.B1(n_91),
.B2(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_113),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_108),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_116),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_112),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_111),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_111),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_95),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_91),
.Y(n_132)
);

AND2x4_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_117),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_95),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_109),
.B1(n_114),
.B2(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_109),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

XNOR2x2_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_127),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_127),
.B1(n_128),
.B2(n_124),
.Y(n_145)
);

OAI221xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_102),
.B1(n_43),
.B2(n_40),
.C(n_90),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_130),
.B1(n_40),
.B2(n_128),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_130),
.B1(n_128),
.B2(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_128),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_133),
.B(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_137),
.Y(n_153)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_145),
.Y(n_154)
);

NAND2x1_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_137),
.Y(n_155)
);

AOI31xp33_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_139),
.A3(n_60),
.B(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_139),
.Y(n_159)
);

AOI321xp33_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_146),
.A3(n_144),
.B1(n_97),
.B2(n_90),
.C(n_84),
.Y(n_160)
);

OAI321xp33_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_80),
.A3(n_125),
.B1(n_97),
.B2(n_66),
.C(n_88),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_158),
.A3(n_151),
.B1(n_152),
.B2(n_153),
.C(n_155),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_133),
.B1(n_88),
.B2(n_117),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_66),
.B1(n_88),
.B2(n_81),
.C(n_4),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_1),
.C(n_2),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_117),
.B1(n_131),
.B2(n_81),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_81),
.C(n_131),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_131),
.C(n_75),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_162),
.B(n_81),
.Y(n_170)
);

OAI211xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_3),
.Y(n_172)
);

NOR4xp75_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_167),
.B1(n_161),
.B2(n_11),
.C(n_12),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_74),
.C(n_10),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_74),
.B1(n_106),
.B2(n_101),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

OAI221xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.C(n_17),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_R g180 ( 
.A(n_173),
.B(n_19),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_106),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_106),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_176),
.B1(n_101),
.B2(n_96),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

NAND4xp25_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_20),
.C(n_22),
.D(n_24),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_190),
.Y(n_192)
);

OAI22x1_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_185),
.B1(n_179),
.B2(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_191),
.B1(n_193),
.B2(n_187),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_186),
.B1(n_188),
.B2(n_191),
.Y(n_196)
);


endmodule