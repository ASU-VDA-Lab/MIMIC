module fake_jpeg_30816_n_78 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_32),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_28),
.B1(n_26),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_56),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_10),
.A3(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_58),
.B(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_0),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_50),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_61),
.B1(n_6),
.B2(n_8),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_3),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_65),
.B1(n_53),
.B2(n_59),
.Y(n_69)
);

XNOR2x1_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_9),
.Y(n_70)
);

OAI21x1_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_70),
.B(n_64),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B1(n_70),
.B2(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_62),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_66),
.C(n_15),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_13),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_17),
.Y(n_78)
);


endmodule