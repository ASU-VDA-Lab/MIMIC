module fake_jpeg_24526_n_20 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_20;

wire n_13;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

AND2x2_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_9),
.Y(n_11)
);

BUFx2_ASAP7_75t_SL g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.C(n_8),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_0),
.B(n_2),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_4),
.B(n_5),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_18),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_10),
.C(n_0),
.Y(n_20)
);


endmodule