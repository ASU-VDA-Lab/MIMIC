module fake_netlist_1_12366_n_724 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_724);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_724;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g108 ( .A(n_83), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_39), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_58), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_100), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_86), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
BUFx5_ASAP7_75t_L g116 ( .A(n_73), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_3), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_54), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_28), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_49), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_18), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_50), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_68), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_102), .Y(n_124) );
INVxp33_ASAP7_75t_L g125 ( .A(n_55), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_1), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_94), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_85), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_20), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_44), .Y(n_130) );
OR2x2_ASAP7_75t_L g131 ( .A(n_23), .B(n_18), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_4), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_74), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_35), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_66), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_67), .Y(n_136) );
NOR2xp67_ASAP7_75t_L g137 ( .A(n_13), .B(n_5), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_26), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_88), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_47), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_12), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_75), .Y(n_143) );
INVxp33_ASAP7_75t_SL g144 ( .A(n_16), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_27), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_96), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_33), .Y(n_147) );
INVxp67_ASAP7_75t_SL g148 ( .A(n_57), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_31), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_56), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_87), .Y(n_152) );
AOI22x1_ASAP7_75t_SL g153 ( .A1(n_138), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_153) );
INVx5_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_151), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
INVxp67_ASAP7_75t_SL g159 ( .A(n_115), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_109), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_150), .B(n_0), .Y(n_162) );
AND2x6_ASAP7_75t_L g163 ( .A(n_110), .B(n_29), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_114), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_116), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_119), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_116), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_119), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_129), .B(n_2), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_163), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_160), .B(n_122), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_172), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_157), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_157), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_154), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_161), .Y(n_181) );
INVx6_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_163), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_172), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_167), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_160), .B(n_122), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_166), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_158), .B(n_125), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_154), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_158), .B(n_133), .Y(n_192) );
INVx1_ASAP7_75t_SL g193 ( .A(n_164), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
AND2x6_ASAP7_75t_L g195 ( .A(n_162), .B(n_123), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_156), .B(n_133), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_159), .B(n_111), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_160), .B(n_156), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_176), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_176), .Y(n_200) );
NOR2x2_ASAP7_75t_L g201 ( .A(n_185), .B(n_153), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_190), .B(n_164), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_190), .B(n_162), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_195), .B(n_162), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_195), .B(n_162), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_195), .B(n_162), .Y(n_210) );
BUFx12f_ASAP7_75t_L g211 ( .A(n_195), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_197), .B(n_176), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_195), .A2(n_172), .B1(n_163), .B2(n_159), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_198), .A2(n_168), .B(n_170), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_176), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_193), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_184), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_184), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_195), .B(n_160), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_195), .B(n_160), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_195), .B(n_165), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_197), .B(n_172), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_193), .B(n_165), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_184), .B(n_172), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_184), .Y(n_226) );
NOR3xp33_ASAP7_75t_SL g227 ( .A(n_192), .B(n_121), .C(n_140), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_174), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_197), .B(n_169), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_173), .Y(n_230) );
NOR2x2_ASAP7_75t_L g231 ( .A(n_192), .B(n_153), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_177), .B(n_171), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_178), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_205), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_224), .B(n_198), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_216), .Y(n_236) );
HB1xp67_ASAP7_75t_SL g237 ( .A(n_208), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_199), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_211), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g241 ( .A1(n_203), .A2(n_196), .B(n_175), .C(n_186), .Y(n_241) );
INVxp67_ASAP7_75t_SL g242 ( .A(n_208), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_208), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_204), .A2(n_194), .B(n_173), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_205), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_211), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_205), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_212), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_219), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_229), .A2(n_196), .B(n_194), .C(n_173), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_206), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_206), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_206), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_233), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_200), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_212), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_200), .A2(n_194), .B(n_186), .C(n_175), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_223), .B(n_177), .Y(n_260) );
CKINVDCx11_ASAP7_75t_R g261 ( .A(n_212), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_212), .B(n_144), .Y(n_262) );
AND3x1_ASAP7_75t_SL g263 ( .A(n_231), .B(n_115), .C(n_117), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_233), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_260), .A2(n_232), .B1(n_213), .B2(n_225), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_251), .A2(n_209), .B(n_204), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_249), .B(n_212), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_243), .Y(n_268) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_259), .A2(n_169), .A3(n_171), .B(n_168), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_234), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_234), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_241), .A2(n_214), .B(n_225), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_234), .A2(n_210), .B(n_209), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_SL g274 ( .A1(n_246), .A2(n_232), .B(n_220), .C(n_219), .Y(n_274) );
OAI21x1_ASAP7_75t_SL g275 ( .A1(n_246), .A2(n_210), .B(n_220), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_264), .B(n_207), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_246), .A2(n_222), .B(n_215), .Y(n_277) );
NOR2xp33_ASAP7_75t_R g278 ( .A(n_261), .B(n_136), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_241), .A2(n_225), .B(n_228), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_243), .Y(n_281) );
OAI221xp5_ASAP7_75t_L g282 ( .A1(n_262), .A2(n_202), .B1(n_227), .B2(n_223), .C(n_131), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_248), .Y(n_283) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_244), .A2(n_124), .B(n_135), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_248), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_244), .A2(n_228), .B(n_222), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_264), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_236), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_274), .A2(n_254), .B(n_253), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g290 ( .A1(n_278), .A2(n_236), .B1(n_249), .B2(n_262), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_288), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_283), .A2(n_254), .B(n_253), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_283), .A2(n_254), .B(n_253), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_282), .A2(n_256), .B1(n_238), .B2(n_239), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_288), .B(n_258), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_270), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_282), .A2(n_260), .B1(n_235), .B2(n_258), .C(n_132), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_265), .A2(n_266), .B(n_271), .C(n_285), .Y(n_299) );
AOI221xp5_ASAP7_75t_SL g300 ( .A1(n_265), .A2(n_235), .B1(n_238), .B2(n_239), .C(n_256), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_283), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_270), .A2(n_237), .B1(n_264), .B2(n_257), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_271), .Y(n_303) );
OAI22xp5_ASAP7_75t_SL g304 ( .A1(n_276), .A2(n_201), .B1(n_263), .B2(n_139), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_280), .A2(n_257), .B(n_255), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_267), .A2(n_131), .B1(n_257), .B2(n_137), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_280), .A2(n_255), .B(n_252), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
CKINVDCx14_ASAP7_75t_R g310 ( .A(n_267), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_291), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_291), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_301), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_301), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_297), .B(n_285), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_303), .B(n_284), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_299), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
NAND2x1_ASAP7_75t_L g320 ( .A(n_305), .B(n_287), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_296), .B(n_269), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_305), .Y(n_322) );
INVx4_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_310), .B(n_284), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_309), .B(n_268), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_299), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_295), .A2(n_237), .B1(n_287), .B2(n_242), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
NOR2x1_ASAP7_75t_L g331 ( .A(n_302), .B(n_284), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_300), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_269), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_289), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_310), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_292), .B(n_269), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_313), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_315), .Y(n_339) );
AOI21x1_ASAP7_75t_L g340 ( .A1(n_335), .A2(n_284), .B(n_272), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_324), .A2(n_307), .B(n_298), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_321), .B(n_307), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_313), .B(n_269), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_315), .B(n_290), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_337), .A2(n_304), .B(n_117), .C(n_145), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_336), .A2(n_126), .B1(n_326), .B2(n_317), .C(n_333), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_313), .B(n_269), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_324), .B(n_287), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_314), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_311), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_269), .Y(n_352) );
INVx5_ASAP7_75t_SL g353 ( .A(n_325), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_312), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_316), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_284), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_334), .B(n_272), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_337), .B(n_263), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_323), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_334), .B(n_116), .Y(n_362) );
AND4x1_ASAP7_75t_L g363 ( .A(n_331), .B(n_147), .C(n_135), .D(n_124), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_317), .B(n_272), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_318), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_323), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
INVx5_ASAP7_75t_L g368 ( .A(n_323), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
OAI33xp33_ASAP7_75t_L g370 ( .A1(n_326), .A2(n_123), .A3(n_147), .B1(n_113), .B2(n_112), .B3(n_143), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_322), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_327), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_318), .B(n_268), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_328), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_333), .B(n_129), .Y(n_376) );
NOR3xp33_ASAP7_75t_SL g377 ( .A(n_329), .B(n_140), .C(n_118), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_331), .A2(n_268), .B1(n_281), .B2(n_242), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_333), .A2(n_325), .B1(n_323), .B2(n_318), .Y(n_380) );
NAND2xp33_ASAP7_75t_SL g381 ( .A(n_320), .B(n_245), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_339), .B(n_333), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_357), .B(n_333), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_358), .B(n_333), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_352), .B(n_319), .Y(n_385) );
OR2x6_ASAP7_75t_L g386 ( .A(n_366), .B(n_332), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_330), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_354), .B(n_319), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_352), .B(n_319), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_362), .B(n_332), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_362), .B(n_375), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_344), .B(n_330), .Y(n_392) );
INVx3_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_344), .B(n_335), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_378), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_342), .A2(n_325), .B1(n_141), .B2(n_116), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_116), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_348), .B(n_325), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_366), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_360), .B(n_141), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_343), .B(n_320), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_343), .B(n_266), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_355), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_359), .B(n_108), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_359), .B(n_155), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_155), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_369), .B(n_128), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_373), .B(n_130), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_364), .B(n_155), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_345), .A3(n_379), .B(n_361), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_373), .B(n_134), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_365), .B(n_142), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_371), .B(n_3), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_365), .B(n_155), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_346), .A2(n_363), .B1(n_347), .B2(n_377), .C(n_376), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_368), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_372), .B(n_4), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_350), .Y(n_419) );
AND2x4_ASAP7_75t_SL g420 ( .A(n_361), .B(n_281), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_350), .Y(n_421) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_361), .B(n_252), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_338), .B(n_155), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_338), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_349), .B(n_155), .Y(n_425) );
NOR2x1_ASAP7_75t_SL g426 ( .A(n_368), .B(n_245), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_367), .B(n_166), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_370), .A2(n_163), .B1(n_275), .B2(n_148), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_349), .B(n_155), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_340), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_368), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_349), .B(n_279), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_349), .B(n_279), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_351), .B(n_5), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_340), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_380), .B(n_279), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_351), .B(n_6), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_353), .B(n_286), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_374), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_353), .B(n_6), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_341), .B(n_7), .Y(n_442) );
NOR2xp33_ASAP7_75t_R g443 ( .A(n_368), .B(n_7), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_368), .B(n_118), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_353), .B(n_286), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_374), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_353), .B(n_8), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_356), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_399), .B(n_356), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_399), .B(n_341), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_405), .B(n_8), .Y(n_451) );
NAND2x1_ASAP7_75t_L g452 ( .A(n_400), .B(n_381), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_405), .B(n_9), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_385), .B(n_9), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_404), .B(n_10), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_395), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_400), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_397), .B(n_10), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_385), .B(n_11), .Y(n_459) );
NAND2x1_ASAP7_75t_L g460 ( .A(n_393), .B(n_275), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_387), .B(n_11), .Y(n_461) );
NOR2xp67_ASAP7_75t_SL g462 ( .A(n_417), .B(n_245), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_431), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_416), .A2(n_281), .B1(n_247), .B2(n_245), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_387), .B(n_391), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_431), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_418), .A2(n_442), .B1(n_401), .B2(n_402), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_417), .B(n_245), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_386), .B(n_12), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_434), .B(n_13), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_397), .B(n_14), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_393), .A2(n_120), .B1(n_146), .B2(n_149), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_443), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_392), .B(n_14), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_388), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_389), .B(n_15), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_391), .B(n_15), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_411), .B(n_393), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_389), .B(n_16), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_384), .B(n_17), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_392), .B(n_17), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_384), .B(n_19), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_448), .Y(n_484) );
NOR3xp33_ASAP7_75t_L g485 ( .A(n_437), .B(n_127), .C(n_170), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_448), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_394), .B(n_20), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_398), .Y(n_488) );
NOR2xp33_ASAP7_75t_SL g489 ( .A(n_417), .B(n_245), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_413), .B(n_21), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_411), .B(n_120), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_398), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_402), .B(n_21), .Y(n_493) );
NAND4xp25_ASAP7_75t_SL g494 ( .A(n_440), .B(n_22), .C(n_23), .D(n_24), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_394), .B(n_22), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_390), .B(n_24), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_413), .B(n_25), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_382), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_393), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_419), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_408), .B(n_25), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_386), .B(n_26), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_406), .B(n_27), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_390), .B(n_286), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_419), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_424), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_421), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_421), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_446), .B(n_30), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_408), .B(n_166), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_439), .B(n_168), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_406), .B(n_170), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_439), .B(n_32), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_409), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_403), .B(n_252), .Y(n_515) );
AND4x1_ASAP7_75t_L g516 ( .A(n_396), .B(n_273), .C(n_277), .D(n_152), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_409), .B(n_146), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_403), .B(n_252), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_446), .B(n_34), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_383), .B(n_439), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_420), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_415), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_424), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_441), .B(n_36), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_412), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_424), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_412), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_441), .B(n_37), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_430), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_383), .B(n_149), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_441), .B(n_38), .Y(n_531) );
OAI221xp5_ASAP7_75t_SL g532 ( .A1(n_467), .A2(n_447), .B1(n_440), .B2(n_386), .C(n_414), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_456), .Y(n_533) );
OAI322xp33_ASAP7_75t_L g534 ( .A1(n_479), .A2(n_447), .A3(n_430), .B1(n_435), .B2(n_427), .C1(n_407), .C2(n_410), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_469), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_465), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_491), .A2(n_444), .B(n_425), .C(n_429), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_484), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_476), .B(n_415), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_486), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_500), .B(n_435), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_488), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_491), .A2(n_429), .B1(n_425), .B2(n_433), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_479), .B(n_422), .Y(n_544) );
OAI22xp33_ASAP7_75t_SL g545 ( .A1(n_474), .A2(n_386), .B1(n_422), .B2(n_410), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_457), .B(n_420), .Y(n_546) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_452), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_521), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_464), .A2(n_432), .B1(n_433), .B2(n_386), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_492), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_463), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_505), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_507), .B(n_508), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_471), .A2(n_427), .B1(n_432), .B2(n_436), .C(n_428), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_466), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_498), .B(n_436), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_520), .Y(n_557) );
OAI31xp33_ASAP7_75t_L g558 ( .A1(n_464), .A2(n_420), .A3(n_438), .B(n_445), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_470), .A2(n_445), .B1(n_438), .B2(n_423), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_522), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_487), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_470), .A2(n_423), .B1(n_407), .B2(n_152), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_455), .B(n_426), .Y(n_563) );
OAI32xp33_ASAP7_75t_L g564 ( .A1(n_468), .A2(n_426), .A3(n_240), .B1(n_255), .B2(n_250), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_487), .Y(n_565) );
OAI21xp33_ASAP7_75t_L g566 ( .A1(n_470), .A2(n_277), .B(n_273), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_529), .B(n_163), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_450), .B(n_40), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_522), .B(n_255), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_485), .B(n_154), .C(n_243), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_495), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_499), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_449), .B(n_41), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_506), .Y(n_574) );
XNOR2x2_ASAP7_75t_L g575 ( .A(n_495), .B(n_496), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_506), .Y(n_576) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_494), .A2(n_247), .B(n_245), .C(n_240), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_502), .B(n_247), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_514), .B(n_163), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_525), .B(n_163), .Y(n_580) );
AOI21xp33_ASAP7_75t_L g581 ( .A1(n_493), .A2(n_42), .B(n_43), .Y(n_581) );
AOI322xp5_ASAP7_75t_L g582 ( .A1(n_496), .A2(n_250), .A3(n_218), .B1(n_217), .B2(n_226), .C1(n_221), .C2(n_207), .Y(n_582) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_485), .B(n_247), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_481), .Y(n_584) );
AND2x2_ASAP7_75t_SL g585 ( .A(n_502), .B(n_247), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_502), .A2(n_240), .B1(n_247), .B2(n_154), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_504), .B(n_45), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_471), .A2(n_154), .B1(n_221), .B2(n_226), .C(n_218), .Y(n_588) );
INVxp33_ASAP7_75t_L g589 ( .A(n_462), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_483), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_475), .A2(n_154), .B1(n_217), .B2(n_215), .C(n_174), .Y(n_591) );
AOI32xp33_ASAP7_75t_L g592 ( .A1(n_454), .A2(n_230), .A3(n_48), .B1(n_51), .B2(n_52), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_499), .A2(n_247), .B(n_154), .C(n_243), .Y(n_593) );
BUFx3_ASAP7_75t_L g594 ( .A(n_468), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_459), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g596 ( .A1(n_482), .A2(n_187), .B(n_181), .C(n_188), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_504), .B(n_46), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_461), .A2(n_59), .B1(n_60), .B2(n_61), .C1(n_62), .C2(n_63), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_529), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_527), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_523), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_523), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_478), .B(n_243), .C(n_183), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_477), .Y(n_604) );
NOR4xp25_ASAP7_75t_L g605 ( .A(n_451), .B(n_64), .C(n_65), .D(n_69), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_480), .A2(n_163), .B1(n_243), .B2(n_183), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_526), .B(n_70), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_526), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_453), .A2(n_174), .B1(n_183), .B2(n_187), .C(n_181), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_532), .A2(n_497), .B1(n_490), .B2(n_458), .C(n_472), .Y(n_610) );
NOR2xp33_ASAP7_75t_SL g611 ( .A(n_585), .B(n_489), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_553), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_604), .A2(n_460), .B1(n_503), .B2(n_530), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_557), .B(n_515), .Y(n_614) );
OAI22xp33_ASAP7_75t_SL g615 ( .A1(n_547), .A2(n_501), .B1(n_517), .B2(n_518), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_555), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_556), .B(n_511), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_556), .B(n_512), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_548), .B(n_531), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_553), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_595), .B(n_516), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_534), .A2(n_473), .B1(n_510), .B2(n_509), .C(n_519), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_536), .B(n_531), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_533), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_561), .B(n_511), .Y(n_625) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_558), .A2(n_524), .B1(n_513), .B2(n_528), .C(n_243), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_535), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_572), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_542), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_560), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_550), .Y(n_631) );
OAI322xp33_ASAP7_75t_L g632 ( .A1(n_575), .A2(n_524), .A3(n_513), .B1(n_183), .B2(n_174), .C1(n_189), .C2(n_179), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_594), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_565), .B(n_71), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_552), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_538), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_541), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_563), .A2(n_183), .B(n_174), .C(n_77), .Y(n_640) );
OAI222xp33_ASAP7_75t_L g641 ( .A1(n_543), .A2(n_72), .B1(n_76), .B2(n_78), .C1(n_79), .C2(n_80), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_541), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_600), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_599), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_571), .B(n_81), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_559), .A2(n_183), .B1(n_174), .B2(n_188), .Y(n_646) );
NAND3xp33_ASAP7_75t_SL g647 ( .A(n_577), .B(n_230), .C(n_84), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_544), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_545), .A2(n_189), .B(n_188), .Y(n_649) );
NAND2xp33_ASAP7_75t_SL g650 ( .A(n_589), .B(n_183), .Y(n_650) );
INVxp33_ASAP7_75t_L g651 ( .A(n_546), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_568), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_551), .B(n_82), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_549), .B(n_174), .C(n_189), .Y(n_654) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_570), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_539), .Y(n_656) );
INVx2_ASAP7_75t_SL g657 ( .A(n_569), .Y(n_657) );
AOI31xp33_ASAP7_75t_L g658 ( .A1(n_578), .A2(n_89), .A3(n_91), .B(n_92), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_584), .B(n_95), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_537), .A2(n_97), .B(n_98), .C(n_99), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_628), .Y(n_661) );
NAND2x1_ASAP7_75t_L g662 ( .A(n_612), .B(n_601), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g663 ( .A1(n_610), .A2(n_592), .B(n_554), .C(n_590), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_616), .B(n_598), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_611), .A2(n_564), .B(n_586), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_633), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_648), .A2(n_566), .B(n_582), .C(n_581), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_655), .B(n_581), .C(n_586), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_615), .A2(n_596), .B(n_605), .C(n_593), .Y(n_669) );
XOR2x2_ASAP7_75t_L g670 ( .A(n_621), .B(n_562), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_621), .A2(n_573), .B1(n_597), .B2(n_603), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_639), .B(n_608), .Y(n_672) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_637), .B(n_602), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_630), .Y(n_674) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_647), .B(n_587), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_637), .B(n_576), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_620), .Y(n_677) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_630), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_642), .B(n_574), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_613), .A2(n_588), .B1(n_591), .B2(n_609), .C(n_580), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_651), .A2(n_607), .B(n_579), .C(n_567), .Y(n_681) );
AO22x1_ASAP7_75t_L g682 ( .A1(n_648), .A2(n_607), .B1(n_567), .B2(n_606), .Y(n_682) );
INVx2_ASAP7_75t_SL g683 ( .A(n_619), .Y(n_683) );
AOI221xp5_ASAP7_75t_SL g684 ( .A1(n_632), .A2(n_101), .B1(n_103), .B2(n_104), .C(n_105), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_652), .Y(n_685) );
OAI32xp33_ASAP7_75t_L g686 ( .A1(n_618), .A2(n_106), .A3(n_179), .B1(n_228), .B2(n_191), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_655), .A2(n_179), .B1(n_228), .B2(n_191), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_644), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_662), .A2(n_658), .B(n_650), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_663), .A2(n_656), .B1(n_629), .B2(n_631), .C(n_627), .Y(n_690) );
AOI211xp5_ASAP7_75t_SL g691 ( .A1(n_664), .A2(n_641), .B(n_626), .C(n_660), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_674), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_678), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_672), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_669), .A2(n_666), .B(n_667), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_677), .B(n_643), .Y(n_696) );
AOI21xp33_ASAP7_75t_SL g697 ( .A1(n_668), .A2(n_654), .B(n_653), .Y(n_697) );
NOR2xp67_ASAP7_75t_L g698 ( .A(n_673), .B(n_635), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_676), .A2(n_641), .B(n_645), .C(n_634), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_670), .A2(n_657), .B1(n_623), .B2(n_614), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g701 ( .A1(n_685), .A2(n_638), .B1(n_636), .B2(n_624), .C1(n_622), .C2(n_625), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_665), .B(n_646), .C(n_640), .D(n_659), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_695), .B(n_675), .C(n_684), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_690), .B(n_661), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_689), .A2(n_672), .B(n_679), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_692), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_698), .B(n_688), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_693), .B(n_679), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_692), .B(n_680), .C(n_682), .Y(n_709) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_706), .Y(n_710) );
OR3x2_ASAP7_75t_L g711 ( .A(n_708), .B(n_702), .C(n_703), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_709), .A2(n_701), .B(n_691), .C(n_697), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_704), .B(n_699), .C(n_694), .Y(n_713) );
AOI322xp5_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_707), .A3(n_700), .B1(n_683), .B2(n_696), .C1(n_671), .C2(n_680), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_712), .B(n_705), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_710), .B(n_687), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_715), .A2(n_711), .B1(n_617), .B2(n_649), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_716), .A2(n_681), .B1(n_686), .B2(n_191), .Y(n_718) );
AOI22xp33_ASAP7_75t_R g719 ( .A1(n_717), .A2(n_714), .B1(n_180), .B2(n_182), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_180), .B1(n_182), .B2(n_715), .C1(n_712), .C2(n_717), .Y(n_721) );
NOR2x1_ASAP7_75t_R g722 ( .A(n_719), .B(n_182), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_722), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_721), .B(n_180), .Y(n_724) );
endmodule