module real_jpeg_23759_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_1),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_31),
.B1(n_36),
.B2(n_39),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_1),
.A2(n_31),
.B1(n_50),
.B2(n_54),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_31),
.B1(n_62),
.B2(n_98),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_50),
.B1(n_54),
.B2(n_58),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_2),
.A2(n_36),
.B1(n_39),
.B2(n_58),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_58),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_4),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_42),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_4),
.A2(n_42),
.B1(n_50),
.B2(n_54),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_4),
.A2(n_53),
.B(n_59),
.C(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_4),
.B(n_49),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_42),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_54),
.B(n_77),
.C(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_4),
.B(n_22),
.C(n_38),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_4),
.B(n_83),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_11),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_4),
.B(n_40),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_20)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_11),
.Y(n_138)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_11),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_127),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_126),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_112),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_112),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_87),
.B2(n_111),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_45),
.B1(n_85),
.B2(n_86),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_18),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_32),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_24),
.B(n_26),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_20),
.A2(n_107),
.B(n_110),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_21),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_22),
.B(n_184),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_24),
.B(n_30),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_24),
.B(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_24),
.A2(n_125),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_24),
.B(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_27),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_27),
.B(n_169),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_43),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_33),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_34),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_34),
.B(n_44),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_35)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_36),
.A2(n_39),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_36),
.B(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_39),
.A2(n_42),
.B(n_78),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_40),
.B(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_42),
.A2(n_52),
.B(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_43),
.B(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_68),
.C(n_73),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_46),
.A2(n_47),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_60),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_54),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_65),
.Y(n_100)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_71),
.B(n_72),
.Y(n_140)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_81),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_80),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_82),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_103),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_95),
.B1(n_101),
.B2(n_102),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_94),
.B(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_110),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_119),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_114),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_119),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_123),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_147),
.B(n_211),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_144),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_129),
.B(n_144),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_139),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_130),
.B(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_132),
.B(n_139),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_133),
.A2(n_135),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_133),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_135),
.Y(n_203)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_206),
.B(n_210),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_193),
.B(n_205),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_173),
.B(n_192),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_151),
.B(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_154),
.B1(n_155),
.B2(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_172),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_163),
.C(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_181),
.B(n_191),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_187),
.B(n_190),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_195),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_207),
.B(n_208),
.Y(n_210)
);


endmodule