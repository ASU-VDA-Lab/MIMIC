module fake_jpeg_5943_n_252 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_30),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

NOR2xp67_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_51),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_47),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_31),
.C(n_32),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_49),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_36),
.B1(n_32),
.B2(n_30),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_71),
.B1(n_49),
.B2(n_36),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_50),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_36),
.B1(n_30),
.B2(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_34),
.B1(n_51),
.B2(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_36),
.B1(n_30),
.B2(n_31),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_88),
.B1(n_58),
.B2(n_14),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_75),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_77),
.B1(n_68),
.B2(n_70),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_47),
.B1(n_30),
.B2(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_63),
.B1(n_62),
.B2(n_34),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_68),
.B1(n_54),
.B2(n_55),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_97),
.B1(n_84),
.B2(n_82),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_80),
.C(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_106),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_80),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_73),
.C(n_83),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_114),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_75),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_34),
.B1(n_50),
.B2(n_17),
.Y(n_152)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_71),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_119),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_88),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_103),
.B1(n_108),
.B2(n_53),
.Y(n_139)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_128),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_99),
.B(n_110),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_103),
.B(n_61),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_86),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_76),
.B1(n_81),
.B2(n_62),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_94),
.B1(n_100),
.B2(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_150),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_14),
.B1(n_25),
.B2(n_85),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_34),
.B1(n_29),
.B2(n_22),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_17),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_153),
.B1(n_120),
.B2(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_120),
.B1(n_114),
.B2(n_128),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_123),
.B(n_119),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_160),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_112),
.C(n_111),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_129),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_145),
.B(n_119),
.C(n_115),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_131),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_50),
.C(n_29),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_167),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_50),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_152),
.B1(n_134),
.B2(n_147),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_172),
.B1(n_141),
.B2(n_144),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_50),
.C(n_29),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_146),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_22),
.B1(n_16),
.B2(n_18),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_155),
.B1(n_167),
.B2(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_190),
.B(n_22),
.Y(n_205)
);

NAND2xp67_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_143),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_169),
.B1(n_172),
.B2(n_149),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_141),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_189),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_174),
.B(n_162),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_198),
.B(n_202),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_161),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_13),
.C(n_18),
.Y(n_213)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_170),
.B(n_163),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_206),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_23),
.B(n_7),
.Y(n_209)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

NAND4xp25_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_183),
.C(n_185),
.D(n_180),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_214),
.B(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_212),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_1),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_13),
.C(n_1),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_6),
.C(n_12),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_192),
.B1(n_202),
.B2(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_13),
.C(n_1),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_5),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_215),
.A2(n_199),
.B1(n_204),
.B2(n_200),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_222),
.C(n_209),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_199),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_221),
.B(n_224),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_5),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_210),
.A2(n_5),
.B1(n_12),
.B2(n_10),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_0),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_218),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_233),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_234),
.B(n_235),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_228),
.B(n_8),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_2),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_220),
.B(n_8),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_227),
.B(n_224),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_242),
.C(n_10),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_9),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_23),
.B(n_9),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_237),
.B(n_3),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_3),
.B1(n_4),
.B2(n_245),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_3),
.B(n_4),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_250),
.Y(n_252)
);


endmodule