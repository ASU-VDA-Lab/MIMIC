module fake_jpeg_18009_n_289 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp67_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_25),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_20),
.B1(n_31),
.B2(n_30),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_59),
.B1(n_62),
.B2(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_68),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_60),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_27),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_33),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_35),
.B(n_43),
.Y(n_87)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_31),
.B1(n_24),
.B2(n_25),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_70),
.B(n_101),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_85),
.B1(n_98),
.B2(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_79),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_95),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_32),
.A3(n_33),
.B1(n_69),
.B2(n_47),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_90),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_94),
.Y(n_119)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_26),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_99),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_39),
.B1(n_43),
.B2(n_31),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_26),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_26),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_22),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_63),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_118),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_1),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_23),
.Y(n_110)
);

NAND2x1p5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_43),
.B1(n_25),
.B2(n_24),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_78),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_30),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_113),
.B(n_121),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_65),
.B1(n_35),
.B2(n_46),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_126),
.B1(n_76),
.B2(n_42),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_34),
.B1(n_30),
.B2(n_24),
.Y(n_116)
);

OAI21x1_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_122),
.B(n_125),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_71),
.B(n_34),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_34),
.B1(n_77),
.B2(n_92),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_84),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_70),
.B(n_46),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_69),
.B1(n_47),
.B2(n_42),
.Y(n_126)
);

OR2x6_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_47),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_71),
.A2(n_33),
.A3(n_32),
.B1(n_22),
.B2(n_37),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_42),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_82),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_140),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_75),
.B1(n_99),
.B2(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_151),
.B1(n_160),
.B2(n_125),
.Y(n_175)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_89),
.B1(n_100),
.B2(n_80),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_145),
.B(n_130),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_149),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_100),
.C(n_22),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_111),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_95),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_81),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_81),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_158),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_113),
.B(n_96),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_159),
.B(n_138),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_167),
.B(n_168),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_109),
.B1(n_118),
.B2(n_119),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_170),
.B1(n_151),
.B2(n_150),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_127),
.B(n_129),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_110),
.B(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_138),
.B1(n_148),
.B2(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_169),
.A2(n_188),
.B1(n_8),
.B2(n_9),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_127),
.B1(n_115),
.B2(n_106),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_125),
.B(n_110),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_175),
.B(n_189),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_147),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_6),
.B(n_7),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_108),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_135),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_108),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_120),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_139),
.A2(n_120),
.B1(n_84),
.B2(n_76),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_67),
.B(n_55),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_190),
.B(n_169),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_144),
.B1(n_139),
.B2(n_160),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_191),
.A2(n_193),
.B1(n_200),
.B2(n_163),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_201),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_197),
.B(n_212),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_149),
.C(n_76),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_209),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_33),
.CI(n_5),
.CON(n_201),
.SN(n_201)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_205),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_210),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_177),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_3),
.B(n_5),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_8),
.B(n_9),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_6),
.C(n_7),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_163),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_161),
.A2(n_186),
.B1(n_185),
.B2(n_174),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_168),
.B1(n_178),
.B2(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_228),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_221),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_179),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_224),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_190),
.B(n_167),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_178),
.B1(n_174),
.B2(n_186),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_185),
.B1(n_182),
.B2(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_180),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_181),
.B1(n_165),
.B2(n_188),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_203),
.B1(n_196),
.B2(n_195),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_195),
.A2(n_189),
.B1(n_164),
.B2(n_10),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_233),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_231),
.A2(n_208),
.B(n_210),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_199),
.B(n_194),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_243),
.B(n_246),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_231),
.B(n_222),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_210),
.B1(n_199),
.B2(n_194),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_223),
.B(n_232),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_209),
.C(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_247),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_201),
.A3(n_198),
.B(n_12),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_225),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_201),
.C(n_11),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_260),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_221),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_234),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_229),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_226),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_248),
.Y(n_263)
);

NAND4xp25_ASAP7_75t_SL g261 ( 
.A(n_259),
.B(n_248),
.C(n_240),
.D(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_265),
.Y(n_274)
);

AOI31xp67_ASAP7_75t_SL g264 ( 
.A1(n_256),
.A2(n_238),
.A3(n_236),
.B(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_268),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_253),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_218),
.B1(n_11),
.B2(n_12),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_14),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_249),
.B(n_251),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_260),
.B1(n_261),
.B2(n_270),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_254),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_272),
.B(n_14),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_266),
.C(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_277),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_282),
.B(n_275),
.C(n_276),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_15),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_15),
.B(n_16),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_278),
.B(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_286),
.B(n_287),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_283),
.Y(n_289)
);


endmodule