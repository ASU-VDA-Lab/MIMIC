module real_aes_7267_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g507 ( .A(n_0), .Y(n_507) );
AOI22xp5_ASAP7_75t_SL g689 ( .A1(n_1), .A2(n_191), .B1(n_347), .B2(n_495), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_2), .Y(n_708) );
XOR2x2_ASAP7_75t_L g710 ( .A(n_2), .B(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_3), .A2(n_14), .B1(n_385), .B2(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g331 ( .A(n_4), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_5), .A2(n_101), .B1(n_381), .B2(n_382), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_6), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g726 ( .A1(n_7), .A2(n_33), .B1(n_184), .B2(n_316), .C1(n_546), .C2(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g490 ( .A(n_8), .Y(n_490) );
INVx1_ASAP7_75t_L g479 ( .A(n_9), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_10), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_11), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_12), .A2(n_66), .B1(n_719), .B2(n_720), .Y(n_718) );
AOI222xp33_ASAP7_75t_L g608 ( .A1(n_13), .A2(n_112), .B1(n_179), .B2(n_316), .C1(n_381), .C2(n_431), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_15), .A2(n_98), .B1(n_276), .B2(n_280), .C(n_285), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_16), .A2(n_64), .B1(n_647), .B2(n_648), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_17), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_18), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_19), .A2(n_146), .B1(n_555), .B2(n_581), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_20), .Y(n_693) );
INVx1_ASAP7_75t_L g500 ( .A(n_21), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_22), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_23), .Y(n_370) );
AO22x2_ASAP7_75t_L g257 ( .A1(n_24), .A2(n_77), .B1(n_249), .B2(n_254), .Y(n_257) );
INVx1_ASAP7_75t_L g678 ( .A(n_24), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_25), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_26), .A2(n_166), .B1(n_393), .B2(n_400), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g345 ( .A1(n_27), .A2(n_221), .B1(n_346), .B2(n_347), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_28), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_29), .A2(n_141), .B1(n_538), .B2(n_638), .Y(n_637) );
XOR2xp5_ASAP7_75t_L g681 ( .A(n_30), .B(n_682), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_31), .A2(n_139), .B1(n_281), .B2(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_32), .A2(n_175), .B1(n_320), .B2(n_386), .Y(n_697) );
INVx1_ASAP7_75t_L g497 ( .A(n_34), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_35), .B(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_36), .A2(n_39), .B1(n_300), .B2(n_535), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_37), .A2(n_406), .B1(n_441), .B2(n_442), .Y(n_405) );
INVx1_ASAP7_75t_L g441 ( .A(n_37), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_38), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_40), .A2(n_152), .B1(n_387), .B2(n_621), .Y(n_620) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_41), .A2(n_82), .B1(n_249), .B2(n_250), .Y(n_259) );
INVx1_ASAP7_75t_L g679 ( .A(n_41), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_42), .A2(n_118), .B1(n_326), .B2(n_365), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_43), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_44), .A2(n_140), .B1(n_346), .B2(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_45), .A2(n_213), .B1(n_297), .B2(n_300), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_46), .A2(n_144), .B1(n_281), .B2(n_420), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_47), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_48), .A2(n_81), .B1(n_291), .B2(n_413), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_49), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_50), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_51), .Y(n_409) );
AOI22xp5_ASAP7_75t_SL g686 ( .A1(n_52), .A2(n_142), .B1(n_579), .B2(n_687), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_53), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_54), .A2(n_87), .B1(n_296), .B2(n_300), .C(n_302), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_55), .A2(n_239), .B1(n_240), .B2(n_328), .Y(n_238) );
INVx1_ASAP7_75t_L g328 ( .A(n_55), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_56), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_57), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_58), .A2(n_217), .B1(n_339), .B2(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_59), .A2(n_131), .B1(n_364), .B2(n_386), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_60), .A2(n_162), .B1(n_504), .B2(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_61), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_62), .A2(n_172), .B1(n_244), .B2(n_414), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_63), .A2(n_168), .B1(n_395), .B2(n_583), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_65), .Y(n_353) );
AOI22xp5_ASAP7_75t_SL g685 ( .A1(n_67), .A2(n_124), .B1(n_260), .B2(n_335), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_68), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_69), .A2(n_183), .B1(n_297), .B2(n_301), .Y(n_698) );
AO22x2_ASAP7_75t_L g563 ( .A1(n_70), .A2(n_564), .B1(n_587), .B2(n_588), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_70), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_71), .A2(n_189), .B1(n_414), .B2(n_581), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_72), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_73), .Y(n_531) );
AOI211xp5_ASAP7_75t_L g528 ( .A1(n_74), .A2(n_529), .B(n_530), .C(n_540), .Y(n_528) );
AOI22xp5_ASAP7_75t_SL g334 ( .A1(n_75), .A2(n_129), .B1(n_281), .B2(n_335), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_76), .A2(n_130), .B1(n_344), .B2(n_393), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_78), .Y(n_461) );
AOI222xp33_ASAP7_75t_L g315 ( .A1(n_79), .A2(n_100), .B1(n_120), .B2(n_316), .C1(n_318), .C2(n_324), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_80), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_83), .A2(n_170), .B1(n_268), .B2(n_292), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_84), .Y(n_432) );
INVx1_ASAP7_75t_L g229 ( .A(n_85), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_86), .A2(n_169), .B1(n_395), .B2(n_396), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_88), .A2(n_119), .B1(n_280), .B2(n_400), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_89), .B(n_517), .Y(n_516) );
AOI22xp5_ASAP7_75t_SL g342 ( .A1(n_90), .A2(n_192), .B1(n_343), .B2(n_344), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_91), .A2(n_158), .B1(n_363), .B2(n_364), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_92), .A2(n_171), .B1(n_551), .B2(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g226 ( .A(n_93), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_94), .A2(n_145), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_95), .A2(n_128), .B1(n_320), .B2(n_326), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_96), .A2(n_223), .B(n_231), .C(n_680), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_97), .A2(n_195), .B1(n_292), .B2(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g455 ( .A(n_99), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_102), .A2(n_196), .B1(n_267), .B2(n_586), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_103), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_104), .A2(n_149), .B1(n_278), .B2(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g509 ( .A(n_105), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_106), .A2(n_208), .B1(n_657), .B2(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g521 ( .A(n_107), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_108), .A2(n_115), .B1(n_386), .B2(n_543), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_109), .Y(n_428) );
INVx1_ASAP7_75t_L g289 ( .A(n_110), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_111), .A2(n_486), .B1(n_522), .B2(n_523), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_111), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_113), .A2(n_198), .B1(n_653), .B2(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g480 ( .A(n_114), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_116), .A2(n_190), .B1(n_292), .B2(n_401), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_117), .A2(n_218), .B1(n_723), .B2(n_724), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_121), .A2(n_165), .B1(n_243), .B2(n_260), .C(n_265), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_122), .A2(n_155), .B1(n_365), .B2(n_381), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_123), .A2(n_177), .B1(n_537), .B2(n_538), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_125), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_126), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g230 ( .A(n_127), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_132), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_133), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_134), .A2(n_173), .B1(n_291), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_135), .A2(n_199), .B1(n_502), .B2(n_504), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_136), .Y(n_526) );
AND2x6_ASAP7_75t_L g225 ( .A(n_137), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_137), .Y(n_672) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_138), .A2(n_187), .B1(n_249), .B2(n_250), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_143), .A2(n_205), .B1(n_339), .B2(n_396), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_147), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_148), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_150), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_151), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_153), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_154), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_156), .A2(n_209), .B1(n_585), .B2(n_586), .Y(n_584) );
AO22x1_ASAP7_75t_L g265 ( .A1(n_157), .A2(n_185), .B1(n_266), .B2(n_270), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_159), .A2(n_202), .B1(n_344), .B2(n_393), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_160), .Y(n_628) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_161), .A2(n_201), .B1(n_249), .B2(n_254), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_163), .A2(n_203), .B1(n_514), .B2(n_546), .Y(n_573) );
INVx1_ASAP7_75t_L g562 ( .A(n_164), .Y(n_562) );
INVx1_ASAP7_75t_L g452 ( .A(n_167), .Y(n_452) );
INVx1_ASAP7_75t_L g476 ( .A(n_174), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_176), .A2(n_204), .B1(n_260), .B2(n_579), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_178), .B(n_347), .Y(n_466) );
INVx1_ASAP7_75t_L g515 ( .A(n_180), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_181), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_182), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_186), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_187), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_188), .B(n_300), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_193), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_194), .Y(n_569) );
INVx1_ASAP7_75t_L g519 ( .A(n_197), .Y(n_519) );
INVx1_ASAP7_75t_L g286 ( .A(n_200), .Y(n_286) );
INVx1_ASAP7_75t_L g675 ( .A(n_201), .Y(n_675) );
INVx1_ASAP7_75t_L g493 ( .A(n_206), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_207), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_210), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_211), .Y(n_307) );
INVx1_ASAP7_75t_L g249 ( .A(n_212), .Y(n_249) );
INVx1_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_214), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_215), .Y(n_436) );
INVx1_ASAP7_75t_L g512 ( .A(n_216), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_219), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_220), .A2(n_632), .B1(n_661), .B2(n_662), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_220), .Y(n_661) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_226), .Y(n_671) );
OA21x2_ASAP7_75t_L g706 ( .A1(n_227), .A2(n_670), .B(n_707), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_593), .B1(n_665), .B2(n_666), .C(n_667), .Y(n_231) );
INVx1_ASAP7_75t_L g665 ( .A(n_232), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B1(n_446), .B2(n_592), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B1(n_373), .B2(n_445), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_329), .B1(n_371), .B2(n_372), .Y(n_236) );
INVx1_ASAP7_75t_L g371 ( .A(n_237), .Y(n_371) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND4x1_ASAP7_75t_L g241 ( .A(n_242), .B(n_275), .C(n_295), .D(n_315), .Y(n_241) );
INVx1_ASAP7_75t_SL g489 ( .A(n_243), .Y(n_489) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g416 ( .A(n_244), .Y(n_416) );
BUFx3_ASAP7_75t_L g647 ( .A(n_244), .Y(n_647) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g340 ( .A(n_245), .Y(n_340) );
BUFx2_ASAP7_75t_SL g687 ( .A(n_245), .Y(n_687) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
AND2x6_ASAP7_75t_L g262 ( .A(n_246), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g278 ( .A(n_246), .B(n_279), .Y(n_278) );
AND2x6_ASAP7_75t_L g317 ( .A(n_246), .B(n_312), .Y(n_317) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
AND2x2_ASAP7_75t_L g269 ( .A(n_247), .B(n_253), .Y(n_269) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_248), .B(n_253), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_248), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g305 ( .A(n_248), .B(n_257), .Y(n_305) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g254 ( .A(n_251), .Y(n_254) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
INVx1_ASAP7_75t_L g323 ( .A(n_253), .Y(n_323) );
AND2x4_ASAP7_75t_L g268 ( .A(n_255), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g272 ( .A(n_255), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g282 ( .A(n_255), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_255), .B(n_283), .Y(n_477) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
OR2x2_ASAP7_75t_L g264 ( .A(n_256), .B(n_259), .Y(n_264) );
AND2x2_ASAP7_75t_L g279 ( .A(n_256), .B(n_259), .Y(n_279) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g312 ( .A(n_257), .B(n_259), .Y(n_312) );
INVx1_ASAP7_75t_L g306 ( .A(n_258), .Y(n_306) );
AND2x2_ASAP7_75t_L g322 ( .A(n_258), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g294 ( .A(n_259), .Y(n_294) );
INVx1_ASAP7_75t_L g558 ( .A(n_260), .Y(n_558) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx4_ASAP7_75t_L g343 ( .A(n_261), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_261), .A2(n_409), .B1(n_410), .B2(n_411), .C(n_412), .Y(n_408) );
INVx2_ASAP7_75t_SL g492 ( .A(n_261), .Y(n_492) );
INVx4_ASAP7_75t_L g723 ( .A(n_261), .Y(n_723) );
INVx11_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx11_ASAP7_75t_L g397 ( .A(n_262), .Y(n_397) );
AND2x4_ASAP7_75t_L g299 ( .A(n_263), .B(n_269), .Y(n_299) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g359 ( .A(n_264), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_268), .Y(n_346) );
BUFx3_ASAP7_75t_L g420 ( .A(n_268), .Y(n_420) );
INVx2_ASAP7_75t_L g464 ( .A(n_268), .Y(n_464) );
BUFx3_ASAP7_75t_L g583 ( .A(n_268), .Y(n_583) );
AND2x6_ASAP7_75t_L g301 ( .A(n_269), .B(n_279), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_269), .B(n_279), .Y(n_352) );
INVx1_ASAP7_75t_L g360 ( .A(n_269), .Y(n_360) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g410 ( .A(n_271), .Y(n_410) );
BUFx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx3_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
INVx1_ASAP7_75t_L g473 ( .A(n_272), .Y(n_473) );
BUFx3_ASAP7_75t_L g495 ( .A(n_272), .Y(n_495) );
BUFx2_ASAP7_75t_L g553 ( .A(n_272), .Y(n_553) );
BUFx3_ASAP7_75t_L g586 ( .A(n_272), .Y(n_586) );
AND2x2_ASAP7_75t_L g347 ( .A(n_273), .B(n_306), .Y(n_347) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x6_ASAP7_75t_L g293 ( .A(n_274), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g400 ( .A(n_277), .Y(n_400) );
OAI22xp5_ASAP7_75t_SL g467 ( .A1(n_277), .A2(n_340), .B1(n_468), .B2(n_469), .Y(n_467) );
OAI221xp5_ASAP7_75t_SL g496 ( .A1(n_277), .A2(n_497), .B1(n_498), .B2(n_500), .C(n_501), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_277), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_556) );
INVx2_ASAP7_75t_L g655 ( .A(n_277), .Y(n_655) );
INVx6_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx3_ASAP7_75t_L g579 ( .A(n_278), .Y(n_579) );
BUFx3_ASAP7_75t_L g724 ( .A(n_278), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_279), .B(n_283), .Y(n_288) );
AND2x2_ASAP7_75t_L g337 ( .A(n_279), .B(n_283), .Y(n_337) );
BUFx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx3_ASAP7_75t_L g393 ( .A(n_282), .Y(n_393) );
BUFx3_ASAP7_75t_L g659 ( .A(n_282), .Y(n_659) );
BUFx3_ASAP7_75t_L g717 ( .A(n_282), .Y(n_717) );
INVx1_ASAP7_75t_L g314 ( .A(n_284), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B1(n_289), .B2(n_290), .Y(n_285) );
BUFx2_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_288), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_291), .Y(n_290) );
BUFx4f_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
BUFx2_ASAP7_75t_L g581 ( .A(n_292), .Y(n_581) );
INVx6_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g504 ( .A(n_293), .Y(n_504) );
INVx1_ASAP7_75t_L g388 ( .A(n_294), .Y(n_388) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx5_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g535 ( .A(n_298), .Y(n_535) );
INVx2_ASAP7_75t_L g606 ( .A(n_298), .Y(n_606) );
INVx2_ASAP7_75t_L g619 ( .A(n_298), .Y(n_619) );
INVx4_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx4f_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_307), .B2(n_308), .Y(n_302) );
INVx4_ASAP7_75t_L g355 ( .A(n_304), .Y(n_355) );
BUFx3_ASAP7_75t_L g439 ( .A(n_304), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_304), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x4_ASAP7_75t_L g321 ( .A(n_305), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g326 ( .A(n_305), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g387 ( .A(n_305), .B(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_308), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_308), .A2(n_519), .B1(n_520), .B2(n_521), .Y(n_518) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
CKINVDCx16_ASAP7_75t_R g309 ( .A(n_310), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_310), .A2(n_520), .B1(n_575), .B2(n_576), .Y(n_574) );
OR2x6_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g365 ( .A(n_312), .B(n_314), .Y(n_365) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g433 ( .A(n_316), .Y(n_433) );
INVx2_ASAP7_75t_SL g511 ( .A(n_316), .Y(n_511) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx4_ASAP7_75t_L g367 ( .A(n_317), .Y(n_367) );
INVx2_ASAP7_75t_L g379 ( .A(n_317), .Y(n_379) );
INVx2_ASAP7_75t_SL g460 ( .A(n_317), .Y(n_460) );
BUFx3_ASAP7_75t_L g529 ( .A(n_317), .Y(n_529) );
INVx2_ASAP7_75t_L g694 ( .A(n_317), .Y(n_694) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_319), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_458) );
INVx4_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g369 ( .A(n_320), .Y(n_369) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx4f_ASAP7_75t_SL g385 ( .A(n_321), .Y(n_385) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_321), .Y(n_431) );
BUFx2_ASAP7_75t_L g514 ( .A(n_321), .Y(n_514) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_321), .Y(n_543) );
INVx1_ASAP7_75t_L g327 ( .A(n_323), .Y(n_327) );
INVx2_ASAP7_75t_L g435 ( .A(n_324), .Y(n_435) );
BUFx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
BUFx12f_ASAP7_75t_L g381 ( .A(n_326), .Y(n_381) );
INVx1_ASAP7_75t_SL g372 ( .A(n_329), .Y(n_372) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
XNOR2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND3x1_ASAP7_75t_SL g332 ( .A(n_333), .B(n_341), .C(n_348), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_338), .Y(n_333) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx5_ASAP7_75t_L g401 ( .A(n_336), .Y(n_401) );
INVx2_ASAP7_75t_L g414 ( .A(n_336), .Y(n_414) );
BUFx3_ASAP7_75t_L g503 ( .A(n_336), .Y(n_503) );
INVx1_ASAP7_75t_L g555 ( .A(n_336), .Y(n_555) );
INVx8_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g395 ( .A(n_340), .Y(n_395) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
BUFx2_ASAP7_75t_L g660 ( .A(n_344), .Y(n_660) );
INVx4_ASAP7_75t_L g552 ( .A(n_346), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_357), .C(n_366), .Y(n_348) );
OAI22xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_353), .B1(n_354), .B2(n_356), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_350), .A2(n_425), .B1(n_426), .B2(n_428), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_350), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g456 ( .A(n_352), .Y(n_456) );
INVx3_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g520 ( .A(n_355), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_361), .B(n_362), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g427 ( .A(n_359), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_359), .A2(n_452), .B(n_453), .Y(n_451) );
BUFx4f_ASAP7_75t_L g517 ( .A(n_363), .Y(n_517) );
INVx1_ASAP7_75t_SL g539 ( .A(n_364), .Y(n_539) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_SL g382 ( .A(n_365), .Y(n_382) );
BUFx3_ASAP7_75t_L g621 ( .A(n_365), .Y(n_621) );
BUFx2_ASAP7_75t_SL g727 ( .A(n_365), .Y(n_727) );
OAI22xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B1(n_369), .B2(n_370), .Y(n_366) );
INVx1_ASAP7_75t_L g445 ( .A(n_373), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_404), .B1(n_443), .B2(n_444), .Y(n_373) );
INVx3_ASAP7_75t_SL g443 ( .A(n_374), .Y(n_443) );
XOR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_403), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_376), .B(n_390), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_383), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_380), .Y(n_377) );
OAI21xp5_ASAP7_75t_SL g613 ( .A1(n_379), .A2(n_614), .B(n_615), .Y(n_613) );
OAI222xp33_ASAP7_75t_L g640 ( .A1(n_379), .A2(n_430), .B1(n_435), .B2(n_641), .C1(n_642), .C2(n_643), .Y(n_640) );
INVx2_ASAP7_75t_L g547 ( .A(n_381), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_389), .Y(n_383) );
BUFx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g537 ( .A(n_387), .Y(n_537) );
INVx1_ASAP7_75t_L g639 ( .A(n_387), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_398), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx5_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_397), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_SL g585 ( .A(n_397), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
BUFx2_ASAP7_75t_L g650 ( .A(n_401), .Y(n_650) );
INVx3_ASAP7_75t_L g444 ( .A(n_404), .Y(n_444) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_407), .B(n_423), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_415), .Y(n_407) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_417), .B1(n_418), .B2(n_421), .C(n_422), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_429), .C(n_437), .Y(n_423) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g508 ( .A(n_427), .Y(n_508) );
INVx2_ASAP7_75t_L g568 ( .A(n_427), .Y(n_568) );
OAI222xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_433), .B2(n_434), .C1(n_435), .C2(n_436), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g592 ( .A(n_446), .Y(n_592) );
XNOR2xp5_ASAP7_75t_SL g446 ( .A(n_447), .B(n_481), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
XNOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_480), .Y(n_448) );
AND3x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_462), .C(n_470), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .C(n_458), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_456), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
INVx2_ASAP7_75t_L g533 ( .A(n_456), .Y(n_533) );
OA211x2_ASAP7_75t_L g603 ( .A1(n_456), .A2(n_604), .B(n_605), .C(n_607), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
OAI21xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_465), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g648 ( .A(n_464), .Y(n_648) );
INVx2_ASAP7_75t_L g719 ( .A(n_464), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .C(n_478), .Y(n_470) );
INVx1_ASAP7_75t_L g720 ( .A(n_473), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g499 ( .A(n_477), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_524), .B2(n_591), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g523 ( .A(n_486), .Y(n_523) );
AND2x2_ASAP7_75t_SL g486 ( .A(n_487), .B(n_505), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
OAI221xp5_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_490), .B1(n_491), .B2(n_493), .C(n_494), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_489), .A2(n_498), .B1(n_561), .B2(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .C(n_518), .Y(n_505) );
OAI221xp5_ASAP7_75t_SL g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_515), .C(n_516), .Y(n_510) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g591 ( .A(n_524), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_563), .B1(n_589), .B2(n_590), .Y(n_524) );
INVx2_ASAP7_75t_L g589 ( .A(n_525), .Y(n_589) );
XNOR2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_548), .Y(n_527) );
INVx3_ASAP7_75t_L g572 ( .A(n_529), .Y(n_572) );
OAI211xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_534), .C(n_536), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_532), .A2(n_568), .B1(n_635), .B2(n_636), .C(n_637), .Y(n_634) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_544), .B2(n_545), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_556), .C(n_560), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g590 ( .A(n_563), .Y(n_590) );
INVx1_ASAP7_75t_SL g587 ( .A(n_564), .Y(n_587) );
AND2x2_ASAP7_75t_SL g564 ( .A(n_565), .B(n_577), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .C(n_574), .Y(n_565) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B(n_573), .Y(n_570) );
AND4x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .C(n_582), .D(n_584), .Y(n_577) );
INVx1_ASAP7_75t_L g654 ( .A(n_585), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g666 ( .A(n_593), .Y(n_666) );
AOI22xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_631), .B1(n_663), .B2(n_664), .Y(n_593) );
INVx1_ASAP7_75t_L g663 ( .A(n_594), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_610), .B1(n_629), .B2(n_630), .Y(n_594) );
INVx2_ASAP7_75t_SL g629 ( .A(n_595), .Y(n_629) );
XOR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_609), .Y(n_595) );
NAND4xp75_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .C(n_603), .D(n_608), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx4_ASAP7_75t_SL g630 ( .A(n_610), .Y(n_630) );
XOR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_628), .Y(n_610) );
NAND3x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_622), .C(n_625), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .C(n_620), .Y(n_616) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g664 ( .A(n_631), .Y(n_664) );
INVx1_ASAP7_75t_SL g662 ( .A(n_632), .Y(n_662) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_644), .Y(n_632) );
NOR2xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_640), .Y(n_633) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_651), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_652), .B(n_656), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .Y(n_668) );
OR2x2_ASAP7_75t_SL g730 ( .A(n_669), .B(n_674), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_671), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_671), .B(n_703), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g703 ( .A(n_672), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_699), .A3(n_700), .B1(n_704), .B2(n_708), .C1(n_709), .C2(n_728), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND4xp75_ASAP7_75t_SL g684 ( .A(n_685), .B(n_686), .C(n_688), .D(n_691), .Y(n_684) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_696), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_695), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_705), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND4xp75_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .C(n_721), .D(n_726), .Y(n_711) );
AND2x2_ASAP7_75t_SL g712 ( .A(n_713), .B(n_714), .Y(n_712) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
endmodule