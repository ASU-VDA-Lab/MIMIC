module fake_jpeg_4628_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_24),
.B(n_19),
.C(n_28),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_60),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_19),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_20),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_36),
.B1(n_35),
.B2(n_17),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_69),
.B1(n_76),
.B2(n_21),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_82),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_36),
.B1(n_35),
.B2(n_17),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_24),
.B1(n_16),
.B2(n_31),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_56),
.B1(n_22),
.B2(n_52),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_31),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_84),
.B(n_25),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_17),
.B1(n_40),
.B2(n_39),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_28),
.B1(n_22),
.B2(n_16),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_39),
.C(n_20),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_30),
.C(n_58),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_27),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_23),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_46),
.B1(n_42),
.B2(n_47),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_96),
.B1(n_99),
.B2(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_94),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_93),
.A2(n_101),
.B(n_70),
.Y(n_128)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_57),
.B1(n_48),
.B2(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_100),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_31),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_22),
.B1(n_29),
.B2(n_25),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_55),
.B(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_106),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_2),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_66),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_21),
.B1(n_15),
.B2(n_18),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_71),
.B1(n_84),
.B2(n_83),
.Y(n_130)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_116),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_79),
.C(n_70),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_91),
.C(n_55),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_72),
.B1(n_78),
.B2(n_64),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_130),
.B1(n_97),
.B2(n_99),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_117),
.B(n_118),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_83),
.B1(n_78),
.B2(n_64),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_89),
.B1(n_92),
.B2(n_107),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_71),
.B(n_50),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_97),
.B(n_93),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_127),
.B1(n_120),
.B2(n_132),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_111),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_149),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_144),
.B1(n_150),
.B2(n_122),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_92),
.B1(n_106),
.B2(n_105),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_75),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_131),
.C(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_125),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_159),
.C(n_160),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_123),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_125),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_150),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_138),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_125),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_113),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_146),
.C(n_170),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_143),
.B(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_180),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_137),
.B(n_153),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_140),
.B1(n_149),
.B2(n_155),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_134),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_106),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_158),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_197),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_159),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_167),
.C(n_160),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_142),
.C(n_144),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_155),
.C(n_119),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_206),
.C(n_184),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_209),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_187),
.B1(n_179),
.B2(n_185),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_213),
.B1(n_181),
.B2(n_198),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_94),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_186),
.B(n_177),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_199),
.A2(n_185),
.B1(n_208),
.B2(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_59),
.C(n_53),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_220),
.B(n_172),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_200),
.A2(n_190),
.B1(n_177),
.B2(n_178),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_214),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_146),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_226),
.C(n_227),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_75),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_100),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_229),
.B(n_231),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_14),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_210),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_53),
.A3(n_21),
.B1(n_18),
.B2(n_15),
.C1(n_8),
.C2(n_10),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_239),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_219),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_211),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_228),
.B(n_218),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_242),
.B(n_2),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_215),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_245),
.B1(n_80),
.B2(n_241),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_80),
.B1(n_18),
.B2(n_15),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_235),
.C(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_2),
.C(n_3),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_250),
.B(n_3),
.C(n_4),
.D(n_6),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_80),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_253),
.B(n_4),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_249),
.C(n_8),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_12),
.C(n_13),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_12),
.Y(n_258)
);


endmodule