module fake_jpeg_1004_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

AOI21xp33_ASAP7_75t_SL g14 ( 
.A1(n_8),
.A2(n_0),
.B(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_17),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_6),
.B1(n_12),
.B2(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_20),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_20),
.C(n_22),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_28),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_4),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_28),
.B1(n_21),
.B2(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_30),
.B(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_37),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_32),
.C(n_4),
.Y(n_38)
);

NOR2xp67_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_35),
.Y(n_42)
);


endmodule