module real_aes_7861_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1205;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1170;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_792;
wire n_905;
wire n_518;
wire n_673;
wire n_1067;
wire n_878;
wire n_1192;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_1110;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1218;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_1217;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1123;
wire n_549;
wire n_571;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_1034;
wire n_1219;
wire n_952;
wire n_429;
wire n_1166;
wire n_1137;
wire n_448;
wire n_752;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_1220;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_528;
wire n_1078;
wire n_495;
wire n_578;
wire n_994;
wire n_1072;
wire n_938;
wire n_744;
wire n_1128;
wire n_935;
wire n_1098;
wire n_824;
wire n_1199;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_1213;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_1182;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_1189;
wire n_1180;
wire n_517;
wire n_931;
wire n_780;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1210;
wire n_1082;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_1025;
wire n_1168;
wire n_1148;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_725;
wire n_973;
wire n_504;
wire n_671;
wire n_1081;
wire n_960;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1207;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1196;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_1215;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_1100;
wire n_1167;
wire n_1174;
wire n_1193;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_1198;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_1212;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_1145;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1202;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_713;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_1179;
wire n_1201;
wire n_1171;
wire n_569;
wire n_563;
wire n_785;
wire n_997;
wire n_1203;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1136;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_1014;
wire n_1028;
wire n_1033;
wire n_1083;
wire n_727;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_1216;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_1127;
wire n_435;
wire n_972;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1187;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_1204;
wire n_486;
wire n_930;
wire n_1209;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_831;
wire n_487;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1071;
wire n_1052;
wire n_630;
wire n_1214;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_1208;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_717;
wire n_456;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_1172;
wire n_459;
wire n_558;
wire n_823;
wire n_863;
wire n_998;
wire n_1175;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_686;
wire n_776;
wire n_1190;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_1159;
wire n_1156;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_1211;
wire n_650;
wire n_710;
wire n_743;
wire n_1040;
wire n_703;
wire n_1097;
wire n_500;
wire n_601;
wire n_652;
wire n_661;
wire n_463;
wire n_1101;
wire n_804;
wire n_1076;
wire n_447;
wire n_1102;
wire n_1185;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_SL g970 ( .A1(n_0), .A2(n_69), .B1(n_971), .B2(n_973), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_1), .A2(n_313), .B1(n_686), .B2(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_2), .A2(n_322), .B1(n_995), .B2(n_1137), .Y(n_1214) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_3), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_4), .Y(n_854) );
INVx1_ASAP7_75t_L g1200 ( .A(n_5), .Y(n_1200) );
OA22x2_ASAP7_75t_L g1201 ( .A1(n_5), .A2(n_1200), .B1(n_1202), .B2(n_1218), .Y(n_1201) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_6), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_7), .A2(n_95), .B1(n_555), .B2(n_1012), .Y(n_1216) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_8), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_9), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_10), .A2(n_63), .B1(n_701), .B2(n_975), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g1091 ( .A1(n_11), .A2(n_21), .B1(n_774), .B2(n_1092), .C(n_1093), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_12), .A2(n_299), .B1(n_789), .B2(n_1077), .C(n_1078), .Y(n_1076) );
AOI22x1_ASAP7_75t_L g1122 ( .A1(n_13), .A2(n_1123), .B1(n_1151), .B2(n_1152), .Y(n_1122) );
INVx1_ASAP7_75t_L g1151 ( .A(n_13), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_14), .A2(n_155), .B1(n_555), .B2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_15), .Y(n_861) );
AO22x2_ASAP7_75t_L g431 ( .A1(n_16), .A2(n_247), .B1(n_423), .B2(n_428), .Y(n_431) );
INVx1_ASAP7_75t_L g1167 ( .A(n_16), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_17), .A2(n_180), .B1(n_417), .B2(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g1036 ( .A(n_18), .Y(n_1036) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_19), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_20), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_22), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_23), .A2(n_317), .B1(n_588), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_24), .A2(n_112), .B1(n_717), .B2(n_802), .Y(n_897) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_25), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_26), .Y(n_952) );
AOI222xp33_ASAP7_75t_L g974 ( .A1(n_27), .A2(n_64), .B1(n_169), .B2(n_491), .C1(n_526), .C2(n_975), .Y(n_974) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_28), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_29), .A2(n_271), .B1(n_631), .B2(n_632), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_30), .A2(n_176), .B1(n_538), .B2(n_703), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_31), .B(n_614), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_32), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_33), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_34), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_35), .A2(n_380), .B1(n_792), .B2(n_886), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_36), .A2(n_383), .B1(n_695), .B2(n_821), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_37), .A2(n_382), .B1(n_717), .B2(n_946), .Y(n_1217) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_38), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_39), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_40), .Y(n_947) );
AOI222xp33_ASAP7_75t_L g1067 ( .A1(n_41), .A2(n_68), .B1(n_369), .B2(n_489), .C1(n_973), .C2(n_1068), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_42), .A2(n_140), .B1(n_548), .B2(n_879), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g1211 ( .A(n_43), .Y(n_1211) );
CKINVDCx20_ASAP7_75t_R g990 ( .A(n_44), .Y(n_990) );
AO22x2_ASAP7_75t_L g433 ( .A1(n_45), .A2(n_124), .B1(n_423), .B2(n_424), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_46), .A2(n_1075), .B1(n_1097), .B2(n_1098), .Y(n_1074) );
INVx1_ASAP7_75t_L g1097 ( .A(n_46), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_47), .A2(n_393), .B1(n_455), .B2(n_724), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_48), .A2(n_232), .B1(n_626), .B2(n_794), .Y(n_1187) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_49), .A2(n_413), .B1(n_514), .B2(n_515), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_49), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_50), .A2(n_273), .B1(n_434), .B2(n_548), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_51), .A2(n_65), .B1(n_457), .B2(n_632), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_52), .A2(n_181), .B1(n_964), .B2(n_1012), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_53), .A2(n_304), .B1(n_555), .B2(n_649), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_54), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_55), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_56), .A2(n_211), .B1(n_417), .B2(n_434), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_57), .A2(n_323), .B1(n_527), .B2(n_541), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_58), .A2(n_240), .B1(n_495), .B2(n_527), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_59), .B(n_775), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g1145 ( .A(n_60), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_61), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_62), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_66), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_67), .A2(n_396), .B1(n_628), .B2(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_70), .A2(n_266), .B1(n_631), .B2(n_632), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_71), .A2(n_312), .B1(n_635), .B2(n_638), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_72), .A2(n_892), .B1(n_919), .B2(n_920), .Y(n_891) );
INVx1_ASAP7_75t_L g919 ( .A(n_72), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_73), .A2(n_147), .B1(n_725), .B2(n_1137), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_74), .A2(n_348), .B1(n_447), .B2(n_902), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_75), .A2(n_598), .B1(n_641), .B2(n_642), .Y(n_597) );
INVx1_ASAP7_75t_L g641 ( .A(n_75), .Y(n_641) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_76), .A2(n_300), .B1(n_551), .B2(n_552), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_77), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_78), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_79), .A2(n_206), .B1(n_624), .B2(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_80), .A2(n_170), .B1(n_455), .B2(n_1047), .Y(n_1215) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_81), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_82), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_83), .A2(n_118), .B1(n_548), .B2(n_580), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_84), .Y(n_771) );
INVx1_ASAP7_75t_L g968 ( .A(n_85), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_86), .A2(n_113), .B1(n_792), .B2(n_995), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_87), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_88), .A2(n_276), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_89), .A2(n_308), .B1(n_366), .B2(n_489), .C1(n_614), .C2(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_90), .A2(n_285), .B1(n_527), .B2(n_541), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_91), .A2(n_343), .B1(n_502), .B2(n_526), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_92), .A2(n_321), .B1(n_470), .B2(n_546), .Y(n_1066) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_93), .Y(n_492) );
INVx1_ASAP7_75t_L g645 ( .A(n_94), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_96), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_97), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1140 ( .A(n_98), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_99), .A2(n_150), .B1(n_845), .B2(n_1029), .Y(n_1028) );
AO22x2_ASAP7_75t_L g427 ( .A1(n_100), .A2(n_277), .B1(n_423), .B2(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g1164 ( .A(n_100), .Y(n_1164) );
CKINVDCx20_ASAP7_75t_R g1106 ( .A(n_101), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_102), .A2(n_103), .B1(n_470), .B2(n_588), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_104), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_105), .A2(n_122), .B1(n_582), .B2(n_633), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_106), .A2(n_252), .B1(n_503), .B2(n_541), .Y(n_750) );
OA22x2_ASAP7_75t_L g925 ( .A1(n_107), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_107), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_108), .A2(n_168), .B1(n_792), .B2(n_794), .Y(n_791) );
AOI222xp33_ASAP7_75t_L g1096 ( .A1(n_109), .A2(n_121), .B1(n_154), .B2(n_489), .C1(n_494), .C2(n_1068), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_110), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_111), .Y(n_918) );
INVx1_ASAP7_75t_L g738 ( .A(n_114), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_115), .A2(n_358), .B1(n_695), .B2(n_696), .C(n_697), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_116), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_117), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_119), .A2(n_204), .B1(n_538), .B2(n_611), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_120), .A2(n_237), .B1(n_631), .B2(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_123), .A2(n_172), .B1(n_466), .B2(n_552), .Y(n_853) );
INVx1_ASAP7_75t_L g1168 ( .A(n_124), .Y(n_1168) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_125), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_126), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_127), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_128), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_129), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g1205 ( .A(n_130), .Y(n_1205) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_131), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_132), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g1134 ( .A(n_133), .Y(n_1134) );
CKINVDCx20_ASAP7_75t_R g1180 ( .A(n_134), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_135), .A2(n_316), .B1(n_546), .B2(n_803), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_136), .A2(n_298), .B1(n_624), .B2(n_900), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g1141 ( .A(n_137), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_138), .A2(n_339), .B1(n_691), .B2(n_789), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_139), .A2(n_250), .B1(n_725), .B2(n_902), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_141), .A2(n_258), .B1(n_775), .B2(n_821), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_142), .A2(n_336), .B1(n_436), .B2(n_548), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_143), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_144), .B(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_145), .A2(n_198), .B1(n_573), .B2(n_703), .Y(n_1111) );
AOI22xp33_ASAP7_75t_SL g1114 ( .A1(n_146), .A2(n_331), .B1(n_588), .B2(n_886), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_148), .A2(n_192), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_149), .A2(n_361), .B1(n_503), .B2(n_573), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_151), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_152), .A2(n_340), .B1(n_495), .B2(n_777), .Y(n_1040) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_153), .A2(n_355), .B1(n_538), .B2(n_541), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g1182 ( .A1(n_156), .A2(n_214), .B1(n_777), .B2(n_973), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_157), .A2(n_359), .B1(n_626), .B2(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_158), .A2(n_338), .B1(n_1131), .B2(n_1132), .Y(n_1130) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_159), .A2(n_341), .B1(n_631), .B2(n_632), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_160), .A2(n_221), .B1(n_557), .B2(n_1047), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_161), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_162), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_163), .B(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_164), .A2(n_226), .B1(n_649), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_165), .A2(n_263), .B1(n_640), .B2(n_961), .Y(n_960) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_166), .Y(n_767) );
AND2x6_ASAP7_75t_L g401 ( .A(n_167), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1161 ( .A(n_167), .Y(n_1161) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_171), .A2(n_188), .B1(n_470), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_173), .A2(n_305), .B1(n_778), .B2(n_1027), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_174), .A2(n_196), .B1(n_546), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_175), .A2(n_288), .B1(n_582), .B2(n_583), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_177), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g1094 ( .A(n_178), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_179), .A2(n_287), .B1(n_441), .B2(n_457), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_182), .A2(n_307), .B1(n_526), .B2(n_527), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g1044 ( .A(n_183), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_184), .A2(n_335), .B1(n_586), .B2(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g1110 ( .A(n_185), .B(n_695), .Y(n_1110) );
AO22x2_ASAP7_75t_L g422 ( .A1(n_186), .A2(n_264), .B1(n_423), .B2(n_424), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g1165 ( .A(n_186), .B(n_1166), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_187), .B(n_913), .Y(n_912) );
CKINVDCx20_ASAP7_75t_R g1147 ( .A(n_189), .Y(n_1147) );
AOI22xp33_ASAP7_75t_SL g1117 ( .A1(n_190), .A2(n_283), .B1(n_946), .B2(n_1012), .Y(n_1117) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_191), .Y(n_800) );
AOI211xp5_ASAP7_75t_L g769 ( .A1(n_193), .A2(n_523), .B(n_770), .C(n_780), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_194), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_195), .A2(n_379), .B1(n_635), .B2(n_638), .Y(n_1049) );
AOI22xp33_ASAP7_75t_SL g1107 ( .A1(n_197), .A2(n_294), .B1(n_502), .B2(n_541), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_199), .A2(n_205), .B1(n_557), .B2(n_959), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_200), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_201), .Y(n_982) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_202), .Y(n_984) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_203), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_207), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_208), .A2(n_249), .B1(n_633), .B2(n_692), .Y(n_849) );
AOI22xp33_ASAP7_75t_SL g1116 ( .A1(n_209), .A2(n_225), .B1(n_633), .B2(n_720), .Y(n_1116) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_210), .A2(n_253), .B1(n_559), .B2(n_588), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_212), .A2(n_399), .B(n_407), .C(n_1169), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g1208 ( .A(n_213), .Y(n_1208) );
CKINVDCx20_ASAP7_75t_R g1090 ( .A(n_215), .Y(n_1090) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_216), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_217), .A2(n_346), .B1(n_724), .B2(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_218), .A2(n_397), .B1(n_466), .B2(n_692), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_219), .B(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_220), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_222), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_223), .A2(n_388), .B1(n_588), .B2(n_763), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g1178 ( .A(n_224), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_227), .A2(n_320), .B1(n_465), .B2(n_763), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_228), .A2(n_330), .B1(n_457), .B2(n_551), .Y(n_852) );
AOI22xp33_ASAP7_75t_SL g1113 ( .A1(n_229), .A2(n_377), .B1(n_455), .B2(n_626), .Y(n_1113) );
CKINVDCx20_ASAP7_75t_R g1060 ( .A(n_230), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_231), .B(n_614), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_233), .A2(n_280), .B1(n_546), .B2(n_548), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_234), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_235), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g1129 ( .A(n_236), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_238), .A2(n_246), .B1(n_502), .B2(n_987), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_239), .A2(n_360), .B1(n_436), .B2(n_1051), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_241), .Y(n_687) );
XNOR2x2_ASAP7_75t_L g955 ( .A(n_242), .B(n_956), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_243), .A2(n_279), .B1(n_470), .B2(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_244), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_245), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_248), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_251), .A2(n_296), .B1(n_611), .B2(n_913), .Y(n_1209) );
OA22x2_ASAP7_75t_L g561 ( .A1(n_254), .A2(n_562), .B1(n_563), .B2(n_589), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_254), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_255), .A2(n_392), .B1(n_447), .B2(n_828), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_256), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_257), .B(n_696), .Y(n_1109) );
XNOR2x2_ASAP7_75t_L g1007 ( .A(n_259), .B(n_1008), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_260), .A2(n_386), .B1(n_559), .B2(n_789), .Y(n_1186) );
INVx2_ASAP7_75t_L g406 ( .A(n_261), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_262), .A2(n_713), .B1(n_739), .B2(n_740), .Y(n_712) );
INVx1_ASAP7_75t_L g739 ( .A(n_262), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g997 ( .A1(n_265), .A2(n_278), .B1(n_635), .B2(n_879), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_267), .A2(n_1171), .B1(n_1172), .B2(n_1191), .Y(n_1170) );
CKINVDCx20_ASAP7_75t_R g1191 ( .A(n_267), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_268), .B(n_845), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_269), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g819 ( .A1(n_270), .A2(n_301), .B1(n_542), .B2(n_777), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_272), .A2(n_394), .B1(n_466), .B2(n_559), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_274), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_275), .A2(n_390), .B1(n_555), .B2(n_557), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_281), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g1080 ( .A(n_282), .Y(n_1080) );
CKINVDCx20_ASAP7_75t_R g1206 ( .A(n_284), .Y(n_1206) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_286), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_289), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_290), .A2(n_387), .B1(n_626), .B2(n_628), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_291), .A2(n_391), .B1(n_881), .B2(n_946), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_292), .A2(n_670), .B1(n_704), .B2(n_705), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_292), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_293), .A2(n_374), .B1(n_440), .B2(n_447), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_295), .Y(n_951) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_297), .Y(n_566) );
OA22x2_ASAP7_75t_L g810 ( .A1(n_302), .A2(n_811), .B1(n_812), .B2(n_833), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_302), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_303), .B(n_534), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_306), .A2(n_332), .B1(n_885), .B2(n_886), .Y(n_884) );
INVx1_ASAP7_75t_L g423 ( .A(n_309), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_309), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_310), .A2(n_389), .B1(n_548), .B2(n_582), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g938 ( .A(n_311), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_314), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_315), .Y(n_1150) );
CKINVDCx20_ASAP7_75t_R g907 ( .A(n_318), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_319), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g1082 ( .A1(n_324), .A2(n_342), .B1(n_635), .B2(n_1083), .C(n_1086), .Y(n_1082) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_325), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_326), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_327), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g1177 ( .A(n_328), .Y(n_1177) );
INVx1_ASAP7_75t_L g728 ( .A(n_329), .Y(n_728) );
INVx1_ASAP7_75t_L g905 ( .A(n_333), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_334), .B(n_1062), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_337), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_344), .A2(n_376), .B1(n_546), .B2(n_559), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_345), .A2(n_365), .B1(n_539), .B2(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g405 ( .A(n_347), .B(n_406), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g1212 ( .A(n_349), .Y(n_1212) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_350), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g1118 ( .A(n_351), .Y(n_1118) );
INVx1_ASAP7_75t_L g402 ( .A(n_352), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_353), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g1087 ( .A(n_354), .Y(n_1087) );
OA22x2_ASAP7_75t_L g517 ( .A1(n_356), .A2(n_518), .B1(n_519), .B2(n_560), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_356), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_357), .B(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_362), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_363), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_364), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g1126 ( .A(n_367), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_368), .Y(n_781) );
INVx1_ASAP7_75t_L g999 ( .A(n_370), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_371), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_372), .B(n_778), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_373), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_375), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_378), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g1135 ( .A(n_381), .Y(n_1135) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_384), .Y(n_677) );
INVx1_ASAP7_75t_L g764 ( .A(n_385), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_395), .Y(n_616) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_402), .Y(n_1160) );
OAI21xp5_ASAP7_75t_L g1198 ( .A1(n_403), .A2(n_1159), .B(n_1199), .Y(n_1198) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_1003), .B1(n_1154), .B2(n_1155), .C(n_1156), .Y(n_407) );
INVxp67_ASAP7_75t_L g1154 ( .A(n_408), .Y(n_1154) );
XOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_707), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_592), .B2(n_706), .Y(n_409) );
INVx2_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
OA22x2_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_516), .B1(n_590), .B2(n_591), .Y(n_411) );
INVx1_ASAP7_75t_L g590 ( .A(n_412), .Y(n_590) );
INVx1_ASAP7_75t_L g515 ( .A(n_413), .Y(n_515) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_414), .B(n_473), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_452), .C(n_462), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_439), .Y(n_415) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g624 ( .A(n_418), .Y(n_624) );
INVx3_ASAP7_75t_L g790 ( .A(n_418), .Y(n_790) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_418), .Y(n_964) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g547 ( .A(n_419), .Y(n_547) );
BUFx2_ASAP7_75t_SL g946 ( .A(n_419), .Y(n_946) );
BUFx2_ASAP7_75t_SL g1051 ( .A(n_419), .Y(n_1051) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_429), .Y(n_419) );
AND2x6_ASAP7_75t_L g436 ( .A(n_420), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g457 ( .A(n_420), .B(n_446), .Y(n_457) );
AND2x6_ASAP7_75t_L g491 ( .A(n_420), .B(n_484), .Y(n_491) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_426), .Y(n_420) );
AND2x2_ASAP7_75t_L g467 ( .A(n_421), .B(n_427), .Y(n_467) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g444 ( .A(n_422), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_422), .B(n_427), .Y(n_451) );
AND2x2_ASAP7_75t_L g477 ( .A(n_422), .B(n_431), .Y(n_477) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_425), .Y(n_428) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g445 ( .A(n_427), .Y(n_445) );
INVx1_ASAP7_75t_L g498 ( .A(n_427), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_429), .B(n_444), .Y(n_461) );
AND2x4_ASAP7_75t_L g466 ( .A(n_429), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g471 ( .A(n_429), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g549 ( .A(n_429), .B(n_444), .Y(n_549) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
OR2x2_ASAP7_75t_L g438 ( .A(n_430), .B(n_433), .Y(n_438) );
AND2x2_ASAP7_75t_L g446 ( .A(n_430), .B(n_433), .Y(n_446) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g484 ( .A(n_431), .B(n_433), .Y(n_484) );
INVx1_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
AND2x2_ASAP7_75t_L g497 ( .A(n_432), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g450 ( .A(n_433), .Y(n_450) );
INVx2_ASAP7_75t_L g950 ( .A(n_434), .Y(n_950) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx5_ASAP7_75t_SL g692 ( .A(n_435), .Y(n_692) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_435), .Y(n_825) );
INVx2_ASAP7_75t_L g959 ( .A(n_435), .Y(n_959) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_435), .Y(n_1085) );
INVx4_ASAP7_75t_L g1131 ( .A(n_435), .Y(n_1131) );
INVx11_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx11_ASAP7_75t_L g556 ( .A(n_436), .Y(n_556) );
AND2x4_ASAP7_75t_L g536 ( .A(n_437), .B(n_467), .Y(n_536) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g508 ( .A(n_438), .B(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx4_ASAP7_75t_L g551 ( .A(n_442), .Y(n_551) );
INVx5_ASAP7_75t_L g586 ( .A(n_442), .Y(n_586) );
BUFx3_ASAP7_75t_L g627 ( .A(n_442), .Y(n_627) );
INVx3_ASAP7_75t_L g761 ( .A(n_442), .Y(n_761) );
INVx2_ASAP7_75t_L g828 ( .A(n_442), .Y(n_828) );
INVx8_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_444), .B(n_446), .Y(n_679) );
INVx1_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_446), .B(n_467), .Y(n_513) );
AND2x6_ASAP7_75t_L g532 ( .A(n_446), .B(n_467), .Y(n_532) );
INVx1_ASAP7_75t_L g1081 ( .A(n_447), .Y(n_1081) );
BUFx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g628 ( .A(n_448), .Y(n_628) );
BUFx4f_ASAP7_75t_SL g725 ( .A(n_448), .Y(n_725) );
BUFx2_ASAP7_75t_L g763 ( .A(n_448), .Y(n_763) );
BUFx2_ASAP7_75t_L g886 ( .A(n_448), .Y(n_886) );
INVx6_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g552 ( .A(n_449), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_449), .A2(n_482), .B1(n_575), .B2(n_576), .Y(n_574) );
INVx1_ASAP7_75t_SL g794 ( .A(n_449), .Y(n_794) );
INVx1_ASAP7_75t_L g995 ( .A(n_449), .Y(n_995) );
OR2x6_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g540 ( .A(n_450), .Y(n_540) );
INVx1_ASAP7_75t_L g472 ( .A(n_451), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_458), .B2(n_459), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g557 ( .A(n_456), .Y(n_557) );
INVx2_ASAP7_75t_L g686 ( .A(n_456), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_456), .A2(n_953), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
INVx2_ASAP7_75t_L g1057 ( .A(n_456), .Y(n_1057) );
INVx6_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g582 ( .A(n_457), .Y(n_582) );
BUFx3_ASAP7_75t_L g631 ( .A(n_457), .Y(n_631) );
BUFx3_ASAP7_75t_L g1089 ( .A(n_457), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_459), .A2(n_684), .B1(n_685), .B2(n_687), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_459), .A2(n_685), .B1(n_796), .B2(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g953 ( .A(n_460), .Y(n_953) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_468), .B2(n_469), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_464), .A2(n_689), .B1(n_690), .B2(n_693), .Y(n_688) );
INVx1_ASAP7_75t_L g831 ( .A(n_464), .Y(n_831) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g588 ( .A(n_466), .Y(n_588) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_466), .Y(n_637) );
INVx2_ASAP7_75t_L g718 ( .A(n_466), .Y(n_718) );
BUFx3_ASAP7_75t_L g885 ( .A(n_466), .Y(n_885) );
INVx1_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g559 ( .A(n_471), .Y(n_559) );
BUFx3_ASAP7_75t_L g640 ( .A(n_471), .Y(n_640) );
BUFx3_ASAP7_75t_L g803 ( .A(n_471), .Y(n_803) );
BUFx2_ASAP7_75t_SL g881 ( .A(n_471), .Y(n_881) );
BUFx2_ASAP7_75t_SL g1012 ( .A(n_471), .Y(n_1012) );
BUFx3_ASAP7_75t_L g1077 ( .A(n_471), .Y(n_1077) );
AND2x2_ASAP7_75t_L g651 ( .A(n_472), .B(n_478), .Y(n_651) );
NOR3xp33_ASAP7_75t_SL g473 ( .A(n_474), .B(n_487), .C(n_505), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_479), .B2(n_480), .Y(n_474) );
INVx4_ASAP7_75t_L g618 ( .A(n_476), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_476), .A2(n_482), .B1(n_698), .B2(n_699), .Y(n_697) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_476), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_476), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
BUFx3_ASAP7_75t_L g875 ( .A(n_476), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_476), .A2(n_620), .B1(n_1205), .B2(n_1206), .Y(n_1204) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x4_ASAP7_75t_L g496 ( .A(n_477), .B(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g503 ( .A(n_477), .B(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g539 ( .A(n_477), .B(n_540), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_480), .A2(n_617), .B1(n_989), .B2(n_990), .Y(n_988) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g620 ( .A(n_481), .Y(n_620) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_482), .Y(n_1043) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g542 ( .A(n_484), .B(n_486), .Y(n_542) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_492), .B1(n_493), .B2(n_499), .C(n_500), .Y(n_487) );
OAI221xp5_ASAP7_75t_SL g608 ( .A1(n_488), .A2(n_609), .B1(n_610), .B2(n_612), .C(n_613), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g730 ( .A1(n_488), .A2(n_731), .B1(n_732), .B2(n_733), .C(n_734), .Y(n_730) );
OAI21xp33_ASAP7_75t_SL g1038 ( .A1(n_488), .A2(n_1039), .B(n_1040), .Y(n_1038) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI21xp5_ASAP7_75t_SL g748 ( .A1(n_490), .A2(n_749), .B(n_750), .Y(n_748) );
BUFx2_ASAP7_75t_L g985 ( .A(n_490), .Y(n_985) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g523 ( .A(n_491), .Y(n_523) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_491), .Y(n_580) );
INVx2_ASAP7_75t_L g815 ( .A(n_491), .Y(n_815) );
INVx2_ASAP7_75t_SL g909 ( .A(n_491), .Y(n_909) );
INVx2_ASAP7_75t_L g1105 ( .A(n_491), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_493), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_493), .A2(n_909), .B1(n_910), .B2(n_911), .C(n_912), .Y(n_908) );
OAI222xp33_ASAP7_75t_L g1142 ( .A1(n_493), .A2(n_1143), .B1(n_1144), .B2(n_1145), .C1(n_1146), .C2(n_1147), .Y(n_1142) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g753 ( .A(n_494), .Y(n_753) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g873 ( .A(n_495), .Y(n_873) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx4f_ASAP7_75t_SL g526 ( .A(n_496), .Y(n_526) );
BUFx2_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_496), .Y(n_611) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_496), .Y(n_703) );
INVx1_ASAP7_75t_L g504 ( .A(n_498), .Y(n_504) );
BUFx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx3_ASAP7_75t_L g614 ( .A(n_502), .Y(n_614) );
INVx2_ASAP7_75t_L g914 ( .A(n_502), .Y(n_914) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx12f_ASAP7_75t_L g527 ( .A(n_503), .Y(n_527) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_503), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_510), .B2(n_511), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_507), .A2(n_607), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g869 ( .A(n_507), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_507), .A2(n_511), .B1(n_1211), .B2(n_1212), .Y(n_1210) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx3_ASAP7_75t_L g567 ( .A(n_508), .Y(n_567) );
INVx2_ASAP7_75t_L g603 ( .A(n_508), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_508), .A2(n_607), .B1(n_656), .B2(n_657), .C(n_658), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_511), .A2(n_868), .B1(n_1036), .B2(n_1037), .Y(n_1035) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_SL g569 ( .A(n_512), .Y(n_569) );
INVx1_ASAP7_75t_L g747 ( .A(n_512), .Y(n_747) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g607 ( .A(n_513), .Y(n_607) );
INVx1_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
XOR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_561), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_517), .A2(n_643), .B1(n_644), .B2(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_517), .Y(n_667) );
INVx1_ASAP7_75t_L g560 ( .A(n_519), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_543), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g520 ( .A(n_521), .B(n_528), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_524), .B(n_525), .Y(n_521) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_522), .A2(n_661), .B(n_662), .Y(n_660) );
OAI21xp33_ASAP7_75t_L g933 ( .A1(n_522), .A2(n_934), .B(n_935), .Y(n_933) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g785 ( .A(n_527), .Y(n_785) );
BUFx4f_ASAP7_75t_SL g1068 ( .A(n_527), .Y(n_1068) );
NAND3xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .C(n_537), .Y(n_528) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_SL g821 ( .A(n_531), .Y(n_821) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g696 ( .A(n_532), .Y(n_696) );
BUFx2_ASAP7_75t_L g845 ( .A(n_532), .Y(n_845) );
BUFx4f_ASAP7_75t_L g1092 ( .A(n_532), .Y(n_1092) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_534), .Y(n_695) );
INVx5_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g775 ( .A(n_535), .Y(n_775) );
INVx2_ASAP7_75t_L g1029 ( .A(n_535), .Y(n_1029) );
INVx2_ASAP7_75t_L g1062 ( .A(n_535), .Y(n_1062) );
INVx4_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g573 ( .A(n_539), .Y(n_573) );
BUFx2_ASAP7_75t_L g777 ( .A(n_539), .Y(n_777) );
INVx1_ASAP7_75t_L g972 ( .A(n_539), .Y(n_972) );
BUFx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_542), .Y(n_659) );
BUFx2_ASAP7_75t_SL g973 ( .A(n_542), .Y(n_973) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_553), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .Y(n_544) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g649 ( .A(n_547), .Y(n_649) );
BUFx2_ASAP7_75t_L g896 ( .A(n_548), .Y(n_896) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
BUFx3_ASAP7_75t_L g965 ( .A(n_549), .Y(n_965) );
BUFx3_ASAP7_75t_L g1047 ( .A(n_549), .Y(n_1047) );
INVx2_ASAP7_75t_L g793 ( .A(n_551), .Y(n_793) );
BUFx6f_ASAP7_75t_L g902 ( .A(n_551), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_558), .Y(n_553) );
INVx4_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI21xp33_ASAP7_75t_SL g570 ( .A1(n_556), .A2(n_571), .B(n_572), .Y(n_570) );
INVx4_ASAP7_75t_L g720 ( .A(n_556), .Y(n_720) );
INVx2_ASAP7_75t_SL g879 ( .A(n_556), .Y(n_879) );
INVx3_ASAP7_75t_L g900 ( .A(n_556), .Y(n_900) );
INVx2_ASAP7_75t_L g589 ( .A(n_563), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_577), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_570), .C(n_574), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_567), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_569), .A2(n_905), .B1(n_906), .B2(n_907), .Y(n_904) );
OA211x2_ASAP7_75t_L g1059 ( .A1(n_569), .A2(n_1060), .B(n_1061), .C(n_1063), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_584), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx2_ASAP7_75t_L g860 ( .A(n_580), .Y(n_860) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_580), .Y(n_1144) );
INVx1_ASAP7_75t_L g732 ( .A(n_583), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_586), .Y(n_724) );
BUFx2_ASAP7_75t_L g1137 ( .A(n_586), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_588), .Y(n_1128) );
INVx1_ASAP7_75t_L g706 ( .A(n_592), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_663), .B2(n_664), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_597), .B1(n_643), .B2(n_644), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g642 ( .A(n_598), .Y(n_642) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_621), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_608), .C(n_615), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_600) );
OAI22xp5_ASAP7_75t_SL g930 ( .A1(n_602), .A2(n_605), .B1(n_931), .B2(n_932), .Y(n_930) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g906 ( .A(n_603), .Y(n_906) );
INVx1_ASAP7_75t_SL g981 ( .A(n_603), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_605), .A2(n_867), .B1(n_868), .B2(n_870), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_605), .A2(n_980), .B1(n_981), .B2(n_982), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_605), .A2(n_868), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx3_ASAP7_75t_L g772 ( .A(n_607), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_610), .A2(n_875), .B1(n_937), .B2(n_938), .Y(n_936) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g1146 ( .A(n_614), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_619), .B2(n_620), .Y(n_615) );
INVx3_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g917 ( .A(n_618), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_620), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_620), .A2(n_916), .B1(n_917), .B2(n_918), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_620), .A2(n_917), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_620), .A2(n_917), .B1(n_1149), .B2(n_1150), .Y(n_1148) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_629), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVxp67_ASAP7_75t_L g681 ( .A(n_628), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
BUFx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx4_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g961 ( .A(n_636), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_636), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
INVx4_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_639), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_672) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_640), .Y(n_1132) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
XNOR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NOR4xp75_ASAP7_75t_L g646 ( .A(n_647), .B(n_652), .C(n_655), .D(n_660), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVxp67_ASAP7_75t_L g674 ( .A(n_649), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_SL g779 ( .A(n_659), .Y(n_779) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI22xp5_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_666), .B1(n_668), .B2(n_669), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g705 ( .A(n_670), .Y(n_705) );
AND4x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_682), .C(n_694), .D(n_700), .Y(n_670) );
NOR2xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_676), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_680), .B2(n_681), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_678), .A2(n_1079), .B1(n_1080), .B2(n_1081), .Y(n_1078) );
BUFx2_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_688), .Y(n_682) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g1016 ( .A(n_692), .Y(n_1016) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx4_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g987 ( .A(n_703), .Y(n_987) );
INVx2_ASAP7_75t_L g1176 ( .A(n_703), .Y(n_1176) );
XOR2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_806), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_SL g709 ( .A1(n_710), .A2(n_766), .B1(n_804), .B2(n_805), .Y(n_709) );
INVx1_ASAP7_75t_L g804 ( .A(n_710), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_741), .B2(n_765), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g740 ( .A(n_713), .Y(n_740) );
AND2x2_ASAP7_75t_SL g713 ( .A(n_714), .B(n_726), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_721), .Y(n_714) );
NAND2xp33_ASAP7_75t_SL g715 ( .A(n_716), .B(n_719), .Y(n_715) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_718), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .C(n_735), .Y(n_726) );
INVx1_ASAP7_75t_L g765 ( .A(n_741), .Y(n_765) );
XOR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_764), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_755), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .C(n_751), .Y(n_743) );
OA211x2_ASAP7_75t_L g967 ( .A1(n_747), .A2(n_968), .B(n_969), .C(n_970), .Y(n_967) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx2_ASAP7_75t_L g805 ( .A(n_766), .Y(n_805) );
XNOR2x1_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_786), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B(n_773), .C(n_776), .Y(n_770) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_795), .C(n_798), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI221xp5_ASAP7_75t_SL g1125 ( .A1(n_790), .A2(n_1126), .B1(n_1127), .B2(n_1129), .C(n_1130), .Y(n_1125) );
INVx3_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
BUFx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
XNOR2xp5_ASAP7_75t_SL g806 ( .A(n_807), .B(n_889), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_834), .B2(n_835), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_SL g833 ( .A(n_812), .Y(n_833) );
NAND3x1_ASAP7_75t_L g812 ( .A(n_813), .B(n_822), .C(n_829), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_818), .Y(n_813) );
OAI21xp5_ASAP7_75t_SL g814 ( .A1(n_815), .A2(n_816), .B(n_817), .Y(n_814) );
OAI21xp5_ASAP7_75t_SL g839 ( .A1(n_815), .A2(n_840), .B(n_841), .Y(n_839) );
OAI21xp5_ASAP7_75t_SL g1022 ( .A1(n_815), .A2(n_1023), .B(n_1024), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_826), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AND2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_832), .Y(n_829) );
INVx2_ASAP7_75t_SL g834 ( .A(n_835), .Y(n_834) );
AO22x2_ASAP7_75t_SL g835 ( .A1(n_836), .A2(n_855), .B1(n_856), .B2(n_888), .Y(n_835) );
INVx3_ASAP7_75t_L g888 ( .A(n_836), .Y(n_888) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_854), .Y(n_836) );
NAND2x1_ASAP7_75t_SL g837 ( .A(n_838), .B(n_847), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_842), .Y(n_838) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .C(n_846), .Y(n_842) );
NOR2x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_851), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
XOR2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_887), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_876), .Y(n_857) );
NOR3xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_866), .C(n_871), .Y(n_858) );
OAI221xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B1(n_862), .B2(n_864), .C(n_865), .Y(n_859) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
BUFx4f_ASAP7_75t_L g975 ( .A(n_863), .Y(n_975) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_873), .B1(n_874), .B2(n_875), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_882), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
INVx1_ASAP7_75t_SL g948 ( .A(n_881), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_921), .B1(n_1001), .B2(n_1002), .Y(n_889) );
INVx2_ASAP7_75t_L g1001 ( .A(n_890), .Y(n_1001) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g920 ( .A(n_892), .Y(n_920) );
AND2x2_ASAP7_75t_SL g892 ( .A(n_893), .B(n_903), .Y(n_892) );
NOR2xp33_ASAP7_75t_SL g893 ( .A(n_894), .B(n_898), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_895), .B(n_897), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_901), .Y(n_898) );
NOR3xp33_ASAP7_75t_L g903 ( .A(n_904), .B(n_908), .C(n_915), .Y(n_903) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_SL g1041 ( .A1(n_914), .A2(n_1042), .B1(n_1043), .B2(n_1044), .Y(n_1041) );
INVx1_ASAP7_75t_L g1002 ( .A(n_921), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B1(n_976), .B2(n_1000), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_925), .B1(n_954), .B2(n_955), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_SL g927 ( .A(n_928), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_929), .B(n_939), .Y(n_928) );
NOR3xp33_ASAP7_75t_L g929 ( .A(n_930), .B(n_933), .C(n_936), .Y(n_929) );
NOR3xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_943), .C(n_949), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_944), .A2(n_945), .B1(n_947), .B2(n_948), .Y(n_943) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_951), .B1(n_952), .B2(n_953), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_953), .A2(n_1087), .B1(n_1088), .B2(n_1090), .Y(n_1086) );
OAI221xp5_ASAP7_75t_SL g1133 ( .A1(n_953), .A2(n_1088), .B1(n_1134), .B2(n_1135), .C(n_1136), .Y(n_1133) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NAND4xp75_ASAP7_75t_L g956 ( .A(n_957), .B(n_962), .C(n_967), .D(n_974), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_958), .B(n_960), .Y(n_957) );
AND2x2_ASAP7_75t_L g962 ( .A(n_963), .B(n_966), .Y(n_962) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g1027 ( .A(n_972), .Y(n_1027) );
INVx1_ASAP7_75t_L g1179 ( .A(n_975), .Y(n_1179) );
INVx1_ASAP7_75t_L g1000 ( .A(n_976), .Y(n_1000) );
XOR2x2_ASAP7_75t_L g976 ( .A(n_977), .B(n_999), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_991), .Y(n_977) );
NOR3xp33_ASAP7_75t_L g978 ( .A(n_979), .B(n_983), .C(n_988), .Y(n_978) );
OAI21xp33_ASAP7_75t_L g983 ( .A1(n_984), .A2(n_985), .B(n_986), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_996), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1003), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B1(n_1122), .B2(n_1153), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_1006), .A2(n_1072), .B1(n_1120), .B2(n_1121), .Y(n_1005) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1006), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1030), .B1(n_1070), .B2(n_1071), .Y(n_1006) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1007), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1099 ( .A1(n_1007), .A2(n_1070), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
NAND2xp5_ASAP7_75t_SL g1008 ( .A(n_1009), .B(n_1021), .Y(n_1008) );
NOR3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1014), .C(n_1018), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1013), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1025), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1028), .Y(n_1025) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1030), .Y(n_1071) );
XNOR2xp5_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1052), .Y(n_1030) );
XNOR2x1_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1045), .Y(n_1033) );
NOR3xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1038), .C(n_1041), .Y(n_1034) );
AND4x1_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1048), .C(n_1049), .D(n_1050), .Y(n_1045) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
XOR2x2_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1069), .Y(n_1053) );
NAND4xp75_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1059), .C(n_1064), .D(n_1067), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1058), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1066), .Y(n_1064) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1072), .Y(n_1120) );
OAI22xp5_ASAP7_75t_SL g1072 ( .A1(n_1073), .A2(n_1074), .B1(n_1099), .B2(n_1119), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1075), .Y(n_1098) );
AND4x1_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1082), .C(n_1091), .D(n_1096), .Y(n_1075) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx3_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1099), .Y(n_1119) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
XOR2x2_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1118), .Y(n_1101) );
NAND3x1_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1112), .C(n_1115), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1108), .Y(n_1103) );
OAI21xp5_ASAP7_75t_SL g1104 ( .A1(n_1105), .A2(n_1106), .B(n_1107), .Y(n_1104) );
OAI21xp33_ASAP7_75t_L g1207 ( .A1(n_1105), .A2(n_1208), .B(n_1209), .Y(n_1207) );
NAND3xp33_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .C(n_1111), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1122), .Y(n_1153) );
INVx1_ASAP7_75t_SL g1152 ( .A(n_1123), .Y(n_1152) );
AND2x2_ASAP7_75t_SL g1123 ( .A(n_1124), .B(n_1138), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1133), .Y(n_1124) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NOR3xp33_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1142), .C(n_1148), .Y(n_1138) );
OAI222xp33_ASAP7_75t_L g1175 ( .A1(n_1144), .A2(n_1176), .B1(n_1177), .B2(n_1178), .C1(n_1179), .C2(n_1180), .Y(n_1175) );
INVx1_ASAP7_75t_SL g1156 ( .A(n_1157), .Y(n_1156) );
NOR2x1_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1162), .Y(n_1157) );
OR2x2_ASAP7_75t_SL g1221 ( .A(n_1158), .B(n_1163), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1161), .Y(n_1158) );
CKINVDCx20_ASAP7_75t_R g1193 ( .A(n_1159), .Y(n_1193) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1160), .B(n_1196), .Y(n_1199) );
CKINVDCx16_ASAP7_75t_R g1196 ( .A(n_1161), .Y(n_1196) );
CKINVDCx20_ASAP7_75t_R g1162 ( .A(n_1163), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1165), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1168), .Y(n_1166) );
OAI322xp33_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1192), .A3(n_1194), .B1(n_1197), .B2(n_1200), .C1(n_1201), .C2(n_1219), .Y(n_1169) );
CKINVDCx20_ASAP7_75t_R g1171 ( .A(n_1172), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1184), .Y(n_1173) );
NOR2x1_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1181), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1183), .Y(n_1181) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1188), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1187), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
CKINVDCx16_ASAP7_75t_R g1197 ( .A(n_1198), .Y(n_1197) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1202), .Y(n_1218) );
NAND2x1_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1213), .Y(n_1202) );
NOR3xp33_ASAP7_75t_SL g1203 ( .A(n_1204), .B(n_1207), .C(n_1210), .Y(n_1203) );
AND4x1_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1215), .C(n_1216), .D(n_1217), .Y(n_1213) );
CKINVDCx20_ASAP7_75t_R g1219 ( .A(n_1220), .Y(n_1219) );
CKINVDCx20_ASAP7_75t_R g1220 ( .A(n_1221), .Y(n_1220) );
endmodule