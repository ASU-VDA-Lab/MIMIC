module fake_aes_8961_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
HB1xp67_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NAND2xp33_ASAP7_75t_L g4 ( .A(n_1), .B(n_0), .Y(n_4) );
OAI21x1_ASAP7_75t_SL g5 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_5) );
NAND2x1p5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_0), .Y(n_7) );
INVxp67_ASAP7_75t_SL g8 ( .A(n_6), .Y(n_8) );
OAI22xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_5), .B1(n_1), .B2(n_2), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_2), .Y(n_10) );
OAI211xp5_ASAP7_75t_SL g11 ( .A1(n_10), .A2(n_7), .B(n_2), .C(n_0), .Y(n_11) );
OA22x2_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_7), .B1(n_9), .B2(n_2), .Y(n_12) );
AOI21xp33_ASAP7_75t_SL g13 ( .A1(n_12), .A2(n_7), .B(n_6), .Y(n_13) );
endmodule