module fake_jpeg_4959_n_69 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_43;
wire n_37;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_38),
.B1(n_39),
.B2(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_54),
.Y(n_57)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_32),
.B1(n_42),
.B2(n_8),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_35),
.B(n_5),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_9),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_16),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_54),
.B1(n_50),
.B2(n_52),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_61),
.B(n_57),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_21),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_24),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_27),
.Y(n_69)
);


endmodule