module fake_jpeg_12660_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_1),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_59),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_63),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_48),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_20),
.C(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_75),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_46),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_5),
.B(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_10),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_44),
.B1(n_42),
.B2(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_51),
.B1(n_60),
.B2(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_49),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_83),
.C(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_88),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_81),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_68),
.B1(n_64),
.B2(n_70),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_15),
.B(n_17),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_47),
.B1(n_39),
.B2(n_6),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_52),
.C(n_47),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_2),
.B(n_5),
.C(n_6),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_21),
.B(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_66),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_98),
.B1(n_99),
.B2(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_98),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_97),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_36),
.B(n_84),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_104),
.C(n_92),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_91),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_106),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_116),
.C(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_113),
.B(n_111),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_111),
.C(n_110),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_99),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_94),
.Y(n_121)
);


endmodule