module fake_jpeg_1482_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_55;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx8_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_14),
.B(n_2),
.C(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_4),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_30),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_9),
.B(n_8),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_16),
.B(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_15),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_16),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_19),
.B1(n_8),
.B2(n_16),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_37),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_33),
.B(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_28),
.C(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_28),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_39),
.B(n_35),
.Y(n_47)
);

AOI21x1_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_48),
.B(n_41),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_39),
.B(n_33),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_46),
.C(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B(n_55),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_46),
.B(n_27),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_55),
.B(n_52),
.Y(n_58)
);

AOI221xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_57),
.B1(n_52),
.B2(n_53),
.C(n_34),
.Y(n_59)
);


endmodule