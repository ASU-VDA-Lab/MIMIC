module fake_jpeg_5436_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_31),
.Y(n_38)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_37),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_29),
.B1(n_36),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_62),
.B1(n_19),
.B2(n_22),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_56),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_21),
.B(n_23),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_66),
.B(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_53),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_29),
.B1(n_14),
.B2(n_22),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_22),
.B(n_17),
.C(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_28),
.B1(n_27),
.B2(n_16),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_50),
.B1(n_42),
.B2(n_20),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_44),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_49),
.CI(n_20),
.CON(n_76),
.SN(n_76)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_41),
.B1(n_44),
.B2(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_86),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_52),
.B1(n_26),
.B2(n_20),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_65),
.B1(n_55),
.B2(n_63),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_104),
.B(n_82),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_100),
.Y(n_113)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_106),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_65),
.B(n_64),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_116),
.B(n_119),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_115),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_79),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_112),
.C(n_118),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_74),
.C(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_56),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_104),
.C(n_93),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_94),
.C(n_105),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_105),
.A3(n_90),
.B1(n_106),
.B2(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_133),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_89),
.C(n_90),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_61),
.C(n_68),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_112),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_84),
.B1(n_66),
.B2(n_59),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_124),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_120),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_101),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_142),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_116),
.B1(n_111),
.B2(n_59),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_146),
.B1(n_129),
.B2(n_32),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_61),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_145),
.B(n_132),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_68),
.B(n_67),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_138),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_52),
.B1(n_32),
.B2(n_26),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_52),
.B1(n_32),
.B2(n_2),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_13),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_140),
.B(n_13),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_143),
.B(n_140),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_159),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_151),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_164),
.B(n_0),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_151),
.B1(n_147),
.B2(n_161),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_1),
.C(n_4),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_6),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_171),
.B(n_166),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_165),
.B(n_8),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_172),
.B(n_7),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_8),
.B(n_9),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_9),
.C(n_11),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_176),
.B(n_11),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_11),
.Y(n_180)
);


endmodule