module fake_jpeg_9666_n_63 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_11),
.B1(n_23),
.B2(n_22),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_29),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_1),
.C(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_44),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_25),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_48),
.C(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_30),
.B1(n_28),
.B2(n_13),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_49),
.B(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

AO21x2_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_30),
.B(n_4),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_54),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_5),
.C(n_6),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_7),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_45),
.C(n_49),
.Y(n_61)
);

OAI321xp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_49),
.A3(n_51),
.B1(n_20),
.B2(n_21),
.C(n_12),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_42),
.B1(n_14),
.B2(n_24),
.Y(n_63)
);


endmodule