module real_jpeg_11986_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_292;
wire n_288;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_30),
.B1(n_33),
.B2(n_54),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_79),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_79),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_30),
.B1(n_33),
.B2(n_79),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_74),
.B1(n_75),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_71),
.B(n_74),
.C(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_5),
.B(n_81),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_5),
.B(n_60),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_SL g211 ( 
.A1(n_5),
.A2(n_60),
.B(n_197),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_5),
.B(n_30),
.C(n_48),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_141),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_5),
.B(n_87),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_45),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_9),
.A2(n_30),
.B1(n_33),
.B2(n_45),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_9),
.A2(n_45),
.B1(n_74),
.B2(n_75),
.Y(n_289)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_74),
.B1(n_75),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_144),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_144),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_11),
.A2(n_30),
.B1(n_33),
.B2(n_144),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_74),
.B1(n_75),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_13),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_132),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_132),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_13),
.A2(n_30),
.B1(n_33),
.B2(n_132),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_14),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_14),
.A2(n_32),
.B1(n_74),
.B2(n_75),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_14),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_14),
.A2(n_32),
.B1(n_60),
.B2(n_61),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_15),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_15),
.A2(n_38),
.B1(n_60),
.B2(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_15),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_15),
.A2(n_38),
.B1(n_74),
.B2(n_75),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_275),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_133),
.B(n_274),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_19),
.B(n_111),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_83),
.B2(n_110),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_20),
.B(n_84),
.C(n_95),
.Y(n_277)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.C(n_68),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_22),
.A2(n_23),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_263)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_27),
.A2(n_35),
.B(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_28),
.A2(n_121),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_28),
.A2(n_34),
.B(n_159),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_28),
.A2(n_158),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_29),
.A2(n_123),
.B(n_158),
.Y(n_200)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_51)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_33),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_35),
.A2(n_36),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_35),
.A2(n_120),
.B(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_35),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_35),
.A2(n_36),
.B1(n_226),
.B2(n_234),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_36),
.B(n_37),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_36),
.B(n_141),
.Y(n_232)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_42),
.A2(n_51),
.B(n_92),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_44),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_SL g198 ( 
.A(n_43),
.B(n_57),
.C(n_61),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_44),
.A2(n_58),
.B(n_196),
.C(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_44),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_53),
.B(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_46),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_46),
.A2(n_52),
.B1(n_192),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_46),
.A2(n_52),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_46),
.A2(n_52),
.B1(n_213),
.B2(n_223),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_51),
.B(n_141),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_51),
.A2(n_151),
.B(n_152),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_52),
.B(n_93),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_68),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_59),
.B(n_63),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_56),
.A2(n_65),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_56),
.A2(n_65),
.B1(n_147),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_56),
.A2(n_65),
.B1(n_169),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_66)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_61),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_60),
.A2(n_72),
.B(n_141),
.Y(n_162)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_65),
.A2(n_148),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_65),
.A2(n_128),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_67),
.B(n_87),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_78),
.B(n_80),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_70),
.B1(n_78),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_69),
.A2(n_70),
.B1(n_131),
.B2(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_70),
.A2(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_81),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_95),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B(n_94),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_87),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_88),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_90),
.A2(n_151),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_94),
.B(n_279),
.CI(n_280),
.CON(n_278),
.SN(n_278)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_103),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g279 ( 
.A1(n_96),
.A2(n_97),
.B(n_105),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_102),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_109),
.B(n_139),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_117),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_116),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_117),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.C(n_129),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_118),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_124),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_265)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_268),
.B(n_273),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_181),
.B(n_259),
.C(n_267),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_170),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_136),
.B(n_170),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_154),
.C(n_163),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_149),
.C(n_153),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_155),
.B1(n_163),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_168),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_171),
.B(n_179),
.C(n_180),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_173),
.B(n_174),
.C(n_177),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_257),
.B(n_258),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_201),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_184),
.B(n_187),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_193),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_199),
.B1(n_200),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_214),
.B(n_256),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_212),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_250),
.B(n_255),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_240),
.B(n_249),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_229),
.B(n_239),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_221),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_238),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_245),
.C(n_248),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_254),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_266),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_292),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_278),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_278),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_288),
.B2(n_291),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);


endmodule