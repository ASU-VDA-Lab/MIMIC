module fake_netlist_5_729_n_2257 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2257);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2257;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_2248;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_315;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2044;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_158),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_48),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_129),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_8),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_41),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_212),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_92),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_120),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_61),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_27),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_77),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_119),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_35),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_165),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_18),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_193),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_104),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_91),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_125),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_68),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_150),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_23),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_80),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_67),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_114),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_68),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_1),
.Y(n_258)
);

BUFx8_ASAP7_75t_SL g259 ( 
.A(n_61),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_57),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_62),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_29),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_4),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_26),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_111),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_130),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_204),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_113),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_122),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_17),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_54),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_11),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_219),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_157),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_55),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_148),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_107),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_170),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_168),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_121),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_79),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_64),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_64),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_210),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_17),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_183),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_66),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_117),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_8),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_93),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_187),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_154),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_139),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_211),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_2),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_19),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_96),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_69),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_73),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_41),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_208),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_5),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_6),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_145),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_110),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_73),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_71),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_189),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_18),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_62),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_3),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_74),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_137),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_172),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_105),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_131),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_14),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_97),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_63),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_29),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_28),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_141),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_101),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_67),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_43),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_21),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_197),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_12),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_56),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_102),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_45),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_207),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_25),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_22),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_6),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_36),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_134),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_28),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_72),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_59),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_98),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_95),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_40),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_76),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_24),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_220),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_209),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_63),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_146),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_60),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_133),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_13),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_40),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_205),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_143),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_49),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_202),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_27),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_194),
.Y(n_365)
);

INVx4_ASAP7_75t_R g366 ( 
.A(n_82),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_37),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_159),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_185),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_109),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_87),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_2),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_106),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_83),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_51),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_88),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_45),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_80),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_116),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_181),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_78),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_196),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_66),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_21),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_37),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_153),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_74),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_100),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_54),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_55),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_25),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_16),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_51),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_53),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_180),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_84),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_3),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_15),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_58),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_57),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_152),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_5),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_155),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_24),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_59),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_200),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_13),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_216),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_72),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_188),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_88),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_144),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_169),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_162),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_84),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_164),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_26),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_56),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_123),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_214),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_179),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_174),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_126),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_77),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_79),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_76),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_43),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_30),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_140),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_177),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_167),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_128),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_86),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_176),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_201),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_20),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_0),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_49),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_78),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_22),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_46),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_7),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_115),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_225),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_267),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_260),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_259),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_268),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_299),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_300),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_403),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_384),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_232),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_234),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_299),
.B(n_0),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_235),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_351),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_421),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_236),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_229),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_229),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_302),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_240),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_360),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_233),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_242),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_427),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_286),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_228),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_238),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_233),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_286),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_286),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_360),
.Y(n_484)
);

CKINVDCx14_ASAP7_75t_R g485 ( 
.A(n_273),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_302),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_443),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_244),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_286),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_252),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_277),
.B(n_338),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_286),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_269),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_265),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_271),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_239),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_276),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_283),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_241),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_443),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_286),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_288),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_243),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_313),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_290),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_313),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_292),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_296),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_313),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_297),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_298),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_306),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_253),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_313),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_231),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_314),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_277),
.B(n_1),
.Y(n_517)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_239),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_338),
.B(n_4),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_313),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_313),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_387),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_387),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_387),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_320),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_321),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_387),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_231),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_273),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_324),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_387),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_328),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_269),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_247),
.B(n_7),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_387),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_343),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_389),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_347),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_389),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_273),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_389),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_389),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_348),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_251),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_251),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_389),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_352),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_254),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_263),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_353),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_419),
.B(n_9),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_355),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_361),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_439),
.Y(n_557)
);

CKINVDCx14_ASAP7_75t_R g558 ( 
.A(n_273),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_363),
.Y(n_559)
);

INVxp33_ASAP7_75t_L g560 ( 
.A(n_255),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_365),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_368),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_327),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_493),
.B(n_327),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_491),
.B(n_419),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_455),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_R g568 ( 
.A(n_485),
.B(n_369),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_478),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_445),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_460),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_450),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_533),
.B(n_327),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_478),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_457),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_515),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_515),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_534),
.B(n_422),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_459),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_482),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_483),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_483),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_534),
.B(n_422),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_463),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_470),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_489),
.B(n_439),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_515),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_476),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_475),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_528),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_489),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_488),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_528),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_492),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_492),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_528),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_501),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_504),
.Y(n_600)
);

BUFx8_ASAP7_75t_L g601 ( 
.A(n_540),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_504),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_506),
.B(n_247),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_464),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_477),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_490),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_509),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_494),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_486),
.B(n_439),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_495),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_509),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_497),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_491),
.B(n_370),
.Y(n_614)
);

OA21x2_ASAP7_75t_L g615 ( 
.A1(n_514),
.A2(n_521),
.B(n_520),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_553),
.B(n_514),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_520),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_R g618 ( 
.A(n_558),
.B(n_379),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_521),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_522),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_498),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_461),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_467),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_522),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_523),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_523),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_502),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_524),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_527),
.B(n_380),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_505),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_468),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_527),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_508),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_531),
.B(n_386),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_531),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_535),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_512),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_535),
.B(n_401),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_516),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_479),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_525),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_537),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_486),
.B(n_275),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_461),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_539),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_539),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_530),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_446),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_532),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_549),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_541),
.B(n_412),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_552),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_542),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_542),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_587),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_587),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_606),
.B(n_564),
.Y(n_662)
);

INVx5_ASAP7_75t_L g663 ( 
.A(n_651),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_615),
.Y(n_664)
);

INVx4_ASAP7_75t_SL g665 ( 
.A(n_604),
.Y(n_665)
);

INVx6_ASAP7_75t_L g666 ( 
.A(n_601),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_617),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_603),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_579),
.B(n_555),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_579),
.B(n_584),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_603),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_615),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_603),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_579),
.B(n_500),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_579),
.B(n_556),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_651),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_579),
.B(n_559),
.Y(n_677)
);

INVxp33_ASAP7_75t_L g678 ( 
.A(n_606),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_568),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_610),
.B(n_256),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_614),
.B(n_503),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_646),
.B(n_484),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_565),
.B(n_564),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_646),
.B(n_500),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_584),
.B(n_563),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_651),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_565),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_651),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_641),
.B(n_480),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_584),
.B(n_614),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_616),
.B(n_451),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_584),
.B(n_543),
.Y(n_692)
);

NAND3x1_ASAP7_75t_L g693 ( 
.A(n_566),
.B(n_458),
.C(n_517),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_615),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_604),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_615),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_566),
.A2(n_565),
.B1(n_573),
.B2(n_472),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_615),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_573),
.B(n_517),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_584),
.B(n_543),
.Y(n_700)
);

AND2x6_ASAP7_75t_L g701 ( 
.A(n_573),
.B(n_247),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_616),
.B(n_499),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_604),
.B(n_226),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_617),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_630),
.B(n_547),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_604),
.B(n_226),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_567),
.B(n_448),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_594),
.Y(n_708)
);

INVxp67_ASAP7_75t_SL g709 ( 
.A(n_630),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_569),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_641),
.B(n_513),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_590),
.B(n_550),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_569),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_574),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_574),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_617),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_622),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_635),
.B(n_639),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_635),
.B(n_247),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_575),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_575),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_570),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_639),
.B(n_547),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_624),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_645),
.B(n_519),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_655),
.B(n_280),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_655),
.B(n_227),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_576),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_581),
.Y(n_729)
);

INVx4_ASAP7_75t_SL g730 ( 
.A(n_581),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_582),
.B(n_227),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_582),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_590),
.B(n_551),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_583),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_571),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_594),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_592),
.B(n_231),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_592),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_595),
.B(n_231),
.Y(n_740)
);

INVx6_ASAP7_75t_L g741 ( 
.A(n_601),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_571),
.B(n_519),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_595),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_596),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_624),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_596),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_601),
.B(n_280),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_601),
.B(n_281),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_624),
.Y(n_750)
);

NAND2x1p5_ASAP7_75t_L g751 ( 
.A(n_598),
.B(n_295),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_598),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_599),
.A2(n_257),
.B1(n_289),
.B2(n_230),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_599),
.A2(n_257),
.B1(n_289),
.B2(n_230),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_600),
.B(n_231),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_600),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_629),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_602),
.A2(n_407),
.B1(n_359),
.B2(n_262),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_602),
.B(n_548),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_594),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_580),
.B(n_447),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_585),
.B(n_452),
.Y(n_762)
);

INVx5_ASAP7_75t_L g763 ( 
.A(n_577),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_SL g764 ( 
.A(n_601),
.B(n_487),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_629),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_572),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_568),
.B(n_529),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_608),
.B(n_548),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_622),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_629),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_577),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_608),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_612),
.A2(n_407),
.B1(n_359),
.B2(n_262),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_647),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_586),
.A2(n_510),
.B1(n_511),
.B2(n_507),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_612),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_618),
.B(n_529),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_619),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_619),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_620),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_620),
.B(n_237),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_625),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_625),
.B(n_554),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_647),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_618),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_605),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_626),
.B(n_554),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_626),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_628),
.B(n_237),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_589),
.B(n_518),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_628),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_593),
.B(n_546),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_633),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_648),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_633),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_607),
.B(n_560),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_636),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_636),
.B(n_231),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_609),
.B(n_281),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_637),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_637),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_643),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_643),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_648),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_605),
.B(n_474),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_644),
.Y(n_807)
);

BUFx10_ASAP7_75t_L g808 ( 
.A(n_611),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_644),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_613),
.B(n_526),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_621),
.B(n_282),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_649),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_649),
.B(n_248),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_658),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_658),
.Y(n_815)
);

AO22x2_ASAP7_75t_L g816 ( 
.A1(n_645),
.A2(n_258),
.B1(n_266),
.B2(n_255),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_709),
.B(n_627),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_691),
.A2(n_449),
.B(n_454),
.C(n_446),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_SL g819 ( 
.A1(n_691),
.A2(n_309),
.B(n_357),
.C(n_282),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_673),
.B(n_481),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_695),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_690),
.B(n_631),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_718),
.B(n_634),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_718),
.B(n_638),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_698),
.B(n_640),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_698),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_683),
.B(n_678),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_681),
.B(n_642),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_668),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_681),
.B(n_687),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_702),
.B(n_650),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_660),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_698),
.B(n_653),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_698),
.B(n_654),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_SL g836 ( 
.A1(n_725),
.A2(n_462),
.B1(n_453),
.B2(n_304),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_702),
.B(n_656),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_774),
.B(n_623),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_687),
.B(n_536),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_661),
.A2(n_454),
.B(n_456),
.C(n_449),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_670),
.A2(n_246),
.B(n_577),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_671),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_683),
.B(n_538),
.Y(n_843)
);

NOR2x1p5_ASAP7_75t_L g844 ( 
.A(n_679),
.B(n_261),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_693),
.A2(n_544),
.B1(n_561),
.B2(n_408),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_662),
.B(n_623),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_729),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_678),
.B(n_632),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_684),
.B(n_632),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_729),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_727),
.B(n_248),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_673),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_727),
.B(n_249),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_693),
.A2(n_420),
.B1(n_423),
.B2(n_414),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_735),
.Y(n_855)
);

NOR2xp67_ASAP7_75t_L g856 ( 
.A(n_679),
.B(n_496),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_727),
.B(n_249),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_735),
.B(n_250),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_699),
.A2(n_357),
.B1(n_373),
.B2(n_309),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_782),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_782),
.B(n_705),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_717),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_710),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_791),
.B(n_545),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_723),
.B(n_250),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_668),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_713),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_714),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_793),
.B(n_261),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_668),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_664),
.B(n_373),
.Y(n_871)
);

OAI221xp5_ASAP7_75t_L g872 ( 
.A1(n_697),
.A2(n_330),
.B1(n_378),
.B2(n_325),
.C(n_323),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_797),
.B(n_432),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_699),
.A2(n_272),
.B1(n_294),
.B2(n_284),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_664),
.B(n_429),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_667),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_715),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_786),
.B(n_557),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_699),
.B(n_272),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_733),
.B(n_264),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_664),
.B(n_429),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_699),
.B(n_284),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_672),
.B(n_431),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_703),
.B(n_294),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_672),
.A2(n_465),
.B(n_456),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_728),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_SL g887 ( 
.A(n_680),
.B(n_307),
.C(n_278),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_769),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_785),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_703),
.B(n_310),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_703),
.B(n_310),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_672),
.B(n_431),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_706),
.B(n_319),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_694),
.A2(n_301),
.B1(n_245),
.B2(n_364),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_706),
.B(n_319),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_670),
.B(n_322),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_736),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_706),
.B(n_322),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_733),
.B(n_270),
.Y(n_899)
);

AND2x2_ASAP7_75t_SL g900 ( 
.A(n_725),
.B(n_329),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_667),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_680),
.A2(n_382),
.B1(n_388),
.B2(n_395),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_711),
.B(n_279),
.C(n_274),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_720),
.B(n_329),
.Y(n_904)
);

INVxp33_ASAP7_75t_L g905 ( 
.A(n_682),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_732),
.B(n_333),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_734),
.B(n_333),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_694),
.B(n_465),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_739),
.B(n_336),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_774),
.B(n_666),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_704),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_743),
.B(n_336),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_744),
.Y(n_913)
);

AO22x1_ASAP7_75t_L g914 ( 
.A1(n_701),
.A2(n_334),
.B1(n_330),
.B2(n_325),
.Y(n_914)
);

NAND3xp33_ASAP7_75t_L g915 ( 
.A(n_711),
.B(n_293),
.C(n_285),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_SL g916 ( 
.A1(n_676),
.A2(n_406),
.B(n_382),
.C(n_388),
.Y(n_916)
);

INVx8_ASAP7_75t_L g917 ( 
.A(n_806),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_747),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_704),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_716),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_752),
.B(n_395),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_756),
.B(n_406),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_669),
.A2(n_677),
.B1(n_685),
.B2(n_675),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_726),
.A2(n_557),
.B(n_562),
.C(n_245),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_772),
.B(n_410),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_689),
.B(n_800),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_776),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_800),
.B(n_303),
.Y(n_928)
);

BUFx8_ASAP7_75t_L g929 ( 
.A(n_736),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_778),
.B(n_779),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_716),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_780),
.B(n_789),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_792),
.B(n_410),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_796),
.B(n_413),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_801),
.B(n_413),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_SL g936 ( 
.A(n_666),
.B(n_416),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_724),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_674),
.A2(n_430),
.B1(n_416),
.B2(n_434),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_712),
.B(n_312),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_802),
.B(n_430),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_804),
.B(n_434),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_807),
.B(n_435),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_724),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_742),
.B(n_312),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_694),
.B(n_696),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_809),
.B(n_435),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_745),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_812),
.B(n_444),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_696),
.B(n_444),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_696),
.B(n_652),
.Y(n_950)
);

AND2x6_ASAP7_75t_SL g951 ( 
.A(n_761),
.B(n_258),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_686),
.B(n_658),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_668),
.B(n_466),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_674),
.A2(n_466),
.B1(n_469),
.B2(n_473),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_688),
.B(n_657),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_721),
.B(n_657),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_721),
.B(n_657),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_811),
.B(n_308),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_721),
.B(n_652),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_721),
.B(n_652),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_811),
.B(n_742),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_794),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_751),
.B(n_311),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_751),
.A2(n_469),
.B1(n_471),
.B2(n_473),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_748),
.B(n_562),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_726),
.A2(n_471),
.B(n_287),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_806),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_761),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_701),
.A2(n_301),
.B1(n_287),
.B2(n_291),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_665),
.B(n_390),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_794),
.B(n_798),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_742),
.B(n_390),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_798),
.B(n_803),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_798),
.B(n_578),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_742),
.B(n_315),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_798),
.B(n_803),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_767),
.B(n_438),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_803),
.B(n_588),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_692),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_SL g980 ( 
.A1(n_722),
.A2(n_411),
.B1(n_394),
.B2(n_383),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_803),
.B(n_700),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_745),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_701),
.B(n_588),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_701),
.A2(n_266),
.B1(n_291),
.B2(n_305),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_746),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_701),
.B(n_588),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_719),
.A2(n_438),
.B(n_318),
.C(n_323),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_831),
.B(n_701),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_876),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_827),
.B(n_665),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_861),
.B(n_762),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_827),
.B(n_665),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_862),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_823),
.B(n_762),
.Y(n_994)
);

BUFx10_ASAP7_75t_L g995 ( 
.A(n_843),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_823),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_833),
.B(n_731),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_864),
.B(n_816),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_827),
.B(n_885),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_833),
.B(n_979),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_876),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_847),
.B(n_748),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_SL g1003 ( 
.A1(n_832),
.A2(n_346),
.B1(n_377),
.B2(n_810),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_901),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_827),
.B(n_728),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_901),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_880),
.B(n_731),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_985),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_911),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_911),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_862),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_821),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_880),
.B(n_731),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_888),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_863),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_867),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_850),
.B(n_749),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_868),
.Y(n_1018)
);

INVxp33_ASAP7_75t_SL g1019 ( 
.A(n_829),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_962),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_855),
.B(n_749),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_848),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_830),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_985),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_830),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_872),
.A2(n_813),
.B(n_781),
.C(n_790),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_962),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_962),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_919),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_830),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_899),
.B(n_781),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_962),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_899),
.B(n_781),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_817),
.B(n_790),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_828),
.B(n_816),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_888),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_877),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_968),
.B(n_810),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_923),
.A2(n_719),
.B1(n_777),
.B2(n_786),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_900),
.A2(n_816),
.B1(n_790),
.B2(n_813),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_SL g1041 ( 
.A(n_832),
.B(n_775),
.C(n_766),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_860),
.B(n_813),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_897),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_830),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_837),
.B(n_783),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_846),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_900),
.B(n_806),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_852),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_866),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_913),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_837),
.B(n_806),
.C(n_787),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_829),
.B(n_764),
.C(n_754),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_838),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_852),
.B(n_707),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_824),
.B(n_728),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_838),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_926),
.B(n_783),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_918),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_838),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_820),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_917),
.B(n_666),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_926),
.B(n_783),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_886),
.B(n_741),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_825),
.B(n_826),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_866),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_919),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_887),
.B(n_741),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_939),
.B(n_808),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_927),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_894),
.B(n_795),
.Y(n_1070)
);

BUFx12f_ASAP7_75t_L g1071 ( 
.A(n_889),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_R g1072 ( 
.A(n_889),
.B(n_741),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_842),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_894),
.B(n_795),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_930),
.B(n_795),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_920),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_932),
.B(n_760),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_822),
.B(n_760),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_920),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_869),
.B(n_808),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_910),
.B(n_730),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_929),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_910),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_839),
.B(n_808),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_822),
.B(n_760),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_SL g1086 ( 
.A(n_980),
.B(n_317),
.C(n_316),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_931),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_851),
.B(n_746),
.Y(n_1088)
);

BUFx4f_ASAP7_75t_L g1089 ( 
.A(n_910),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_820),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_870),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_931),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_SL g1093 ( 
.A(n_967),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_970),
.B(n_730),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_853),
.B(n_746),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_849),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_977),
.B(n_753),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_929),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_857),
.B(n_928),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_970),
.B(n_730),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_870),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_937),
.Y(n_1102)
);

NAND2x1_ASAP7_75t_L g1103 ( 
.A(n_937),
.B(n_771),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_943),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_943),
.Y(n_1105)
);

AO22x1_ASAP7_75t_L g1106 ( 
.A1(n_961),
.A2(n_331),
.B1(n_326),
.B2(n_332),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_928),
.B(n_663),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_958),
.B(n_663),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_971),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_947),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_973),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_878),
.B(n_90),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_917),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_947),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_917),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_SL g1116 ( 
.A(n_843),
.B(n_839),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_982),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_958),
.B(n_663),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_982),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_950),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_SL g1121 ( 
.A(n_856),
.B(n_335),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_945),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_952),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_945),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_966),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_896),
.Y(n_1126)
);

INVx6_ASAP7_75t_L g1127 ( 
.A(n_844),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_951),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_966),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_976),
.Y(n_1130)
);

OR2x2_ASAP7_75t_SL g1131 ( 
.A(n_903),
.B(n_305),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_983),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_836),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_955),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_986),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_884),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_961),
.B(n_758),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_879),
.B(n_663),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_882),
.B(n_858),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_956),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_905),
.B(n_337),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_975),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_845),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_826),
.A2(n_815),
.B1(n_814),
.B2(n_759),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_944),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_834),
.A2(n_768),
.B1(n_784),
.B2(n_788),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_896),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_972),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_890),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_965),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_891),
.Y(n_1151)
);

BUFx4_ASAP7_75t_SL g1152 ( 
.A(n_915),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_834),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_975),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_965),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_957),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_893),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_949),
.B(n_773),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_895),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_835),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_835),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_969),
.B(n_663),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_898),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_914),
.Y(n_1164)
);

BUFx8_ASAP7_75t_SL g1165 ( 
.A(n_904),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_859),
.A2(n_805),
.B1(n_757),
.B2(n_750),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_984),
.B(n_750),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_959),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_865),
.B(n_757),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_906),
.B(n_339),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_969),
.B(n_765),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_981),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_960),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_SL g1174 ( 
.A(n_873),
.B(n_341),
.C(n_340),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_907),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_938),
.B(n_94),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_909),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_912),
.Y(n_1178)
);

INVx5_ASAP7_75t_L g1179 ( 
.A(n_908),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_953),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1116),
.A2(n_963),
.B1(n_854),
.B2(n_902),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_999),
.A2(n_908),
.B(n_875),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1019),
.A2(n_984),
.B1(n_883),
.B2(n_875),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1007),
.A2(n_881),
.B(n_871),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_993),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1125),
.A2(n_881),
.B(n_871),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1038),
.B(n_987),
.Y(n_1187)
);

AO21x1_ASAP7_75t_L g1188 ( 
.A1(n_1064),
.A2(n_874),
.B(n_883),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1013),
.A2(n_892),
.B(n_818),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1019),
.A2(n_892),
.B1(n_964),
.B2(n_841),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_991),
.B(n_921),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1096),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_993),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1125),
.A2(n_978),
.B(n_974),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1135),
.A2(n_953),
.B(n_924),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_988),
.A2(n_1112),
.B(n_1017),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1022),
.A2(n_925),
.B(n_922),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_998),
.B(n_1068),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_999),
.A2(n_840),
.B(n_954),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1075),
.A2(n_934),
.B(n_933),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_998),
.B(n_935),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_994),
.B(n_940),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1129),
.A2(n_942),
.B(n_941),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1099),
.B(n_948),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1031),
.A2(n_946),
.B(n_819),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1175),
.B(n_765),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_996),
.Y(n_1207)
);

OAI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1121),
.A2(n_349),
.B(n_344),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1129),
.A2(n_805),
.B(n_770),
.Y(n_1209)
);

AOI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1133),
.A2(n_819),
.B(n_936),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1077),
.A2(n_799),
.B(n_738),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_SL g1212 ( 
.A1(n_1000),
.A2(n_334),
.B(n_318),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1012),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1033),
.B(n_770),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1026),
.A2(n_400),
.A3(n_345),
.B(n_358),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_989),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1064),
.A2(n_597),
.B(n_591),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1057),
.A2(n_597),
.B(n_591),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1135),
.A2(n_771),
.B(n_591),
.Y(n_1220)
);

NOR2x1_ASAP7_75t_SL g1221 ( 
.A(n_1061),
.B(n_708),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1101),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_L g1223 ( 
.A(n_1124),
.B(n_740),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_SL g1224 ( 
.A1(n_1112),
.A2(n_916),
.B(n_366),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1070),
.A2(n_799),
.B(n_738),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1045),
.B(n_771),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1074),
.A2(n_708),
.B(n_737),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1176),
.A2(n_397),
.B(n_345),
.C(n_358),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1122),
.A2(n_916),
.B(n_755),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_SL g1230 ( 
.A1(n_1126),
.A2(n_342),
.B(n_364),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1122),
.A2(n_755),
.B(n_740),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1011),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1153),
.B(n_1160),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_989),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1130),
.A2(n_1147),
.B(n_1120),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1130),
.A2(n_597),
.B(n_409),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1163),
.B(n_350),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1101),
.Y(n_1238)
);

CKINVDCx14_ASAP7_75t_R g1239 ( 
.A(n_1072),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1078),
.A2(n_1085),
.B(n_1062),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1068),
.B(n_354),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_L g1242 ( 
.A(n_1071),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1026),
.A2(n_399),
.A3(n_426),
.B(n_342),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1003),
.B(n_356),
.C(n_362),
.Y(n_1244)
);

CKINVDCx6p67_ASAP7_75t_R g1245 ( 
.A(n_1071),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1171),
.A2(n_755),
.B(n_740),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1034),
.A2(n_708),
.B(n_737),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1120),
.A2(n_708),
.B(n_737),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1142),
.A2(n_740),
.B1(n_755),
.B2(n_404),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1139),
.A2(n_755),
.B(n_740),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1080),
.B(n_367),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1153),
.B(n_708),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1176),
.A2(n_400),
.B(n_371),
.C(n_440),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1107),
.A2(n_737),
.B(n_763),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1154),
.B(n_372),
.Y(n_1255)
);

BUFx4_ASAP7_75t_SL g1256 ( 
.A(n_1014),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1136),
.B(n_374),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1061),
.B(n_371),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1108),
.A2(n_418),
.B(n_392),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1046),
.B(n_375),
.Y(n_1260)
);

BUFx2_ASAP7_75t_SL g1261 ( 
.A(n_1014),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1130),
.A2(n_378),
.B(n_392),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1149),
.B(n_1151),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1159),
.B(n_376),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1118),
.A2(n_737),
.B(n_763),
.Y(n_1265)
);

NAND2x1p5_ASAP7_75t_L g1266 ( 
.A(n_1101),
.B(n_763),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1147),
.A2(n_393),
.B(n_397),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1180),
.A2(n_424),
.A3(n_393),
.B(n_399),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1147),
.A2(n_409),
.B(n_440),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1145),
.B(n_381),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1133),
.B(n_385),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1158),
.A2(n_755),
.B(n_740),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1087),
.A2(n_418),
.B(n_426),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_997),
.A2(n_763),
.B(n_424),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1087),
.A2(n_1105),
.B(n_1065),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1087),
.A2(n_132),
.B(n_224),
.Y(n_1276)
);

NOR2x1_ASAP7_75t_SL g1277 ( 
.A(n_1061),
.B(n_763),
.Y(n_1277)
);

NOR2xp67_ASAP7_75t_L g1278 ( 
.A(n_1051),
.B(n_99),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1176),
.A2(n_442),
.B(n_441),
.C(n_437),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1015),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1080),
.B(n_391),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1088),
.A2(n_118),
.B(n_223),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1146),
.A2(n_436),
.B(n_433),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1105),
.A2(n_1065),
.B(n_1049),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1041),
.B(n_396),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1105),
.A2(n_103),
.B(n_108),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1040),
.A2(n_428),
.B1(n_425),
.B2(n_417),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1180),
.A2(n_366),
.A3(n_10),
.B(n_12),
.Y(n_1288)
);

INVx5_ASAP7_75t_L g1289 ( 
.A(n_1020),
.Y(n_1289)
);

AOI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1138),
.A2(n_1169),
.B(n_1095),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1126),
.A2(n_178),
.B(n_124),
.Y(n_1291)
);

AO32x2_ASAP7_75t_L g1292 ( 
.A1(n_1164),
.A2(n_9),
.A3(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_1292)
);

BUFx12f_ASAP7_75t_L g1293 ( 
.A(n_1098),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1011),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1049),
.A2(n_222),
.B(n_218),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1049),
.A2(n_217),
.B(n_213),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1055),
.B(n_415),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1065),
.A2(n_206),
.B(n_199),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1123),
.B(n_1134),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1158),
.A2(n_405),
.B(n_402),
.Y(n_1300)
);

O2A1O1Ixp5_ASAP7_75t_L g1301 ( 
.A1(n_1002),
.A2(n_163),
.B(n_198),
.C(n_195),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1091),
.A2(n_160),
.B(n_192),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1137),
.A2(n_398),
.B(n_19),
.C(n_20),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_SL g1304 ( 
.A(n_1084),
.B(n_16),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1091),
.A2(n_186),
.B(n_184),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1036),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1076),
.A2(n_182),
.B(n_173),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1001),
.A2(n_171),
.B(n_166),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1020),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1143),
.B(n_23),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1001),
.A2(n_161),
.B(n_156),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1143),
.A2(n_30),
.B(n_31),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1157),
.B(n_31),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1016),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1091),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1140),
.A2(n_151),
.B(n_149),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1091),
.A2(n_147),
.B(n_142),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1018),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1157),
.B(n_32),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1091),
.A2(n_135),
.B(n_127),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1140),
.A2(n_112),
.B(n_33),
.Y(n_1321)
);

NAND2x1_ASAP7_75t_L g1322 ( 
.A(n_1032),
.B(n_32),
.Y(n_1322)
);

NAND2xp33_ASAP7_75t_SL g1323 ( 
.A(n_1063),
.B(n_1174),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1137),
.B(n_33),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1156),
.A2(n_34),
.B(n_36),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1035),
.B(n_34),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1035),
.B(n_38),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1004),
.A2(n_38),
.B(n_39),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1097),
.B(n_39),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1156),
.A2(n_42),
.B(n_44),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_SL g1331 ( 
.A1(n_1039),
.A2(n_1024),
.B(n_1008),
.C(n_1027),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1037),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1097),
.B(n_42),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1004),
.A2(n_1066),
.B(n_1029),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1006),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1153),
.B(n_44),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1061),
.A2(n_47),
.B(n_50),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1168),
.A2(n_47),
.B(n_50),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1168),
.A2(n_52),
.B(n_53),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1167),
.A2(n_52),
.B(n_58),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1006),
.A2(n_60),
.B(n_65),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1167),
.A2(n_65),
.B(n_69),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1124),
.A2(n_70),
.B(n_71),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1060),
.B(n_70),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1172),
.B(n_75),
.Y(n_1345)
);

CKINVDCx11_ASAP7_75t_R g1346 ( 
.A(n_1242),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1240),
.A2(n_1124),
.B(n_1179),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1216),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1209),
.A2(n_1166),
.B(n_1103),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1213),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1185),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1209),
.A2(n_1144),
.B(n_1066),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1196),
.A2(n_1029),
.B(n_1079),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1271),
.B(n_995),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1193),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1280),
.Y(n_1356)
);

OAI222xp33_ASAP7_75t_L g1357 ( 
.A1(n_1310),
.A2(n_1047),
.B1(n_1128),
.B2(n_1164),
.C1(n_1059),
.C2(n_1056),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1310),
.A2(n_1047),
.B1(n_995),
.B2(n_1128),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1235),
.A2(n_1220),
.B(n_1236),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_SL g1360 ( 
.A1(n_1188),
.A2(n_1180),
.B(n_1164),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1220),
.A2(n_1110),
.B(n_1104),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1271),
.B(n_995),
.Y(n_1362)
);

CKINVDCx16_ASAP7_75t_R g1363 ( 
.A(n_1242),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1236),
.A2(n_1079),
.B(n_1010),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_SL g1365 ( 
.A(n_1293),
.B(n_1082),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1233),
.B(n_1153),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1232),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1314),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1285),
.A2(n_1052),
.B1(n_1106),
.B2(n_1086),
.C(n_1141),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1297),
.A2(n_1148),
.B1(n_1090),
.B2(n_1127),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1234),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1335),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1233),
.B(n_1124),
.Y(n_1373)
);

BUFx8_ASAP7_75t_L g1374 ( 
.A(n_1293),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1275),
.A2(n_1009),
.B(n_1010),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1244),
.A2(n_1128),
.B1(n_1043),
.B2(n_1036),
.Y(n_1376)
);

OAI222xp33_ASAP7_75t_L g1377 ( 
.A1(n_1181),
.A2(n_1324),
.B1(n_1297),
.B2(n_1287),
.C1(n_1336),
.C2(n_1218),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_SL g1378 ( 
.A1(n_1228),
.A2(n_1005),
.B(n_1102),
.C(n_1117),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1205),
.A2(n_1114),
.B(n_1092),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1303),
.A2(n_1150),
.A3(n_1009),
.B(n_1058),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1294),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1256),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1290),
.A2(n_1150),
.B(n_1162),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1200),
.A2(n_1124),
.B(n_1179),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1318),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1335),
.Y(n_1386)
);

AND2x6_ASAP7_75t_L g1387 ( 
.A(n_1222),
.B(n_1153),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1275),
.A2(n_1008),
.B(n_1024),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1332),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1284),
.A2(n_1194),
.B(n_1334),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1207),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1198),
.B(n_1172),
.Y(n_1392)
);

INVx3_ASAP7_75t_SL g1393 ( 
.A(n_1245),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1334),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1285),
.A2(n_1021),
.B1(n_1002),
.B2(n_1017),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1192),
.Y(n_1396)
);

AOI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1214),
.A2(n_1162),
.B(n_1002),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1284),
.A2(n_1008),
.B(n_1024),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1183),
.A2(n_1017),
.B(n_1021),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1194),
.A2(n_1027),
.B(n_1028),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1273),
.Y(n_1401)
);

OAI211xp5_ASAP7_75t_L g1402 ( 
.A1(n_1312),
.A2(n_1342),
.B(n_1340),
.C(n_1300),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1315),
.Y(n_1403)
);

AND2x6_ASAP7_75t_L g1404 ( 
.A(n_1222),
.B(n_1161),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1203),
.A2(n_1073),
.B(n_1050),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1191),
.B(n_1172),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1299),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1186),
.A2(n_1203),
.B(n_1195),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1263),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1184),
.A2(n_1179),
.B(n_1119),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1273),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1303),
.A2(n_1069),
.A3(n_1032),
.B(n_1059),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1202),
.A2(n_1089),
.B1(n_1179),
.B2(n_1155),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1204),
.B(n_1172),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1217),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1262),
.A2(n_1021),
.B(n_1112),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1186),
.A2(n_1028),
.B(n_990),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1331),
.A2(n_1170),
.B(n_1067),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1206),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1306),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1201),
.B(n_1054),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1187),
.B(n_1042),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1255),
.A2(n_1128),
.B1(n_1056),
.B2(n_1148),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1289),
.B(n_1160),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1329),
.B(n_1042),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_R g1426 ( 
.A(n_1239),
.B(n_1082),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1268),
.Y(n_1427)
);

AO31x2_ASAP7_75t_L g1428 ( 
.A1(n_1228),
.A2(n_1032),
.A3(n_1160),
.B(n_1161),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1268),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1224),
.A2(n_992),
.B(n_990),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1262),
.A2(n_1005),
.B(n_992),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1315),
.B(n_1115),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1326),
.B(n_1161),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1333),
.B(n_1054),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1257),
.B(n_1054),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1309),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1189),
.A2(n_1042),
.B(n_1160),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1264),
.B(n_1111),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1214),
.A2(n_1161),
.B(n_1160),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_L g1440 ( 
.A(n_1255),
.B(n_1128),
.C(n_1053),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1217),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1217),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1182),
.A2(n_1161),
.B(n_1119),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1260),
.A2(n_1043),
.B1(n_1089),
.B2(n_1113),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1345),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1313),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1319),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1309),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1308),
.A2(n_1311),
.B(n_1276),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1253),
.B(n_1111),
.Y(n_1450)
);

BUFx8_ASAP7_75t_L g1451 ( 
.A(n_1292),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1308),
.A2(n_1119),
.B(n_1179),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1327),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1311),
.A2(n_1119),
.B(n_1132),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1276),
.A2(n_1119),
.B(n_1132),
.Y(n_1455)
);

AOI221x1_ASAP7_75t_L g1456 ( 
.A1(n_1325),
.A2(n_1173),
.B1(n_1109),
.B2(n_1111),
.C(n_1132),
.Y(n_1456)
);

AO31x2_ASAP7_75t_L g1457 ( 
.A1(n_1253),
.A2(n_1131),
.A3(n_1173),
.B(n_1132),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1199),
.A2(n_1155),
.B(n_1089),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1208),
.A2(n_1127),
.B1(n_1093),
.B2(n_1173),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1215),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1270),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1286),
.A2(n_1298),
.B(n_1295),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1261),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1286),
.A2(n_1173),
.B(n_1109),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1241),
.B(n_1109),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1212),
.A2(n_1131),
.B(n_1093),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_SL g1467 ( 
.A1(n_1331),
.A2(n_1152),
.B(n_1111),
.C(n_1109),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1215),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1267),
.A2(n_1044),
.B(n_1020),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1215),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1309),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1309),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1258),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1267),
.A2(n_1044),
.B(n_1020),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1251),
.B(n_1048),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1190),
.A2(n_1100),
.B(n_1094),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1279),
.B(n_1048),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1279),
.A2(n_1100),
.B(n_1094),
.Y(n_1478)
);

AOI21xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1237),
.A2(n_1113),
.B(n_1165),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1269),
.A2(n_1044),
.B(n_1020),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1243),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1330),
.A2(n_1093),
.B1(n_1083),
.B2(n_1115),
.C(n_1165),
.Y(n_1482)
);

AND2x6_ASAP7_75t_L g1483 ( 
.A(n_1238),
.B(n_1081),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1243),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1328),
.A2(n_1341),
.B(n_1225),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1269),
.A2(n_1044),
.B(n_1023),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1281),
.A2(n_1127),
.B1(n_1083),
.B2(n_1098),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1344),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1243),
.B(n_1100),
.Y(n_1489)
);

OAI22x1_ASAP7_75t_L g1490 ( 
.A1(n_1336),
.A2(n_1081),
.B1(n_1094),
.B2(n_1127),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1296),
.A2(n_1044),
.B(n_1030),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1289),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1197),
.B(n_1048),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1243),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1230),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1289),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1272),
.A2(n_1081),
.B(n_1048),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1304),
.A2(n_1323),
.B1(n_1339),
.B2(n_1338),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1274),
.A2(n_1030),
.B(n_1025),
.Y(n_1499)
);

AND2x4_ASAP7_75t_SL g1500 ( 
.A(n_1238),
.B(n_1258),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1211),
.A2(n_1030),
.B(n_1025),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1343),
.A2(n_75),
.B(n_81),
.C(n_82),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1283),
.B(n_1030),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1328),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1239),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1323),
.B(n_1025),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1296),
.A2(n_1248),
.B(n_1265),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1254),
.A2(n_1025),
.B(n_1023),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1258),
.B(n_1023),
.Y(n_1509)
);

AO31x2_ASAP7_75t_L g1510 ( 
.A1(n_1226),
.A2(n_1023),
.A3(n_83),
.B(n_85),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1341),
.A2(n_81),
.B(n_85),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1304),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1229),
.A2(n_86),
.B(n_87),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1259),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1288),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1283),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1252),
.A2(n_89),
.B(n_1250),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1227),
.A2(n_89),
.B(n_1307),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1420),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1407),
.B(n_1283),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1409),
.A2(n_1278),
.B1(n_1316),
.B2(n_1322),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1432),
.B(n_1289),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1369),
.A2(n_1210),
.B1(n_1321),
.B2(n_1252),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1420),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1453),
.B(n_1288),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1350),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1432),
.B(n_1221),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1348),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1451),
.A2(n_1292),
.B1(n_1337),
.B2(n_1223),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1355),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1346),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1414),
.B(n_1288),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1432),
.B(n_1277),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1392),
.B(n_1292),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1348),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1355),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1402),
.A2(n_1292),
.B1(n_1246),
.B2(n_1231),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1498),
.A2(n_1301),
.B(n_1282),
.C(n_1291),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1367),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1403),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1509),
.B(n_1320),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1356),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1346),
.Y(n_1543)
);

BUFx4f_ASAP7_75t_SL g1544 ( 
.A(n_1374),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1437),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1403),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1381),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1422),
.B(n_1317),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1368),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1512),
.A2(n_1249),
.B1(n_1266),
.B2(n_1302),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1509),
.B(n_1305),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1512),
.A2(n_1247),
.B1(n_1266),
.B2(n_1219),
.Y(n_1552)
);

CKINVDCx6p67_ASAP7_75t_R g1553 ( 
.A(n_1393),
.Y(n_1553)
);

AOI21xp33_ASAP7_75t_L g1554 ( 
.A1(n_1399),
.A2(n_1219),
.B(n_1223),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1422),
.B(n_1219),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1492),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1488),
.B(n_1425),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1425),
.B(n_1354),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1362),
.B(n_1445),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1395),
.A2(n_1414),
.B1(n_1451),
.B2(n_1358),
.Y(n_1560)
);

OR2x6_ASAP7_75t_SL g1561 ( 
.A(n_1505),
.B(n_1440),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1451),
.A2(n_1406),
.B1(n_1446),
.B2(n_1447),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1437),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1426),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1483),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1513),
.A2(n_1389),
.B1(n_1385),
.B2(n_1391),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1351),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1513),
.A2(n_1434),
.B1(n_1423),
.B2(n_1482),
.Y(n_1568)
);

INVx4_ASAP7_75t_SL g1569 ( 
.A(n_1387),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1437),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1513),
.A2(n_1517),
.B1(n_1473),
.B2(n_1357),
.Y(n_1571)
);

INVx4_ASAP7_75t_SL g1572 ( 
.A(n_1387),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1374),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1421),
.A2(n_1487),
.B1(n_1370),
.B2(n_1419),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1461),
.A2(n_1435),
.B1(n_1490),
.B2(n_1438),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1502),
.B(n_1459),
.C(n_1458),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_SL g1577 ( 
.A(n_1509),
.Y(n_1577)
);

AO31x2_ASAP7_75t_L g1578 ( 
.A1(n_1504),
.A2(n_1515),
.A3(n_1468),
.B(n_1460),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1433),
.B(n_1493),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1473),
.A2(n_1365),
.B1(n_1476),
.B2(n_1374),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1452),
.A2(n_1454),
.B(n_1359),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1492),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1351),
.B(n_1465),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1377),
.A2(n_1456),
.B(n_1384),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1418),
.A2(n_1511),
.B1(n_1360),
.B2(n_1478),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1418),
.A2(n_1511),
.B1(n_1360),
.B2(n_1363),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1371),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_SL g1588 ( 
.A1(n_1466),
.A2(n_1450),
.B(n_1497),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_SL g1589 ( 
.A(n_1475),
.B(n_1433),
.C(n_1479),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1372),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1386),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1386),
.B(n_1380),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1405),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1500),
.B(n_1463),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1496),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1366),
.B(n_1490),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1477),
.A2(n_1444),
.B1(n_1466),
.B2(n_1495),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1452),
.A2(n_1454),
.B(n_1359),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1405),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_R g1600 ( 
.A(n_1505),
.B(n_1489),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1382),
.Y(n_1601)
);

AND2x6_ASAP7_75t_SL g1602 ( 
.A(n_1506),
.B(n_1393),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1477),
.A2(n_1418),
.B1(n_1489),
.B2(n_1376),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1396),
.B(n_1366),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1413),
.A2(n_1500),
.B1(n_1467),
.B2(n_1366),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1366),
.A2(n_1424),
.B1(n_1410),
.B2(n_1373),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1427),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1483),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1436),
.B(n_1448),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1449),
.A2(n_1455),
.B(n_1408),
.Y(n_1610)
);

CKINVDCx11_ASAP7_75t_R g1611 ( 
.A(n_1436),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1429),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1448),
.B(n_1471),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_SL g1614 ( 
.A(n_1496),
.B(n_1397),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1503),
.A2(n_1516),
.B1(n_1514),
.B2(n_1387),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1457),
.B(n_1471),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1353),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1503),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1483),
.B(n_1472),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1467),
.A2(n_1404),
.B1(n_1387),
.B2(n_1483),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1380),
.B(n_1456),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1353),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1472),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1387),
.A2(n_1404),
.B1(n_1494),
.B2(n_1481),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1511),
.A2(n_1404),
.B1(n_1387),
.B2(n_1416),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1424),
.A2(n_1373),
.B1(n_1484),
.B2(n_1460),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1457),
.B(n_1412),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1483),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1424),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1483),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1404),
.A2(n_1378),
.B1(n_1373),
.B2(n_1416),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1470),
.A2(n_1416),
.B1(n_1347),
.B2(n_1397),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1379),
.A2(n_1504),
.B1(n_1383),
.B2(n_1501),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1404),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1439),
.B(n_1383),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1404),
.A2(n_1431),
.B1(n_1401),
.B2(n_1411),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1412),
.A2(n_1379),
.B1(n_1443),
.B2(n_1380),
.Y(n_1637)
);

OAI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1379),
.A2(n_1411),
.B1(n_1401),
.B2(n_1439),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1510),
.Y(n_1639)
);

NAND2xp33_ASAP7_75t_R g1640 ( 
.A(n_1431),
.B(n_1485),
.Y(n_1640)
);

NAND2xp33_ASAP7_75t_R g1641 ( 
.A(n_1431),
.B(n_1485),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_R g1642 ( 
.A(n_1485),
.B(n_1430),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1510),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1457),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1457),
.Y(n_1645)
);

OAI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1394),
.A2(n_1499),
.B1(n_1415),
.B2(n_1442),
.Y(n_1646)
);

INVx4_ASAP7_75t_SL g1647 ( 
.A(n_1457),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1510),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1378),
.A2(n_1412),
.B1(n_1380),
.B2(n_1394),
.C(n_1415),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1510),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1412),
.A2(n_1443),
.B1(n_1380),
.B2(n_1518),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1428),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1441),
.A2(n_1442),
.B1(n_1412),
.B2(n_1428),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1430),
.A2(n_1518),
.B1(n_1400),
.B2(n_1398),
.Y(n_1654)
);

AO32x2_ASAP7_75t_L g1655 ( 
.A1(n_1510),
.A2(n_1428),
.A3(n_1408),
.B1(n_1390),
.B2(n_1449),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1428),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1441),
.A2(n_1428),
.B1(n_1352),
.B2(n_1464),
.C(n_1364),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1398),
.B(n_1352),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1375),
.B(n_1361),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1417),
.B(n_1508),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1361),
.B(n_1388),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1388),
.B(n_1364),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1400),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1417),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1464),
.A2(n_1508),
.B1(n_1455),
.B2(n_1486),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1486),
.A2(n_1491),
.B1(n_1474),
.B2(n_1469),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1349),
.B(n_1390),
.Y(n_1667)
);

AO31x2_ASAP7_75t_L g1668 ( 
.A1(n_1507),
.A2(n_1462),
.A3(n_1469),
.B(n_1474),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1480),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1462),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1349),
.A2(n_1019),
.B1(n_832),
.B2(n_837),
.Y(n_1671)
);

CKINVDCx6p67_ASAP7_75t_R g1672 ( 
.A(n_1507),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1346),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1369),
.A2(n_1019),
.B1(n_832),
.B2(n_837),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1381),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1381),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1432),
.B(n_1509),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1346),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1492),
.Y(n_1679)
);

A2O1A1Ixp33_ASAP7_75t_SL g1680 ( 
.A1(n_1354),
.A2(n_829),
.B(n_837),
.C(n_832),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1402),
.A2(n_1019),
.B1(n_837),
.B2(n_832),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1392),
.B(n_1198),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1350),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1407),
.B(n_1324),
.Y(n_1684)
);

NOR2x1_ASAP7_75t_SL g1685 ( 
.A(n_1366),
.B(n_1061),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1381),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1420),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1350),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1407),
.B(n_1409),
.Y(n_1689)
);

CKINVDCx11_ASAP7_75t_R g1690 ( 
.A(n_1346),
.Y(n_1690)
);

OAI211xp5_ASAP7_75t_L g1691 ( 
.A1(n_1674),
.A2(n_1680),
.B(n_1681),
.C(n_1671),
.Y(n_1691)
);

OR2x6_ASAP7_75t_L g1692 ( 
.A(n_1596),
.B(n_1634),
.Y(n_1692)
);

OAI211xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1681),
.A2(n_1575),
.B(n_1586),
.C(n_1597),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1576),
.A2(n_1580),
.B1(n_1571),
.B2(n_1684),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1560),
.A2(n_1689),
.B1(n_1600),
.B2(n_1574),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1538),
.A2(n_1521),
.B(n_1584),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1580),
.A2(n_1571),
.B1(n_1529),
.B2(n_1559),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1574),
.A2(n_1560),
.B1(n_1682),
.B2(n_1568),
.Y(n_1698)
);

AOI222xp33_ASAP7_75t_L g1699 ( 
.A1(n_1562),
.A2(n_1568),
.B1(n_1544),
.B2(n_1537),
.C1(n_1689),
.C2(n_1579),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1526),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1613),
.B(n_1583),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1589),
.A2(n_1541),
.B1(n_1551),
.B2(n_1548),
.Y(n_1702)
);

OAI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1562),
.A2(n_1561),
.B1(n_1604),
.B2(n_1579),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1589),
.A2(n_1529),
.B1(n_1537),
.B2(n_1523),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1547),
.A2(n_1675),
.B1(n_1676),
.B2(n_1686),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1623),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1603),
.A2(n_1605),
.B1(n_1628),
.B2(n_1630),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1556),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1567),
.A2(n_1530),
.B1(n_1536),
.B2(n_1539),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1521),
.A2(n_1584),
.B1(n_1566),
.B2(n_1520),
.C(n_1588),
.Y(n_1710)
);

AOI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1520),
.A2(n_1525),
.B(n_1550),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1586),
.A2(n_1550),
.B1(n_1601),
.B2(n_1687),
.C(n_1585),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1542),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1541),
.A2(n_1551),
.B1(n_1544),
.B2(n_1683),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1624),
.A2(n_1620),
.B1(n_1615),
.B2(n_1596),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1549),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1688),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1566),
.A2(n_1585),
.B1(n_1525),
.B2(n_1532),
.C(n_1639),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1610),
.A2(n_1598),
.B(n_1581),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1690),
.A2(n_1577),
.B1(n_1611),
.B2(n_1677),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1577),
.A2(n_1594),
.B1(n_1532),
.B2(n_1543),
.Y(n_1721)
);

OAI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1596),
.A2(n_1634),
.B1(n_1553),
.B2(n_1531),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1607),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1594),
.A2(n_1519),
.B1(n_1524),
.B2(n_1573),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1631),
.A2(n_1616),
.B1(n_1673),
.B2(n_1678),
.Y(n_1725)
);

BUFx4f_ASAP7_75t_SL g1726 ( 
.A(n_1556),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1555),
.A2(n_1648),
.B1(n_1643),
.B2(n_1650),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1618),
.A2(n_1608),
.B1(n_1565),
.B2(n_1582),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1578),
.Y(n_1729)
);

OAI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1565),
.A2(n_1608),
.B1(n_1556),
.B2(n_1582),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_SL g1731 ( 
.A1(n_1685),
.A2(n_1606),
.B1(n_1645),
.B2(n_1614),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1582),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_SL g1733 ( 
.A1(n_1606),
.A2(n_1627),
.B1(n_1656),
.B2(n_1534),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1528),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1592),
.B(n_1609),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1623),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1527),
.B(n_1623),
.Y(n_1737)
);

OAI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1651),
.A2(n_1625),
.B(n_1637),
.C(n_1649),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1564),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1612),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1587),
.A2(n_1590),
.B1(n_1591),
.B2(n_1535),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1552),
.A2(n_1653),
.B1(n_1649),
.B2(n_1633),
.C(n_1632),
.Y(n_1742)
);

OAI211xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1651),
.A2(n_1637),
.B(n_1592),
.C(n_1625),
.Y(n_1743)
);

AOI22x1_ASAP7_75t_SL g1744 ( 
.A1(n_1595),
.A2(n_1679),
.B1(n_1602),
.B2(n_1546),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1533),
.A2(n_1554),
.B1(n_1644),
.B2(n_1522),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1533),
.A2(n_1554),
.B1(n_1644),
.B2(n_1522),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1595),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1545),
.A2(n_1563),
.B1(n_1570),
.B2(n_1629),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1679),
.B(n_1540),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1629),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1545),
.A2(n_1563),
.B1(n_1570),
.B2(n_1619),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1619),
.A2(n_1621),
.B1(n_1626),
.B2(n_1646),
.Y(n_1752)
);

OAI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1621),
.A2(n_1626),
.B1(n_1633),
.B2(n_1552),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1653),
.B(n_1652),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1569),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1593),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1569),
.A2(n_1572),
.B1(n_1646),
.B2(n_1647),
.Y(n_1757)
);

OAI21xp33_ASAP7_75t_L g1758 ( 
.A1(n_1635),
.A2(n_1632),
.B(n_1654),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1652),
.B(n_1599),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1636),
.A2(n_1665),
.B1(n_1666),
.B2(n_1663),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1647),
.B(n_1658),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1660),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1670),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1664),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1617),
.A2(n_1622),
.B1(n_1672),
.B2(n_1669),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1638),
.B(n_1657),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1657),
.A2(n_1667),
.B1(n_1642),
.B2(n_1662),
.C(n_1661),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1640),
.B(n_1641),
.C(n_1662),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1659),
.A2(n_1638),
.B1(n_1670),
.B2(n_1661),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1655),
.A2(n_1019),
.B1(n_1674),
.B2(n_1003),
.Y(n_1770)
);

OAI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1655),
.A2(n_1674),
.B(n_832),
.C(n_837),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_SL g1772 ( 
.A1(n_1655),
.A2(n_1680),
.B(n_1303),
.C(n_1019),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1668),
.B(n_1655),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1668),
.A2(n_1019),
.B1(n_1674),
.B2(n_1312),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1668),
.A2(n_1019),
.B1(n_1674),
.B2(n_1003),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1674),
.A2(n_1116),
.B1(n_829),
.B2(n_837),
.C(n_832),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1003),
.B2(n_832),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1526),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1684),
.B(n_1579),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1681),
.A2(n_1116),
.B1(n_1019),
.B2(n_1143),
.Y(n_1783)
);

AO31x2_ASAP7_75t_L g1784 ( 
.A1(n_1632),
.A2(n_1633),
.A3(n_1635),
.B(n_1653),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1681),
.A2(n_1019),
.B1(n_1003),
.B2(n_1116),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_SL g1786 ( 
.A1(n_1681),
.A2(n_1019),
.B1(n_1003),
.B2(n_1116),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1674),
.A2(n_829),
.B1(n_837),
.B2(n_832),
.C(n_1312),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1578),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1684),
.B(n_1579),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1003),
.B2(n_832),
.Y(n_1792)
);

INVx11_ASAP7_75t_L g1793 ( 
.A(n_1544),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1681),
.A2(n_837),
.B1(n_832),
.B2(n_899),
.C(n_880),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1519),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_L g1796 ( 
.A1(n_1674),
.A2(n_832),
.B(n_837),
.C(n_829),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1681),
.A2(n_837),
.B(n_832),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1557),
.B(n_1558),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1519),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1681),
.A2(n_837),
.B1(n_832),
.B2(n_899),
.C(n_880),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1003),
.B2(n_832),
.Y(n_1802)
);

CKINVDCx20_ASAP7_75t_R g1803 ( 
.A(n_1690),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1003),
.B2(n_832),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1519),
.Y(n_1805)
);

AOI21xp33_ASAP7_75t_L g1806 ( 
.A1(n_1681),
.A2(n_1680),
.B(n_837),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_829),
.B2(n_837),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1578),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1674),
.A2(n_1116),
.B1(n_829),
.B2(n_837),
.C(n_832),
.Y(n_1809)
);

OA21x2_ASAP7_75t_L g1810 ( 
.A1(n_1584),
.A2(n_1649),
.B(n_1621),
.Y(n_1810)
);

AOI222xp33_ASAP7_75t_L g1811 ( 
.A1(n_1674),
.A2(n_1312),
.B1(n_980),
.B2(n_1402),
.C1(n_899),
.C2(n_880),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_SL g1812 ( 
.A1(n_1681),
.A2(n_1019),
.B1(n_1003),
.B2(n_1116),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1684),
.B(n_1579),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1684),
.B(n_1579),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1681),
.A2(n_837),
.B1(n_832),
.B2(n_899),
.C(n_880),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1556),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1547),
.Y(n_1818)
);

OR2x6_ASAP7_75t_L g1819 ( 
.A(n_1596),
.B(n_1634),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1674),
.B(n_837),
.C(n_832),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_SL g1821 ( 
.A(n_1519),
.Y(n_1821)
);

AOI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1681),
.A2(n_837),
.B1(n_832),
.B2(n_899),
.C(n_880),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1823)
);

AOI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1681),
.A2(n_837),
.B1(n_832),
.B2(n_899),
.C(n_880),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1681),
.A2(n_1116),
.B1(n_1019),
.B2(n_1143),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1674),
.A2(n_1019),
.B1(n_1312),
.B2(n_1681),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1538),
.A2(n_1347),
.B(n_1384),
.Y(n_1827)
);

BUFx12f_ASAP7_75t_L g1828 ( 
.A(n_1690),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1764),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1763),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1782),
.B(n_1791),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1784),
.B(n_1810),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1784),
.B(n_1810),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1756),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1723),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1740),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1820),
.A2(n_1801),
.B1(n_1824),
.B2(n_1822),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1784),
.B(n_1810),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1784),
.B(n_1762),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1733),
.B(n_1751),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1766),
.B(n_1773),
.Y(n_1841)
);

NOR2x1_ASAP7_75t_L g1842 ( 
.A(n_1768),
.B(n_1722),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1692),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1692),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1751),
.B(n_1742),
.Y(n_1845)
);

OA21x2_ASAP7_75t_L g1846 ( 
.A1(n_1696),
.A2(n_1827),
.B(n_1758),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1754),
.B(n_1727),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1727),
.B(n_1769),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1769),
.B(n_1761),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1735),
.B(n_1759),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1719),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1692),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1729),
.Y(n_1853)
);

AND2x4_ASAP7_75t_SL g1854 ( 
.A(n_1757),
.B(n_1819),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1700),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1814),
.B(n_1815),
.Y(n_1856)
);

INVx4_ASAP7_75t_L g1857 ( 
.A(n_1747),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1748),
.B(n_1711),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1748),
.B(n_1790),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1790),
.B(n_1808),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1797),
.A2(n_1816),
.B(n_1794),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1713),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1716),
.B(n_1717),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1767),
.B(n_1753),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1780),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1752),
.B(n_1718),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1752),
.B(n_1738),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1765),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1734),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1760),
.Y(n_1870)
);

INVxp67_ASAP7_75t_SL g1871 ( 
.A(n_1753),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1745),
.B(n_1746),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1741),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1746),
.B(n_1710),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1743),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1772),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1701),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1818),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1699),
.B(n_1704),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1712),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1704),
.B(n_1731),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1715),
.B(n_1703),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1694),
.B(n_1703),
.Y(n_1883)
);

OA21x2_ASAP7_75t_L g1884 ( 
.A1(n_1771),
.A2(n_1806),
.B(n_1698),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1702),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1694),
.B(n_1695),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_1799),
.Y(n_1887)
);

BUFx10_ASAP7_75t_L g1888 ( 
.A(n_1854),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1861),
.A2(n_1796),
.B(n_1809),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1837),
.A2(n_1812),
.B(n_1785),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1847),
.B(n_1721),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1844),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1831),
.B(n_1698),
.Y(n_1893)
);

OAI322xp33_ASAP7_75t_L g1894 ( 
.A1(n_1861),
.A2(n_1777),
.A3(n_1783),
.B1(n_1825),
.B2(n_1770),
.C1(n_1695),
.C2(n_1807),
.Y(n_1894)
);

AO21x1_ASAP7_75t_SL g1895 ( 
.A1(n_1864),
.A2(n_1714),
.B(n_1721),
.Y(n_1895)
);

AO221x2_ASAP7_75t_L g1896 ( 
.A1(n_1883),
.A2(n_1697),
.B1(n_1825),
.B2(n_1783),
.C(n_1725),
.Y(n_1896)
);

AOI33xp33_ASAP7_75t_L g1897 ( 
.A1(n_1875),
.A2(n_1786),
.A3(n_1788),
.B1(n_1826),
.B2(n_1823),
.B3(n_1813),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1877),
.Y(n_1898)
);

OAI31xp33_ASAP7_75t_L g1899 ( 
.A1(n_1879),
.A2(n_1787),
.A3(n_1804),
.B(n_1802),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1847),
.B(n_1839),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1846),
.A2(n_1779),
.B(n_1792),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1830),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1829),
.Y(n_1903)
);

NOR2x1_ASAP7_75t_L g1904 ( 
.A(n_1842),
.B(n_1857),
.Y(n_1904)
);

OAI31xp33_ASAP7_75t_L g1905 ( 
.A1(n_1879),
.A2(n_1691),
.A3(n_1693),
.B(n_1775),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1880),
.A2(n_1813),
.B1(n_1826),
.B2(n_1781),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1866),
.A2(n_1811),
.B1(n_1823),
.B2(n_1776),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1851),
.A2(n_1714),
.B(n_1707),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1831),
.B(n_1725),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1846),
.A2(n_1886),
.B(n_1871),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1862),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1866),
.A2(n_1778),
.B1(n_1776),
.B2(n_1798),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1866),
.A2(n_1744),
.B1(n_1828),
.B2(n_1750),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1880),
.A2(n_1798),
.B1(n_1789),
.B2(n_1788),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1850),
.B(n_1841),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1834),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1834),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1835),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1835),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1842),
.B(n_1722),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1886),
.A2(n_1789),
.B(n_1781),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1883),
.A2(n_1778),
.B1(n_1774),
.B2(n_1724),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1836),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1867),
.A2(n_1774),
.B1(n_1724),
.B2(n_1720),
.Y(n_1924)
);

NAND5xp2_ASAP7_75t_L g1925 ( 
.A(n_1881),
.B(n_1720),
.C(n_1737),
.D(n_1749),
.E(n_1793),
.Y(n_1925)
);

AOI31xp33_ASAP7_75t_L g1926 ( 
.A1(n_1882),
.A2(n_1755),
.A3(n_1805),
.B(n_1795),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1850),
.B(n_1705),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1865),
.Y(n_1928)
);

AOI21x1_ASAP7_75t_L g1929 ( 
.A1(n_1876),
.A2(n_1709),
.B(n_1732),
.Y(n_1929)
);

OR2x6_ASAP7_75t_L g1930 ( 
.A(n_1843),
.B(n_1708),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1878),
.B(n_1800),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_SL g1932 ( 
.A1(n_1881),
.A2(n_1726),
.B1(n_1803),
.B2(n_1821),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1875),
.A2(n_1726),
.B1(n_1730),
.B2(n_1728),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1867),
.A2(n_1821),
.B1(n_1728),
.B2(n_1739),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1852),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1863),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1847),
.B(n_1839),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1839),
.B(n_1706),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1843),
.B(n_1817),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1863),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1863),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1850),
.B(n_1817),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1859),
.B(n_1706),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1885),
.B(n_1730),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1865),
.Y(n_1945)
);

INVxp67_ASAP7_75t_SL g1946 ( 
.A(n_1869),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1841),
.B(n_1736),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1830),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1841),
.B(n_1736),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1859),
.B(n_1708),
.Y(n_1950)
);

AOI322xp5_ASAP7_75t_L g1951 ( 
.A1(n_1867),
.A2(n_1881),
.A3(n_1871),
.B1(n_1845),
.B2(n_1874),
.C1(n_1840),
.C2(n_1870),
.Y(n_1951)
);

OAI211xp5_ASAP7_75t_L g1952 ( 
.A1(n_1864),
.A2(n_1882),
.B(n_1846),
.C(n_1874),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1900),
.B(n_1838),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1900),
.B(n_1838),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1915),
.B(n_1832),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1937),
.B(n_1838),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1915),
.B(n_1832),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1937),
.B(n_1832),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1940),
.B(n_1833),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1940),
.B(n_1833),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1930),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1940),
.B(n_1843),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1938),
.B(n_1833),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1938),
.B(n_1859),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1910),
.B(n_1858),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1930),
.B(n_1843),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1898),
.B(n_1858),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1911),
.B(n_1858),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1936),
.B(n_1846),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1941),
.B(n_1846),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1943),
.B(n_1872),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1943),
.B(n_1872),
.Y(n_1973)
);

NAND2x1p5_ASAP7_75t_L g1974 ( 
.A(n_1904),
.B(n_1843),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1950),
.B(n_1872),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1950),
.B(n_1860),
.Y(n_1976)
);

NOR3xp33_ASAP7_75t_L g1977 ( 
.A(n_1889),
.B(n_1864),
.C(n_1882),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1928),
.B(n_1849),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1928),
.B(n_1849),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1945),
.B(n_1849),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1892),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1916),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1916),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1917),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1917),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1918),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1918),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1919),
.B(n_1855),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1919),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1935),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1923),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1935),
.B(n_1946),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1930),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1947),
.B(n_1853),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1947),
.B(n_1853),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1983),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1989),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1962),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1965),
.B(n_1942),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1983),
.Y(n_2000)
);

NAND2x1_ASAP7_75t_L g2001 ( 
.A(n_1961),
.B(n_1993),
.Y(n_2001)
);

NAND2x1p5_ASAP7_75t_L g2002 ( 
.A(n_1961),
.B(n_1843),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1965),
.B(n_1878),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1953),
.B(n_1891),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1985),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1985),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1975),
.B(n_1942),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1955),
.B(n_1957),
.Y(n_2008)
);

AO21x1_ASAP7_75t_L g2009 ( 
.A1(n_1977),
.A2(n_1920),
.B(n_1905),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1975),
.B(n_1972),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1986),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1986),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1975),
.B(n_1927),
.Y(n_2013)
);

BUFx2_ASAP7_75t_SL g2014 ( 
.A(n_1981),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1953),
.B(n_1891),
.Y(n_2015)
);

OAI21xp33_ASAP7_75t_L g2016 ( 
.A1(n_1977),
.A2(n_1890),
.B(n_1951),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1982),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1953),
.B(n_1930),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1989),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1955),
.B(n_1957),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1991),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1982),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1954),
.B(n_1939),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1972),
.B(n_1927),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1987),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1954),
.B(n_1939),
.Y(n_2026)
);

AOI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_1966),
.A2(n_1896),
.B1(n_1901),
.B2(n_1874),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1991),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1954),
.B(n_1939),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1989),
.Y(n_2030)
);

NAND2x1_ASAP7_75t_L g2031 ( 
.A(n_1961),
.B(n_1948),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1972),
.B(n_1909),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1987),
.Y(n_2033)
);

AOI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1966),
.A2(n_1896),
.B1(n_1906),
.B2(n_1907),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1984),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_L g2036 ( 
.A(n_1993),
.B(n_1952),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1984),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1973),
.B(n_1949),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1956),
.B(n_1888),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1974),
.B(n_1932),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1984),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1984),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1956),
.B(n_1888),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1988),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1988),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1973),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1955),
.B(n_1949),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1993),
.B(n_1902),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_2010),
.B(n_1967),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_2009),
.B(n_1966),
.Y(n_2050)
);

INVxp67_ASAP7_75t_SL g2051 ( 
.A(n_2036),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2004),
.B(n_1956),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2004),
.B(n_1973),
.Y(n_2053)
);

OAI33xp33_ASAP7_75t_L g2054 ( 
.A1(n_2016),
.A2(n_1967),
.A3(n_1968),
.B1(n_1922),
.B2(n_1957),
.B3(n_1995),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2041),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1996),
.Y(n_2056)
);

INVxp67_ASAP7_75t_L g2057 ( 
.A(n_2003),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2000),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2005),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2046),
.B(n_1968),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_2041),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2015),
.B(n_1964),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_2034),
.B(n_1978),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2015),
.B(n_1964),
.Y(n_2064)
);

AND2x4_ASAP7_75t_SL g2065 ( 
.A(n_2048),
.B(n_1888),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2018),
.B(n_1964),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2032),
.B(n_1978),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2027),
.B(n_1978),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2006),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2018),
.B(n_1963),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2009),
.B(n_1931),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2019),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2011),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2019),
.Y(n_2074)
);

INVx3_ASAP7_75t_SL g2075 ( 
.A(n_2040),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2012),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2014),
.B(n_1963),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2013),
.B(n_1958),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_2040),
.B(n_1926),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2014),
.B(n_1963),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2044),
.B(n_1979),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2030),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2024),
.B(n_1958),
.Y(n_2083)
);

OAI31xp33_ASAP7_75t_L g2084 ( 
.A1(n_2002),
.A2(n_1899),
.A3(n_1925),
.B(n_1924),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_1999),
.B(n_1958),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2023),
.B(n_1976),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2045),
.B(n_1979),
.Y(n_2087)
);

NOR2x1_ASAP7_75t_R g2088 ( 
.A(n_2048),
.B(n_1944),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_2025),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2030),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2021),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2028),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2007),
.B(n_1979),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2023),
.B(n_2026),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2017),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2017),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2047),
.B(n_1971),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2026),
.B(n_1976),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2022),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2022),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_R g2101 ( 
.A(n_2048),
.B(n_1929),
.Y(n_2101)
);

NOR2xp67_ASAP7_75t_R g2102 ( 
.A(n_1998),
.B(n_1948),
.Y(n_2102)
);

AOI211xp5_ASAP7_75t_SL g2103 ( 
.A1(n_2071),
.A2(n_1894),
.B(n_1933),
.C(n_1845),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2056),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2056),
.Y(n_2105)
);

OAI322xp33_ASAP7_75t_L g2106 ( 
.A1(n_2050),
.A2(n_2001),
.A3(n_2020),
.B1(n_2008),
.B2(n_2031),
.C1(n_2002),
.C2(n_2047),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2058),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2057),
.B(n_2029),
.Y(n_2108)
);

OAI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2075),
.A2(n_1913),
.B1(n_2001),
.B2(n_2031),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2058),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2089),
.Y(n_2111)
);

OAI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_2075),
.A2(n_1912),
.B1(n_1974),
.B2(n_1914),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_2075),
.Y(n_2113)
);

OAI32xp33_ASAP7_75t_SL g2114 ( 
.A1(n_2054),
.A2(n_1896),
.A3(n_2033),
.B1(n_2008),
.B2(n_2020),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_2088),
.Y(n_2115)
);

NAND3xp33_ASAP7_75t_L g2116 ( 
.A(n_2051),
.B(n_1896),
.C(n_1921),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2079),
.A2(n_1966),
.B1(n_1840),
.B2(n_1845),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2059),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2094),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_2065),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2063),
.A2(n_1966),
.B1(n_1840),
.B2(n_1885),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_2084),
.A2(n_2002),
.B(n_1974),
.C(n_1893),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2094),
.B(n_1998),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2059),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2084),
.B(n_2029),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2068),
.B(n_2038),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2053),
.Y(n_2127)
);

AOI21xp33_ASAP7_75t_SL g2128 ( 
.A1(n_2088),
.A2(n_1974),
.B(n_1884),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2065),
.B(n_2039),
.Y(n_2129)
);

AOI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_2065),
.A2(n_1870),
.B1(n_1884),
.B2(n_1848),
.Y(n_2130)
);

AOI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2077),
.A2(n_1884),
.B1(n_1848),
.B2(n_2043),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2053),
.B(n_1980),
.Y(n_2132)
);

AOI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2077),
.A2(n_1884),
.B1(n_1848),
.B2(n_2043),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2069),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2080),
.A2(n_1884),
.B1(n_2039),
.B2(n_1970),
.Y(n_2135)
);

OAI31xp33_ASAP7_75t_L g2136 ( 
.A1(n_2080),
.A2(n_1934),
.A3(n_1981),
.B(n_1868),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_2066),
.A2(n_1969),
.B1(n_1970),
.B2(n_1962),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2066),
.B(n_1998),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_2095),
.B(n_1897),
.C(n_1873),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_2095),
.A2(n_1908),
.B(n_1969),
.Y(n_2140)
);

OAI32xp33_ASAP7_75t_L g2141 ( 
.A1(n_2060),
.A2(n_1990),
.A3(n_1970),
.B1(n_1969),
.B2(n_1994),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_2062),
.B(n_1962),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2113),
.B(n_2103),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2111),
.B(n_2049),
.Y(n_2144)
);

OAI221xp5_ASAP7_75t_L g2145 ( 
.A1(n_2122),
.A2(n_2096),
.B1(n_2100),
.B2(n_2099),
.C(n_2049),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2104),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_2116),
.B(n_2101),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2123),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2115),
.A2(n_2064),
.B1(n_2062),
.B2(n_2052),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2105),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2113),
.B(n_2052),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2109),
.A2(n_2064),
.B1(n_2087),
.B2(n_2081),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2107),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2123),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2103),
.B(n_2086),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2110),
.Y(n_2156)
);

AOI322xp5_ASAP7_75t_L g2157 ( 
.A1(n_2125),
.A2(n_2070),
.A3(n_2067),
.B1(n_2093),
.B2(n_2098),
.C1(n_2086),
.C2(n_2099),
.Y(n_2157)
);

INVxp67_ASAP7_75t_SL g2158 ( 
.A(n_2129),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2120),
.B(n_2070),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_2108),
.B(n_2085),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2118),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2112),
.A2(n_2096),
.B1(n_2100),
.B2(n_2069),
.Y(n_2162)
);

O2A1O1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_2128),
.A2(n_2076),
.B(n_2073),
.C(n_2092),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2124),
.Y(n_2164)
);

INVxp67_ASAP7_75t_SL g2165 ( 
.A(n_2130),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2134),
.Y(n_2166)
);

AOI221xp5_ASAP7_75t_L g2167 ( 
.A1(n_2114),
.A2(n_2073),
.B1(n_2092),
.B2(n_2076),
.C(n_2091),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2119),
.Y(n_2168)
);

NAND4xp75_ASAP7_75t_SL g2169 ( 
.A(n_2136),
.B(n_1929),
.C(n_2102),
.D(n_2098),
.Y(n_2169)
);

AO22x1_ASAP7_75t_L g2170 ( 
.A1(n_2140),
.A2(n_2091),
.B1(n_1990),
.B2(n_1962),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2126),
.B(n_2085),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2151),
.B(n_2159),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2144),
.Y(n_2173)
);

INVxp67_ASAP7_75t_SL g2174 ( 
.A(n_2158),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2143),
.B(n_2117),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2151),
.Y(n_2176)
);

NOR2xp67_ASAP7_75t_L g2177 ( 
.A(n_2144),
.B(n_2121),
.Y(n_2177)
);

NOR3xp33_ASAP7_75t_SL g2178 ( 
.A(n_2147),
.B(n_2106),
.C(n_2139),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2155),
.B(n_2136),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2146),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_2171),
.B(n_2168),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2159),
.B(n_2127),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2150),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2153),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2165),
.B(n_2131),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_2160),
.B(n_2133),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2149),
.B(n_2132),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2148),
.B(n_2138),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2156),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2160),
.B(n_2135),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_2148),
.Y(n_2191)
);

CKINVDCx16_ASAP7_75t_R g2192 ( 
.A(n_2162),
.Y(n_2192)
);

NOR3xp33_ASAP7_75t_SL g2193 ( 
.A(n_2147),
.B(n_2141),
.C(n_2140),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2161),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2154),
.B(n_2142),
.Y(n_2195)
);

NOR4xp25_ASAP7_75t_L g2196 ( 
.A(n_2175),
.B(n_2174),
.C(n_2173),
.D(n_2179),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_2192),
.B(n_2145),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2191),
.Y(n_2198)
);

INVx1_ASAP7_75t_SL g2199 ( 
.A(n_2172),
.Y(n_2199)
);

AOI211xp5_ASAP7_75t_L g2200 ( 
.A1(n_2185),
.A2(n_2163),
.B(n_2170),
.C(n_2167),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2191),
.Y(n_2201)
);

NOR2x1_ASAP7_75t_L g2202 ( 
.A(n_2184),
.B(n_2169),
.Y(n_2202)
);

NOR4xp25_ASAP7_75t_L g2203 ( 
.A(n_2184),
.B(n_2166),
.C(n_2164),
.D(n_2154),
.Y(n_2203)
);

NOR3xp33_ASAP7_75t_L g2204 ( 
.A(n_2186),
.B(n_2152),
.C(n_2142),
.Y(n_2204)
);

NAND2x1_ASAP7_75t_L g2205 ( 
.A(n_2172),
.B(n_2137),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2176),
.B(n_2157),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_SL g2207 ( 
.A(n_2177),
.B(n_1857),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2188),
.B(n_2178),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2181),
.Y(n_2209)
);

AOI211x1_ASAP7_75t_SL g2210 ( 
.A1(n_2206),
.A2(n_2195),
.B(n_2190),
.C(n_2182),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_2201),
.Y(n_2211)
);

OAI211xp5_ASAP7_75t_SL g2212 ( 
.A1(n_2200),
.A2(n_2193),
.B(n_2181),
.C(n_2183),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_2198),
.B(n_2188),
.Y(n_2213)
);

AOI221xp5_ASAP7_75t_L g2214 ( 
.A1(n_2196),
.A2(n_2189),
.B1(n_2180),
.B2(n_2194),
.C(n_2187),
.Y(n_2214)
);

O2A1O1Ixp5_ASAP7_75t_SL g2215 ( 
.A1(n_2209),
.A2(n_2194),
.B(n_2187),
.C(n_2035),
.Y(n_2215)
);

OAI211xp5_ASAP7_75t_SL g2216 ( 
.A1(n_2197),
.A2(n_2208),
.B(n_2202),
.C(n_2199),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2207),
.B(n_2078),
.Y(n_2217)
);

OAI21xp5_ASAP7_75t_SL g2218 ( 
.A1(n_2204),
.A2(n_2207),
.B(n_2205),
.Y(n_2218)
);

O2A1O1Ixp33_ASAP7_75t_L g2219 ( 
.A1(n_2203),
.A2(n_2060),
.B(n_2078),
.C(n_2083),
.Y(n_2219)
);

OAI221xp5_ASAP7_75t_L g2220 ( 
.A1(n_2196),
.A2(n_2083),
.B1(n_2055),
.B2(n_2061),
.C(n_2082),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2211),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2213),
.B(n_2097),
.Y(n_2222)
);

INVx1_ASAP7_75t_SL g2223 ( 
.A(n_2213),
.Y(n_2223)
);

AND4x1_ASAP7_75t_L g2224 ( 
.A(n_2210),
.B(n_1992),
.C(n_1959),
.D(n_1960),
.Y(n_2224)
);

NAND3xp33_ASAP7_75t_L g2225 ( 
.A(n_2214),
.B(n_2055),
.C(n_2061),
.Y(n_2225)
);

NAND2x1p5_ASAP7_75t_L g2226 ( 
.A(n_2217),
.B(n_1857),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2218),
.B(n_2097),
.Y(n_2227)
);

OAI21xp33_ASAP7_75t_SL g2228 ( 
.A1(n_2215),
.A2(n_2090),
.B(n_2082),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2223),
.B(n_2216),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2221),
.B(n_2219),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2222),
.Y(n_2231)
);

NOR3xp33_ASAP7_75t_L g2232 ( 
.A(n_2227),
.B(n_2212),
.C(n_2220),
.Y(n_2232)
);

INVx2_ASAP7_75t_SL g2233 ( 
.A(n_2226),
.Y(n_2233)
);

INVx1_ASAP7_75t_SL g2234 ( 
.A(n_2225),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2228),
.A2(n_2061),
.B1(n_2055),
.B2(n_2074),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2224),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2229),
.Y(n_2237)
);

AO22x2_ASAP7_75t_L g2238 ( 
.A1(n_2236),
.A2(n_2090),
.B1(n_2082),
.B2(n_2074),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_2229),
.B(n_2072),
.Y(n_2239)
);

NOR3xp33_ASAP7_75t_L g2240 ( 
.A(n_2232),
.B(n_2090),
.C(n_2074),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2230),
.Y(n_2241)
);

NOR3xp33_ASAP7_75t_L g2242 ( 
.A(n_2231),
.B(n_2072),
.C(n_1856),
.Y(n_2242)
);

NAND3xp33_ASAP7_75t_L g2243 ( 
.A(n_2237),
.B(n_2233),
.C(n_2235),
.Y(n_2243)
);

NAND3xp33_ASAP7_75t_L g2244 ( 
.A(n_2239),
.B(n_2234),
.C(n_2072),
.Y(n_2244)
);

AO22x1_ASAP7_75t_L g2245 ( 
.A1(n_2241),
.A2(n_2240),
.B1(n_2242),
.B2(n_2238),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2237),
.Y(n_2246)
);

INVx1_ASAP7_75t_SL g2247 ( 
.A(n_2246),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2243),
.B(n_1997),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2248),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2249),
.B(n_2248),
.Y(n_2250)
);

CKINVDCx20_ASAP7_75t_R g2251 ( 
.A(n_2249),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2250),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2251),
.A2(n_2247),
.B1(n_2244),
.B2(n_2245),
.Y(n_2253)
);

OAI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2253),
.A2(n_1997),
.B(n_2037),
.Y(n_2254)
);

AOI222xp33_ASAP7_75t_L g2255 ( 
.A1(n_2254),
.A2(n_2252),
.B1(n_2042),
.B2(n_1992),
.C1(n_1962),
.C2(n_1887),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_R g2256 ( 
.A1(n_2255),
.A2(n_1895),
.B1(n_1948),
.B2(n_1989),
.C(n_1857),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2256),
.A2(n_1992),
.B1(n_1948),
.B2(n_1960),
.Y(n_2257)
);


endmodule