module fake_jpeg_19316_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_46),
.B(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_47),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_12),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_60),
.B(n_74),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_63),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_72),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_66),
.Y(n_123)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_76),
.Y(n_107)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_78),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_2),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_80),
.B(n_82),
.Y(n_139)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_83),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_3),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

OR2x4_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_16),
.B1(n_28),
.B2(n_36),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_98),
.B1(n_104),
.B2(n_113),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_16),
.B1(n_39),
.B2(n_36),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_57),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_16),
.B1(n_39),
.B2(n_34),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_102),
.A2(n_114),
.B1(n_116),
.B2(n_133),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_16),
.B1(n_24),
.B2(n_33),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_26),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_125),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_26),
.B1(n_22),
.B2(n_33),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_22),
.B1(n_27),
.B2(n_25),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_52),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_81),
.B1(n_79),
.B2(n_49),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_130),
.B1(n_123),
.B2(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_50),
.B(n_20),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_47),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_54),
.A2(n_35),
.B1(n_32),
.B2(n_23),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_56),
.B(n_40),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_136),
.B(n_137),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_44),
.B(n_40),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_85),
.A2(n_35),
.B1(n_32),
.B2(n_23),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_71),
.B1(n_66),
.B2(n_35),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_53),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_140),
.A2(n_146),
.B(n_153),
.Y(n_206)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_40),
.B1(n_29),
.B2(n_32),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_144),
.A2(n_165),
.B(n_97),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_145),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_44),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_100),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_152),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_106),
.B(n_45),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_45),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_106),
.B(n_68),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_68),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_164),
.Y(n_188)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_130),
.A2(n_111),
.B1(n_139),
.B2(n_94),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_110),
.A2(n_75),
.B1(n_51),
.B2(n_53),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_107),
.A2(n_29),
.B1(n_57),
.B2(n_7),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_111),
.A2(n_29),
.B1(n_5),
.B2(n_7),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_169),
.A2(n_171),
.B1(n_180),
.B2(n_182),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_184),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_4),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_173),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_112),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_179),
.B1(n_183),
.B2(n_185),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_92),
.B(n_8),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_175),
.B(n_91),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_8),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_174),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_10),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_186),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_11),
.B1(n_117),
.B2(n_123),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_94),
.A2(n_11),
.B1(n_103),
.B2(n_105),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_131),
.C(n_91),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_103),
.A2(n_11),
.B1(n_105),
.B2(n_120),
.Y(n_182)
);

AO22x2_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_109),
.B1(n_115),
.B2(n_134),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_93),
.B(n_124),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_117),
.A2(n_132),
.B1(n_124),
.B2(n_108),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_189),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_193),
.B(n_225),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_121),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_196),
.A2(n_199),
.B(n_208),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_131),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_197),
.B(n_212),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_115),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_201),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_109),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_141),
.B(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_108),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_119),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_149),
.B(n_119),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_140),
.B(n_150),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_140),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_232),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_181),
.B1(n_148),
.B2(n_159),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_228),
.A2(n_229),
.B1(n_237),
.B2(n_239),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_199),
.A2(n_144),
.B1(n_167),
.B2(n_173),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_230),
.B(n_234),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_171),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_235),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_171),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_162),
.B1(n_172),
.B2(n_183),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_187),
.A2(n_183),
.B1(n_158),
.B2(n_142),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_187),
.A2(n_183),
.B1(n_143),
.B2(n_174),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_244),
.B1(n_256),
.B2(n_196),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_175),
.C(n_176),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_246),
.C(n_248),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_183),
.B1(n_174),
.B2(n_155),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_186),
.C(n_151),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_164),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_189),
.B(n_145),
.C(n_174),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_221),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_202),
.B(n_214),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_225),
.B1(n_197),
.B2(n_200),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_190),
.B1(n_213),
.B2(n_218),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_191),
.B(n_216),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_261),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_208),
.A2(n_220),
.B1(n_190),
.B2(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_205),
.B(n_190),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_265),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_196),
.B1(n_205),
.B2(n_215),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_267),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_213),
.B(n_195),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_268),
.A2(n_258),
.B(n_239),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_195),
.C(n_193),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_275),
.C(n_277),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_198),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_251),
.C(n_236),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_192),
.C(n_223),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_233),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_198),
.B(n_194),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_281),
.B(n_287),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_194),
.B(n_192),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_242),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_240),
.B(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_232),
.B(n_223),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_289),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_202),
.B(n_214),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_237),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_211),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_252),
.B(n_202),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_291),
.B(n_243),
.CI(n_229),
.CON(n_304),
.SN(n_304)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_259),
.B(n_235),
.C(n_231),
.D(n_257),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_275),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_246),
.C(n_258),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_317),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_295),
.B(n_299),
.Y(n_320)
);

BUFx12_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_296),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_263),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_310),
.Y(n_322)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

BUFx12f_ASAP7_75t_SL g306 ( 
.A(n_288),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_306),
.A2(n_316),
.B1(n_311),
.B2(n_283),
.Y(n_331)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_314),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_298),
.B(n_308),
.Y(n_323)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_245),
.C(n_255),
.Y(n_317)
);

OA22x2_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_285),
.B1(n_288),
.B2(n_262),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_329),
.B1(n_331),
.B2(n_338),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_321),
.B(n_272),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_323),
.A2(n_330),
.B(n_312),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_285),
.B1(n_262),
.B2(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_281),
.B(n_280),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_304),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_303),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_333),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_267),
.B1(n_285),
.B2(n_289),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_298),
.A2(n_277),
.B(n_271),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_303),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_272),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_272),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_297),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_316),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_300),
.A2(n_264),
.B1(n_274),
.B2(n_266),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_300),
.A2(n_278),
.B1(n_270),
.B2(n_234),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_339),
.A2(n_301),
.B1(n_302),
.B2(n_273),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_293),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_343),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_356),
.C(n_357),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_317),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_349),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_345),
.A2(n_354),
.B(n_334),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_347),
.B(n_353),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_294),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_319),
.Y(n_358)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

AOI21xp33_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_278),
.B(n_301),
.Y(n_353)
);

A2O1A1O1Ixp25_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_304),
.B(n_292),
.C(n_312),
.D(n_276),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_326),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_302),
.C(n_310),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_309),
.C(n_307),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_363),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_340),
.A2(n_339),
.B1(n_322),
.B2(n_328),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_361),
.A2(n_355),
.B1(n_337),
.B2(n_324),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_296),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_364),
.B(n_340),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_366),
.B(n_273),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_346),
.A2(n_348),
.B(n_334),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_357),
.A2(n_329),
.B1(n_338),
.B2(n_319),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_370),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_356),
.B(n_327),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_378),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_336),
.B(n_318),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_374),
.A2(n_382),
.B(n_305),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_343),
.C(n_359),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_379),
.C(n_381),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_376),
.A2(n_371),
.B1(n_291),
.B2(n_366),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_318),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_341),
.C(n_342),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_349),
.C(n_344),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_369),
.A2(n_337),
.B(n_324),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_375),
.B(n_368),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_386),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_361),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_367),
.C(n_360),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_381),
.C(n_313),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_390),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_360),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_378),
.B(n_376),
.Y(n_392)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_297),
.Y(n_395)
);

AOI321xp33_ASAP7_75t_SL g399 ( 
.A1(n_395),
.A2(n_290),
.A3(n_238),
.B1(n_214),
.B2(n_226),
.C(n_384),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_397),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_383),
.A2(n_390),
.B(n_387),
.Y(n_397)
);

AOI322xp5_ASAP7_75t_L g398 ( 
.A1(n_393),
.A2(n_296),
.A3(n_260),
.B1(n_255),
.B2(n_384),
.C1(n_238),
.C2(n_226),
.Y(n_398)
);

BUFx24_ASAP7_75t_SL g403 ( 
.A(n_398),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_399),
.B(n_401),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_402),
.Y(n_404)
);

NOR3xp33_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_394),
.C(n_400),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_226),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_404),
.Y(n_407)
);


endmodule