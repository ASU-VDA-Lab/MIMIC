module fake_jpeg_27636_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_38),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_43),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_19),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_17),
.B(n_30),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_57),
.C(n_22),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_25),
.B1(n_16),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_38),
.B1(n_24),
.B2(n_26),
.Y(n_69)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_17),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_30),
.C(n_25),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_57),
.C(n_43),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_60),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_35),
.B(n_33),
.C(n_28),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_66),
.B(n_58),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_77),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_41),
.B(n_2),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_41),
.A3(n_27),
.B1(n_22),
.B2(n_38),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_58),
.B(n_46),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_19),
.B1(n_46),
.B2(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_70),
.B(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_47),
.B1(n_49),
.B2(n_43),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_27),
.B1(n_29),
.B2(n_24),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_22),
.B1(n_17),
.B2(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_80),
.B(n_29),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_74),
.B1(n_69),
.B2(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_95),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_92),
.B(n_94),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_3),
.B(n_4),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_3),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_14),
.B(n_12),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_9),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_9),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_59),
.B(n_72),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_4),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_67),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_110),
.Y(n_131)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_118),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_89),
.B1(n_81),
.B2(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_114),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_92),
.B(n_91),
.C(n_88),
.D(n_99),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_103),
.B(n_118),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_96),
.C(n_71),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.C(n_120),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_96),
.B1(n_64),
.B2(n_6),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_115),
.B1(n_106),
.B2(n_105),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_139),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_146),
.C(n_128),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_115),
.B(n_112),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_144),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_107),
.C(n_64),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_152),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_146),
.C(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_134),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_140),
.B(n_143),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_130),
.C(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_125),
.B1(n_148),
.B2(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_166),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_161),
.B(n_7),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_148),
.B1(n_147),
.B2(n_8),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_159),
.C(n_162),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_173),
.B1(n_167),
.B2(n_164),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_8),
.Y(n_176)
);


endmodule