module fake_netlist_1_7145_n_722 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_722);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_722;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g80 ( .A(n_44), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_15), .Y(n_81) );
BUFx3_ASAP7_75t_L g82 ( .A(n_45), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_24), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_64), .Y(n_84) );
INVxp33_ASAP7_75t_L g85 ( .A(n_23), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_63), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_49), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_4), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_74), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_70), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_67), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_54), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_19), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_60), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_79), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_7), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_27), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_26), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_62), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_17), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_78), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_33), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_65), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_9), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_12), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_32), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_34), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_75), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_1), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_36), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_43), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_73), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_42), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_35), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_61), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_31), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_55), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_16), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_68), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_109), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_126), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_84), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_84), .B(n_0), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_118), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_100), .Y(n_139) );
XNOR2xp5_ASAP7_75t_L g140 ( .A(n_101), .B(n_0), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_126), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_108), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_82), .B(n_25), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_120), .B(n_1), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_82), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_90), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_105), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_82), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_80), .B(n_2), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_86), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_96), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_117), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_127), .B(n_3), .Y(n_155) );
CKINVDCx8_ASAP7_75t_R g156 ( .A(n_124), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_104), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_127), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_88), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_96), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_89), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_92), .Y(n_163) );
NOR2xp33_ASAP7_75t_R g164 ( .A(n_89), .B(n_29), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_91), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_87), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_94), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_123), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_91), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_95), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_85), .B(n_3), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_121), .B(n_4), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_95), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_163), .B(n_129), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_135), .B(n_111), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_135), .B(n_111), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
OR2x2_ASAP7_75t_L g179 ( .A(n_145), .B(n_110), .Y(n_179) );
NAND3x1_ASAP7_75t_L g180 ( .A(n_150), .B(n_110), .C(n_128), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_134), .B(n_129), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_133), .B(n_97), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g185 ( .A(n_156), .B(n_139), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_138), .A2(n_128), .B1(n_81), .B2(n_93), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_132), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_152), .B(n_97), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_169), .B(n_112), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_137), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_160), .B(n_127), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_147), .A2(n_112), .B1(n_98), .B2(n_106), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_162), .B(n_125), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_170), .B(n_93), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_171), .B(n_98), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_159), .B(n_99), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
INVx8_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_141), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_136), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_173), .B(n_106), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_143), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_141), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_158), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_159), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_146), .A2(n_114), .B1(n_115), .B2(n_102), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_171), .B(n_114), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_159), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_172), .Y(n_223) );
NAND2xp33_ASAP7_75t_SL g224 ( .A(n_172), .B(n_115), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_142), .B(n_125), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_159), .B(n_122), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_143), .B(n_122), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_166), .B(n_119), .Y(n_228) );
OR2x2_ASAP7_75t_SL g229 ( .A(n_140), .B(n_119), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_157), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_143), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_167), .B(n_116), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_149), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_168), .B(n_116), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_143), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_143), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_130), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_155), .B(n_113), .Y(n_238) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_140), .A2(n_113), .B1(n_107), .B2(n_103), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_144), .Y(n_240) );
AO22x1_ASAP7_75t_L g241 ( .A1(n_227), .A2(n_99), .B1(n_103), .B2(n_107), .Y(n_241) );
NOR3xp33_ASAP7_75t_SL g242 ( .A(n_237), .B(n_154), .C(n_148), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_230), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_176), .B(n_161), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_218), .Y(n_245) );
BUFx12f_ASAP7_75t_L g246 ( .A(n_230), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_176), .B(n_153), .Y(n_247) );
NOR3xp33_ASAP7_75t_SL g248 ( .A(n_237), .B(n_156), .C(n_164), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_209), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_194), .B(n_5), .Y(n_251) );
AND2x6_ASAP7_75t_L g252 ( .A(n_236), .B(n_30), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_177), .B(n_5), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_219), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_204), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_218), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_211), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_223), .B(n_6), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_212), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_202), .B(n_6), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_177), .B(n_7), .Y(n_262) );
NAND2xp33_ASAP7_75t_SL g263 ( .A(n_214), .B(n_8), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_202), .B(n_8), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_180), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_192), .Y(n_267) );
NOR3xp33_ASAP7_75t_SL g268 ( .A(n_199), .B(n_10), .C(n_11), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_224), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_221), .B(n_13), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_189), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_192), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_189), .Y(n_273) );
NAND3xp33_ASAP7_75t_SL g274 ( .A(n_220), .B(n_15), .C(n_18), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_204), .Y(n_275) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_214), .B(n_18), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_221), .B(n_19), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_209), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_214), .B(n_20), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_216), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_219), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_193), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_222), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_217), .Y(n_284) );
NOR3xp33_ASAP7_75t_SL g285 ( .A(n_224), .B(n_20), .C(n_21), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_225), .B(n_22), .C(n_28), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_222), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_193), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_240), .B(n_37), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_198), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_235), .Y(n_291) );
NOR3xp33_ASAP7_75t_SL g292 ( .A(n_174), .B(n_38), .C(n_39), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_182), .B(n_40), .Y(n_293) );
NAND2xp33_ASAP7_75t_SL g294 ( .A(n_235), .B(n_41), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_234), .B(n_46), .Y(n_295) );
NOR2xp33_ASAP7_75t_R g296 ( .A(n_185), .B(n_47), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_198), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g298 ( .A1(n_186), .A2(n_48), .B1(n_50), .B2(n_51), .C(n_52), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_207), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_207), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_175), .B(n_53), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_235), .A2(n_56), .B(n_58), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_210), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_191), .B(n_77), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_210), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_215), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_191), .B(n_66), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_178), .B(n_76), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_215), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_231), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_204), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_244), .B(n_233), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_255), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_261), .B(n_234), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_251), .B(n_201), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_310), .A2(n_231), .B(n_204), .Y(n_316) );
INVx5_ASAP7_75t_L g317 ( .A(n_252), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_258), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_261), .B(n_234), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_261), .B(n_191), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_264), .A2(n_239), .B1(n_213), .B2(n_201), .C(n_233), .Y(n_321) );
O2A1O1Ixp5_ASAP7_75t_L g322 ( .A1(n_241), .A2(n_197), .B(n_226), .C(n_200), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_310), .A2(n_231), .B(n_204), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_272), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_255), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_259), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_243), .B(n_229), .Y(n_327) );
AOI21xp5_ASAP7_75t_SL g328 ( .A1(n_304), .A2(n_236), .B(n_213), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_258), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_246), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_265), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_264), .B(n_213), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_264), .B(n_201), .Y(n_334) );
NOR2x1_ASAP7_75t_SL g335 ( .A(n_244), .B(n_236), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_299), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_255), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_276), .A2(n_180), .B1(n_179), .B2(n_236), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_270), .B(n_232), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_246), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_244), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_276), .B(n_203), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_259), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_253), .A2(n_179), .B(n_197), .C(n_232), .Y(n_344) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_263), .B(n_228), .C(n_208), .Y(n_345) );
INVx4_ASAP7_75t_L g346 ( .A(n_244), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_277), .B(n_181), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_247), .A2(n_183), .B1(n_190), .B2(n_187), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_245), .Y(n_349) );
BUFx12f_ASAP7_75t_L g350 ( .A(n_267), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_297), .A2(n_227), .B(n_188), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_267), .B(n_239), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_301), .A2(n_184), .B(n_195), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_307), .B(n_238), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_308), .A2(n_196), .B(n_206), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_245), .Y(n_356) );
NAND2xp33_ASAP7_75t_L g357 ( .A(n_255), .B(n_227), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_304), .B(n_205), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_247), .B(n_239), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_304), .B(n_205), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_247), .B(n_239), .Y(n_361) );
INVxp67_ASAP7_75t_L g362 ( .A(n_247), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_242), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_259), .B(n_238), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_262), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_307), .B(n_205), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_342), .B(n_279), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_353), .A2(n_302), .B(n_279), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
NAND2xp33_ASAP7_75t_SL g371 ( .A(n_338), .B(n_296), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_320), .B(n_268), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_362), .B(n_229), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_359), .A2(n_274), .B1(n_263), .B2(n_266), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_SL g376 ( .A1(n_348), .A2(n_289), .B(n_293), .C(n_298), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_320), .B(n_260), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_324), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_359), .A2(n_295), .B1(n_245), .B2(n_256), .Y(n_380) );
AND2x6_ASAP7_75t_L g381 ( .A(n_334), .B(n_265), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_257), .B(n_280), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_359), .A2(n_256), .B1(n_249), .B2(n_269), .Y(n_384) );
INVx6_ASAP7_75t_L g385 ( .A(n_341), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_361), .A2(n_279), .B1(n_227), .B2(n_205), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_342), .A2(n_284), .B1(n_297), .B2(n_305), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_318), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_334), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_313), .Y(n_390) );
INVx4_ASAP7_75t_SL g391 ( .A(n_361), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_313), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_361), .B(n_305), .Y(n_393) );
NAND2x1_ASAP7_75t_L g394 ( .A(n_313), .B(n_282), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_312), .Y(n_395) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_315), .A2(n_283), .B(n_256), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_347), .Y(n_397) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_313), .B(n_282), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_312), .Y(n_399) );
NAND2xp33_ASAP7_75t_R g400 ( .A(n_330), .B(n_248), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_375), .A2(n_321), .B1(n_352), .B2(n_312), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_315), .B1(n_350), .B2(n_341), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_379), .A2(n_346), .B1(n_333), .B2(n_314), .Y(n_403) );
NAND3xp33_ASAP7_75t_SL g404 ( .A(n_379), .B(n_363), .C(n_285), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_397), .A2(n_339), .B1(n_344), .B2(n_319), .C(n_362), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_373), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_397), .A2(n_350), .B1(n_346), .B2(n_365), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_373), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_383), .B(n_286), .C(n_292), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_393), .B(n_327), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_367), .B(n_364), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_372), .A2(n_363), .B1(n_343), .B2(n_326), .C(n_354), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_395), .A2(n_335), .B1(n_340), .B2(n_345), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_382), .A2(n_354), .B1(n_366), .B2(n_205), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_378), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
AO21x2_ASAP7_75t_L g418 ( .A1(n_376), .A2(n_369), .B(n_396), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_367), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_378), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_370), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_393), .B(n_328), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_399), .B(n_283), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_387), .A2(n_322), .B(n_358), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_370), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_391), .A2(n_368), .B1(n_389), .B2(n_380), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_391), .A2(n_205), .B1(n_294), .B2(n_227), .Y(n_428) );
AND2x6_ASAP7_75t_L g429 ( .A(n_391), .B(n_360), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_406), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_406), .Y(n_431) );
OAI33xp33_ASAP7_75t_L g432 ( .A1(n_403), .A2(n_377), .A3(n_391), .B1(n_400), .B2(n_371), .B3(n_384), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_406), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_419), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_410), .A2(n_368), .B1(n_385), .B2(n_389), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_412), .B(n_368), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_401), .A2(n_368), .B1(n_381), .B2(n_385), .Y(n_437) );
AOI221xp5_ASAP7_75t_SL g438 ( .A1(n_405), .A2(n_355), .B1(n_388), .B2(n_351), .C(n_357), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_404), .A2(n_368), .B1(n_381), .B2(n_385), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_419), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_421), .B(n_388), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_408), .A2(n_386), .B1(n_385), .B2(n_317), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_412), .B(n_388), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_421), .Y(n_445) );
AOI31xp33_ASAP7_75t_L g446 ( .A1(n_427), .A2(n_294), .A3(n_390), .B(n_392), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_411), .B(n_388), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_410), .A2(n_322), .B(n_369), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_413), .A2(n_241), .B1(n_249), .B2(n_349), .C(n_356), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_422), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_402), .A2(n_381), .B1(n_356), .B2(n_349), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_415), .A2(n_381), .B1(n_252), .B2(n_227), .C1(n_357), .C2(n_317), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
OAI31xp33_ASAP7_75t_SL g455 ( .A1(n_414), .A2(n_390), .A3(n_392), .B(n_381), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_422), .B(n_300), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_409), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_409), .B(n_300), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_416), .B(n_306), .Y(n_461) );
AOI21xp5_ASAP7_75t_SL g462 ( .A1(n_416), .A2(n_337), .B(n_325), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_411), .Y(n_463) );
AOI31xp33_ASAP7_75t_L g464 ( .A1(n_423), .A2(n_381), .A3(n_317), .B(n_250), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_424), .B(n_249), .C(n_398), .Y(n_465) );
OAI21x1_ASAP7_75t_L g466 ( .A1(n_416), .A2(n_398), .B(n_394), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_435), .A2(n_423), .B1(n_428), .B2(n_425), .C(n_417), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_463), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_458), .A2(n_425), .B1(n_426), .B2(n_417), .C(n_418), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_430), .B(n_417), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_455), .B(n_426), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_432), .A2(n_426), .B1(n_418), .B2(n_273), .C(n_282), .Y(n_474) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_449), .A2(n_418), .B(n_323), .Y(n_475) );
OR2x6_ASAP7_75t_L g476 ( .A(n_430), .B(n_420), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_450), .A2(n_381), .B1(n_429), .B2(n_252), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_435), .A2(n_394), .B1(n_273), .B2(n_288), .C(n_303), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_434), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_433), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_433), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_454), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_447), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_440), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_432), .B(n_303), .C(n_290), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_454), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_460), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_459), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_459), .B(n_420), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_445), .B(n_420), .Y(n_494) );
INVx4_ASAP7_75t_L g495 ( .A(n_444), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_451), .B(n_429), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_447), .Y(n_497) );
INVx5_ASAP7_75t_SL g498 ( .A(n_447), .Y(n_498) );
OAI21xp33_ASAP7_75t_SL g499 ( .A1(n_455), .A2(n_317), .B(n_429), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_444), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_444), .Y(n_501) );
OAI31xp33_ASAP7_75t_L g502 ( .A1(n_442), .A2(n_318), .A3(n_332), .B(n_329), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_420), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_451), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_443), .B(n_429), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_456), .B(n_420), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_457), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_456), .Y(n_508) );
AOI31xp33_ASAP7_75t_L g509 ( .A1(n_439), .A2(n_429), .A3(n_250), .B(n_278), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_456), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_456), .B(n_420), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_436), .B(n_306), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_438), .B(n_309), .C(n_254), .Y(n_513) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_441), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_436), .B(n_309), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_457), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_443), .B(n_429), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_466), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_516), .B(n_448), .Y(n_519) );
NOR2xp33_ASAP7_75t_R g520 ( .A(n_473), .B(n_437), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_468), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_504), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_491), .B(n_449), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_491), .B(n_460), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_471), .B(n_461), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_484), .Y(n_526) );
XNOR2x1_ASAP7_75t_L g527 ( .A(n_512), .B(n_448), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_504), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_492), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_492), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_507), .B(n_441), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_490), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_471), .B(n_461), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_472), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_481), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_481), .B(n_442), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_495), .B(n_466), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_482), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_485), .B(n_446), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_470), .B(n_465), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_512), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_487), .B(n_446), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_470), .B(n_483), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_487), .B(n_438), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_482), .B(n_464), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_472), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_486), .B(n_462), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_489), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_489), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_478), .A2(n_450), .B1(n_452), .B2(n_429), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_486), .B(n_462), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_494), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_477), .Y(n_558) );
AOI21xp33_ASAP7_75t_L g559 ( .A1(n_499), .A2(n_464), .B(n_453), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_489), .B(n_332), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_477), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_489), .B(n_290), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_501), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_515), .Y(n_564) );
NAND2xp33_ASAP7_75t_SL g565 ( .A(n_495), .B(n_453), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_479), .B(n_288), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_479), .B(n_429), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_497), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_497), .B(n_288), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_495), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_510), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_517), .B(n_273), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_510), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_517), .B(n_290), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_509), .B(n_329), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_505), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_500), .B(n_252), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_526), .A2(n_499), .B(n_467), .C(n_502), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_571), .B(n_538), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_540), .A2(n_473), .B(n_478), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_522), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_528), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_551), .B(n_469), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_529), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_543), .B(n_495), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_537), .A2(n_473), .B1(n_488), .B2(n_501), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_537), .A2(n_498), .B1(n_493), .B2(n_511), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_540), .A2(n_518), .B(n_493), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_530), .Y(n_590) );
CKINVDCx14_ASAP7_75t_R g591 ( .A(n_521), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_564), .B(n_532), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_565), .A2(n_498), .B1(n_493), .B2(n_511), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_552), .B(n_498), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_550), .B(n_502), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_545), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_565), .A2(n_480), .B1(n_474), .B2(n_518), .C(n_476), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_550), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_542), .Y(n_600) );
AO22x1_ASAP7_75t_L g601 ( .A1(n_521), .A2(n_493), .B1(n_518), .B2(n_500), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_553), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_520), .A2(n_498), .B1(n_506), .B2(n_503), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_524), .B(n_476), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_557), .B(n_508), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_546), .B(n_508), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_524), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_525), .B(n_506), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_559), .A2(n_513), .B(n_476), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_534), .Y(n_610) );
AOI21xp33_ASAP7_75t_SL g611 ( .A1(n_547), .A2(n_476), .B(n_513), .Y(n_611) );
NAND2x1_ASAP7_75t_L g612 ( .A(n_571), .B(n_503), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_575), .A2(n_475), .B(n_303), .C(n_271), .Y(n_613) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_562), .A2(n_475), .B(n_254), .Y(n_614) );
CKINVDCx14_ASAP7_75t_R g615 ( .A(n_520), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_572), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_527), .A2(n_271), .B1(n_287), .B2(n_281), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_525), .B(n_475), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_539), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_527), .B(n_252), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_574), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_576), .B(n_271), .C(n_287), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_519), .Y(n_623) );
INVxp67_ASAP7_75t_R g624 ( .A(n_549), .Y(n_624) );
OAI22xp5_ASAP7_75t_SL g625 ( .A1(n_554), .A2(n_278), .B1(n_252), .B2(n_337), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_541), .A2(n_281), .B(n_316), .C(n_291), .Y(n_626) );
AOI211xp5_ASAP7_75t_L g627 ( .A1(n_544), .A2(n_325), .B(n_337), .C(n_291), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_570), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g629 ( .A1(n_577), .A2(n_325), .B1(n_337), .B2(n_311), .C1(n_255), .C2(n_275), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_582), .Y(n_630) );
NOR2x1_ASAP7_75t_L g631 ( .A(n_599), .B(n_538), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_581), .A2(n_523), .B(n_563), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g633 ( .A(n_586), .B(n_573), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_592), .B(n_555), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_611), .B(n_538), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_596), .B(n_531), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_585), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_590), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_597), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_600), .Y(n_641) );
NAND2xp33_ASAP7_75t_L g642 ( .A(n_622), .B(n_560), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_599), .B(n_580), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_623), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_628), .B(n_533), .Y(n_645) );
NAND2x1_ASAP7_75t_L g646 ( .A(n_580), .B(n_558), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_602), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_617), .A2(n_549), .B(n_567), .C(n_568), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_615), .A2(n_561), .B1(n_556), .B2(n_548), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_616), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_607), .B(n_556), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_591), .A2(n_560), .B1(n_548), .B2(n_536), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_621), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_608), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_606), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_612), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_619), .B(n_536), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_602), .B(n_566), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_606), .B(n_569), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_617), .A2(n_578), .B(n_325), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_618), .B(n_578), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_605), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_610), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_603), .B(n_275), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_604), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_655), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_632), .B(n_595), .C(n_579), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_662), .B(n_584), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_630), .Y(n_669) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_642), .B(n_613), .Y(n_670) );
NOR2xp67_ASAP7_75t_L g671 ( .A(n_656), .B(n_593), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_652), .A2(n_624), .B1(n_588), .B2(n_587), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_664), .A2(n_609), .B(n_627), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_637), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_646), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_638), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_639), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_640), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_664), .A2(n_601), .B(n_589), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_631), .B(n_643), .Y(n_680) );
NAND2xp33_ASAP7_75t_SL g681 ( .A(n_643), .B(n_594), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_644), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_654), .A2(n_620), .B1(n_584), .B2(n_625), .Y(n_683) );
BUFx3_ASAP7_75t_L g684 ( .A(n_658), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g685 ( .A1(n_635), .A2(n_598), .B(n_614), .C(n_626), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_634), .B(n_614), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_657), .B(n_629), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g688 ( .A(n_633), .B(n_629), .Y(n_688) );
AOI311xp33_ASAP7_75t_L g689 ( .A1(n_667), .A2(n_648), .A3(n_657), .B(n_650), .C(n_641), .Y(n_689) );
NOR2xp33_ASAP7_75t_R g690 ( .A(n_681), .B(n_647), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_682), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_667), .A2(n_649), .B1(n_635), .B2(n_636), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_668), .B(n_647), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_687), .B(n_653), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_666), .Y(n_695) );
XOR2xp5_ASAP7_75t_L g696 ( .A(n_688), .B(n_652), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_686), .B(n_659), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_682), .Y(n_698) );
BUFx2_ASAP7_75t_L g699 ( .A(n_680), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_669), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g701 ( .A1(n_672), .A2(n_645), .B1(n_663), .B2(n_665), .C1(n_660), .C2(n_661), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_674), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_681), .A2(n_275), .B1(n_311), .B2(n_651), .C(n_685), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_670), .A2(n_275), .B1(n_311), .B2(n_671), .Y(n_704) );
OAI211xp5_ASAP7_75t_SL g705 ( .A1(n_685), .A2(n_275), .B(n_311), .C(n_673), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_683), .A2(n_311), .B1(n_680), .B2(n_684), .Y(n_706) );
AOI211xp5_ASAP7_75t_L g707 ( .A1(n_679), .A2(n_675), .B(n_676), .C(n_677), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_678), .A2(n_667), .B1(n_672), .B2(n_688), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_696), .A2(n_708), .B(n_707), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_695), .Y(n_710) );
NAND2x1_ASAP7_75t_L g711 ( .A(n_699), .B(n_675), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_698), .A2(n_691), .B(n_705), .C(n_699), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_690), .Y(n_713) );
OAI211xp5_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_689), .B(n_690), .C(n_701), .Y(n_714) );
OAI322xp33_ASAP7_75t_L g715 ( .A1(n_709), .A2(n_692), .A3(n_706), .B1(n_694), .B2(n_704), .C1(n_693), .C2(n_700), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_711), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_716), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_714), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g719 ( .A(n_717), .B(n_715), .Y(n_719) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_718), .Y(n_720) );
OAI221xp5_ASAP7_75t_R g721 ( .A1(n_719), .A2(n_712), .B1(n_703), .B2(n_710), .C(n_697), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_720), .B(n_702), .Y(n_722) );
endmodule