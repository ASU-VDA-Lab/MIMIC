module fake_jpeg_1789_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx8_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_33),
.Y(n_43)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_28),
.B1(n_32),
.B2(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_52),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_49),
.B1(n_37),
.B2(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_23),
.B1(n_13),
.B2(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_14),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_65),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_69),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_50),
.B(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_70),
.Y(n_77)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_22),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_53),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_19),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_37),
.B1(n_35),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_77),
.B1(n_71),
.B2(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_77),
.B1(n_86),
.B2(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_62),
.B(n_55),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_74),
.B(n_67),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_99),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_60),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_54),
.C(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_103),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

OA21x2_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_110),
.B(n_48),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_36),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_94),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_96),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_118),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_110),
.B(n_93),
.CI(n_96),
.CON(n_113),
.SN(n_113)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_102),
.A3(n_37),
.B1(n_12),
.B2(n_5),
.C1(n_9),
.C2(n_4),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_77),
.B1(n_99),
.B2(n_69),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_117),
.B1(n_119),
.B2(n_36),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_61),
.C(n_41),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_111),
.C(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_56),
.B1(n_53),
.B2(n_51),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_104),
.Y(n_122)
);

OAI321xp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_100),
.A3(n_102),
.B1(n_108),
.B2(n_26),
.C(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_114),
.B(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_128),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_117),
.B1(n_116),
.B2(n_113),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_3),
.A3(n_4),
.B1(n_30),
.B2(n_128),
.C1(n_130),
.C2(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.Y(n_137)
);


endmodule