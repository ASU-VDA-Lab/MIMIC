module fake_jpeg_5851_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_39),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_43),
.Y(n_67)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_22),
.B1(n_27),
.B2(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_68),
.B1(n_16),
.B2(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_22),
.B1(n_27),
.B2(n_32),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_19),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_83),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_43),
.B1(n_18),
.B2(n_21),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_53),
.B1(n_57),
.B2(n_31),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_39),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_40),
.B(n_33),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_33),
.B(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_20),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_39),
.C(n_37),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_20),
.B1(n_18),
.B2(n_51),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_39),
.B1(n_16),
.B2(n_17),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_94),
.B1(n_64),
.B2(n_47),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_21),
.B1(n_17),
.B2(n_23),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_114),
.B(n_29),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_66),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_108),
.Y(n_132)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_101),
.Y(n_133)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_112),
.Y(n_123)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_113),
.Y(n_141)
);

AO22x2_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_84),
.B1(n_87),
.B2(n_83),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_83),
.B1(n_77),
.B2(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_69),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_120),
.B1(n_122),
.B2(n_88),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_54),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_63),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_99),
.B1(n_119),
.B2(n_95),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_77),
.B(n_72),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_142),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_37),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_144),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_30),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_140),
.Y(n_165)
);

NAND2x1_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_37),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_120),
.B(n_34),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_82),
.B1(n_74),
.B2(n_81),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_137),
.B1(n_148),
.B2(n_116),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_139),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_71),
.B1(n_58),
.B2(n_79),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_37),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_19),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_73),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_52),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_95),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_101),
.A2(n_57),
.B1(n_30),
.B2(n_19),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_163),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_100),
.C(n_106),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_162),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_140),
.B1(n_134),
.B2(n_30),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_38),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_129),
.C(n_139),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_157),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_76),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_124),
.B1(n_148),
.B2(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_159),
.B(n_169),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_171),
.B(n_31),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_52),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_172),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_49),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_38),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_113),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_49),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_30),
.B1(n_19),
.B2(n_31),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_140),
.B1(n_124),
.B2(n_137),
.Y(n_181)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_70),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_0),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_165),
.B1(n_176),
.B2(n_164),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_185),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_126),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_29),
.B(n_34),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_70),
.B1(n_31),
.B2(n_29),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_171),
.B1(n_155),
.B2(n_25),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_195),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_38),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_152),
.C(n_149),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_201),
.B(n_1),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_206),
.C(n_224),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_215),
.B1(n_201),
.B2(n_183),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_161),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_210),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_161),
.B(n_164),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_221),
.B(n_183),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_165),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_165),
.B1(n_29),
.B2(n_25),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_10),
.C(n_15),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_227),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_189),
.B1(n_182),
.B2(n_178),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_34),
.Y(n_224)
);

AO22x1_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_179),
.B(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_206),
.C(n_205),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_244),
.C(n_10),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_237),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_238),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_182),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_210),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_180),
.B1(n_196),
.B2(n_181),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_246),
.B1(n_204),
.B2(n_3),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_186),
.C(n_202),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_198),
.B1(n_192),
.B2(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_3),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_254),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_216),
.B1(n_221),
.B2(n_213),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_245),
.B1(n_239),
.B2(n_243),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_225),
.CI(n_224),
.CON(n_255),
.SN(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_266),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_240),
.B(n_250),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_249),
.B(n_240),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_268),
.C(n_229),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_9),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_245),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_7),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_270),
.C(n_276),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_229),
.C(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_264),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_252),
.B1(n_257),
.B2(n_251),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_277),
.B(n_265),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_234),
.C(n_244),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_236),
.B(n_239),
.Y(n_277)
);

BUFx12_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_267),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_246),
.B(n_235),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_255),
.C(n_8),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_258),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_284),
.A2(n_285),
.B(n_277),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_292),
.Y(n_305)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_293),
.C(n_294),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_283),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_269),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_235),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_255),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_280),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_279),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_7),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_271),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_296),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_8),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_13),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_302),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_270),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_272),
.B1(n_275),
.B2(n_282),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_287),
.B1(n_276),
.B2(n_278),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_13),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_306),
.A2(n_278),
.B(n_12),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_312),
.B(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_14),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_318),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_315),
.A3(n_311),
.B1(n_320),
.B2(n_317),
.C1(n_305),
.C2(n_299),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_305),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_14),
.B(n_15),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_14),
.Y(n_327)
);


endmodule