module fake_jpeg_608_n_231 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_231);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_66),
.Y(n_89)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_77),
.B1(n_72),
.B2(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_66),
.B1(n_76),
.B2(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_60),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_73),
.B1(n_68),
.B2(n_75),
.Y(n_98)
);

OA22x2_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_76),
.B1(n_60),
.B2(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_56),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_107),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_114),
.B1(n_116),
.B2(n_98),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_100),
.B1(n_59),
.B2(n_2),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_75),
.B1(n_68),
.B2(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_119),
.B1(n_79),
.B2(n_91),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_81),
.B1(n_67),
.B2(n_70),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_76),
.B1(n_73),
.B2(n_63),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_121),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_79),
.B1(n_61),
.B2(n_63),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_55),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_69),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_0),
.Y(n_142)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_140),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_100),
.B1(n_59),
.B2(n_2),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_154)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_7),
.B(n_8),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_124),
.B1(n_122),
.B2(n_118),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_40),
.B(n_36),
.Y(n_171)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_51),
.Y(n_148)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_7),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_1),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_4),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_54),
.C(n_52),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_126),
.C(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_50),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_17),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_147),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_161),
.B1(n_165),
.B2(n_16),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_3),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_159),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_49),
.C(n_48),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_165),
.C(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_6),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_141),
.B(n_47),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_169),
.B(n_139),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_171),
.B1(n_156),
.B2(n_160),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_8),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_144),
.B(n_132),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_144),
.B1(n_139),
.B2(n_11),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_32),
.A3(n_28),
.B1(n_27),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_178),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_179),
.B1(n_183),
.B2(n_185),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_169),
.B(n_170),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_172),
.B(n_158),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_182),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_192)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_171),
.B(n_163),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_194),
.A2(n_202),
.B(n_189),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_181),
.C(n_173),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_197),
.B1(n_193),
.B2(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_198),
.B(n_177),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_184),
.C(n_188),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_200),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_175),
.B1(n_182),
.B2(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_191),
.Y(n_212)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_200),
.B1(n_195),
.B2(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_209),
.C(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_201),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_215),
.B1(n_214),
.B2(n_216),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_220),
.C(n_218),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_223),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_218),
.B(n_217),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_204),
.A3(n_196),
.B1(n_22),
.B2(n_24),
.C(n_21),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_183),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_196),
.Y(n_231)
);


endmodule