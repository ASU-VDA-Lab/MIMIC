module fake_jpeg_30542_n_451 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_57),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_55),
.B(n_87),
.Y(n_120)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_25),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_19),
.B(n_16),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_68),
.Y(n_112)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_80),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_14),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_88),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_13),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_37),
.Y(n_131)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_42),
.B(n_27),
.C(n_30),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_95),
.B(n_129),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_42),
.B1(n_27),
.B2(n_21),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_97),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_99),
.B(n_109),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_51),
.A2(n_42),
.B(n_33),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_105),
.B(n_121),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_117),
.B(n_118),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_38),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_33),
.B(n_30),
.Y(n_121)
);

NAND2x1_ASAP7_75t_L g129 ( 
.A(n_47),
.B(n_74),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_45),
.A2(n_23),
.B1(n_28),
.B2(n_21),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_167)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_68),
.C(n_81),
.Y(n_143)
);

FAx1_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_97),
.CI(n_93),
.CON(n_184),
.SN(n_184)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_87),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_154),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_147),
.A2(n_137),
.B(n_102),
.Y(n_208)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_64),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx12_ASAP7_75t_R g152 ( 
.A(n_96),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_23),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_48),
.B1(n_67),
.B2(n_69),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_156),
.A2(n_161),
.B1(n_166),
.B2(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_159),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_82),
.B1(n_78),
.B2(n_77),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_28),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_169),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_76),
.B1(n_28),
.B2(n_23),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_177),
.B1(n_73),
.B2(n_62),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_37),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_114),
.B(n_36),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_33),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_178),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_95),
.A2(n_58),
.B1(n_46),
.B2(n_53),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_92),
.B(n_34),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_127),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_172),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_141),
.B1(n_108),
.B2(n_107),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_201),
.B1(n_167),
.B2(n_174),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_34),
.B(n_32),
.C(n_124),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_168),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_107),
.B1(n_111),
.B2(n_128),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_159),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_127),
.B1(n_128),
.B2(n_115),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_172),
.A2(n_115),
.B1(n_103),
.B2(n_136),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_98),
.B1(n_137),
.B2(n_102),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_157),
.C(n_151),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_224),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_212),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_151),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_151),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_202),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_206),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_203),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_230),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_186),
.B1(n_208),
.B2(n_188),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_222),
.B(n_227),
.Y(n_239)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_150),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_143),
.C(n_175),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_165),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_226),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_175),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_136),
.B1(n_135),
.B2(n_173),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_198),
.B1(n_164),
.B2(n_145),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_142),
.B1(n_148),
.B2(n_144),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_178),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_188),
.Y(n_257)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_226),
.A2(n_184),
.B1(n_204),
.B2(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_261),
.Y(n_268)
);

AO22x2_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_184),
.B1(n_205),
.B2(n_199),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_236),
.A2(n_260),
.B1(n_222),
.B2(n_228),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_251),
.B1(n_254),
.B2(n_256),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_186),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_247),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_216),
.A2(n_202),
.B1(n_189),
.B2(n_198),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_229),
.B1(n_210),
.B2(n_218),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_176),
.B1(n_190),
.B2(n_145),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_211),
.B(n_190),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_225),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_264),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_253),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_276),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_266),
.B(n_273),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_217),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_269),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_213),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_214),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

AOI32xp33_ASAP7_75t_L g272 ( 
.A1(n_236),
.A2(n_219),
.A3(n_220),
.B1(n_227),
.B2(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_288),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_259),
.B(n_230),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_211),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_275),
.B(n_281),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_248),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_248),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_282),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_236),
.A2(n_193),
.B1(n_215),
.B2(n_98),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_260),
.B1(n_247),
.B2(n_237),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_256),
.B(n_224),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_258),
.B(n_209),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_250),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_236),
.A2(n_215),
.B(n_152),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_289),
.B(n_189),
.Y(n_308)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_233),
.Y(n_287)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_243),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_239),
.A2(n_193),
.B(n_215),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_291),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_195),
.Y(n_291)
);

XOR2x1_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_235),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_294),
.B(n_315),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_300),
.A2(n_316),
.B1(n_318),
.B2(n_320),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_235),
.B(n_255),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_302),
.A2(n_307),
.B(n_308),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_242),
.C(n_245),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_303),
.B(n_306),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_237),
.B1(n_254),
.B2(n_239),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_304),
.A2(n_262),
.B1(n_290),
.B2(n_283),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_242),
.C(n_261),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_289),
.B(n_160),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_267),
.B(n_195),
.Y(n_310)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_162),
.Y(n_314)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_279),
.B(n_124),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_270),
.A2(n_182),
.B1(n_191),
.B2(n_149),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_192),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_284),
.A2(n_268),
.B(n_283),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_281),
.A2(n_182),
.B1(n_153),
.B2(n_164),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_171),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_321),
.B(n_265),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_268),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_337),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_329),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_308),
.A2(n_270),
.B(n_274),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_297),
.A2(n_287),
.B1(n_271),
.B2(n_269),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_325),
.A2(n_328),
.B1(n_330),
.B2(n_334),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_286),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_263),
.B1(n_277),
.B2(n_282),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_263),
.B1(n_276),
.B2(n_288),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_342),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_275),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_298),
.A2(n_283),
.B(n_262),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_341),
.B(n_345),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_291),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_340),
.B(n_305),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_300),
.A2(n_283),
.B(n_285),
.Y(n_341)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_292),
.B1(n_182),
.B2(n_149),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_346),
.A2(n_320),
.B1(n_316),
.B2(n_299),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_301),
.C(n_309),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_350),
.C(n_357),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_301),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_353),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_302),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_361),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_309),
.C(n_312),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_295),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_331),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_360),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_312),
.C(n_313),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_344),
.B(n_296),
.Y(n_360)
);

XNOR2x1_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_295),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_310),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_362),
.B(n_333),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_365),
.C(n_366),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_293),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_343),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_343),
.A2(n_313),
.B1(n_293),
.B2(n_299),
.Y(n_368)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_341),
.B1(n_338),
.B2(n_327),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_367),
.A2(n_346),
.B1(n_332),
.B2(n_327),
.Y(n_372)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_356),
.A2(n_333),
.B1(n_307),
.B2(n_292),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_125),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_376),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_292),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_347),
.B(n_192),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_377),
.B(n_12),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_366),
.A2(n_153),
.B1(n_221),
.B2(n_234),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_380),
.A2(n_387),
.B1(n_350),
.B2(n_361),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_357),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_384),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_234),
.B(n_221),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_383),
.A2(n_385),
.B(n_355),
.Y(n_389)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_179),
.B(n_104),
.Y(n_385)
);

AO22x1_ASAP7_75t_L g387 ( 
.A1(n_365),
.A2(n_104),
.B1(n_135),
.B2(n_138),
.Y(n_387)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_403),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_364),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_392),
.A2(n_393),
.B1(n_395),
.B2(n_398),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_378),
.A2(n_349),
.B1(n_358),
.B2(n_61),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_397),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_358),
.C(n_70),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_401),
.C(n_380),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_400),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_381),
.C(n_386),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_379),
.B(n_386),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_402),
.B(n_382),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_SL g404 ( 
.A(n_401),
.B(n_387),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_407),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_SL g408 ( 
.A(n_396),
.B(n_374),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_408),
.A2(n_414),
.B(n_389),
.Y(n_420)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_409),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_382),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_413),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_403),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_400),
.A2(n_385),
.B1(n_371),
.B2(n_383),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_390),
.A2(n_134),
.B(n_1),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_70),
.C(n_125),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_0),
.C(n_1),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_419),
.B(n_420),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_405),
.A2(n_134),
.B1(n_125),
.B2(n_3),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_423),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_0),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_0),
.Y(n_425)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_425),
.A2(n_426),
.B(n_1),
.Y(n_431)
);

AOI21xp33_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_410),
.B(n_412),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_411),
.C(n_416),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_429),
.B(n_430),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_411),
.C(n_3),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_431),
.Y(n_439)
);

NAND2x1p5_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_4),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_434),
.Y(n_438)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_417),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_435),
.A2(n_422),
.B(n_423),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_5),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_5),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_437),
.B(n_442),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_440),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_6),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_441),
.B(n_433),
.C(n_436),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_445),
.B(n_439),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_446),
.A2(n_447),
.B(n_444),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_438),
.C(n_432),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_435),
.C(n_8),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_7),
.Y(n_451)
);


endmodule