module fake_jpeg_3431_n_469 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_49),
.B(n_50),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_55),
.Y(n_98)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_53),
.Y(n_147)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_59),
.Y(n_101)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g146 ( 
.A(n_58),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_62),
.Y(n_113)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_65),
.B(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_0),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_2),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_91),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_41),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_41),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_96),
.A2(n_24),
.B1(n_39),
.B2(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_24),
.B(n_2),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_97),
.B(n_40),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_39),
.B1(n_30),
.B2(n_32),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_105),
.A2(n_117),
.B1(n_131),
.B2(n_141),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_41),
.B(n_40),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_108),
.A2(n_58),
.B(n_83),
.C(n_80),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_54),
.A2(n_39),
.B1(n_30),
.B2(n_32),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_67),
.A2(n_21),
.B1(n_45),
.B2(n_43),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_122),
.A2(n_124),
.B1(n_130),
.B2(n_132),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_70),
.A2(n_21),
.B1(n_45),
.B2(n_43),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_49),
.A2(n_47),
.B1(n_25),
.B2(n_23),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_32),
.B1(n_26),
.B2(n_40),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_50),
.A2(n_47),
.B1(n_25),
.B2(n_23),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_82),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_53),
.A2(n_31),
.B1(n_41),
.B2(n_34),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_48),
.A2(n_31),
.B1(n_41),
.B2(n_34),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_75),
.B1(n_123),
.B2(n_61),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_65),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_77),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_68),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_69),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_150),
.B1(n_152),
.B2(n_12),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_84),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_87),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_108),
.A2(n_84),
.B(n_78),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_155),
.A2(n_194),
.B(n_192),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_90),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_161),
.B(n_162),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_102),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_163),
.A2(n_180),
.B(n_188),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_52),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_170),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_166),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_179),
.B1(n_139),
.B2(n_123),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_88),
.Y(n_170)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_85),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_71),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_72),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_189),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_57),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_192),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_114),
.B(n_75),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_205),
.C(n_128),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_94),
.B1(n_89),
.B2(n_73),
.Y(n_179)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_104),
.Y(n_183)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx6_ASAP7_75t_SL g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_185),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_101),
.B(n_81),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2x1_ASAP7_75t_SL g188 ( 
.A(n_114),
.B(n_135),
.Y(n_188)
);

INVx2_ASAP7_75t_R g189 ( 
.A(n_110),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_115),
.B(n_8),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_191),
.B(n_195),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_10),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_197),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_133),
.A2(n_11),
.B(n_12),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_113),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_196),
.A2(n_129),
.B1(n_107),
.B2(n_145),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_137),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_120),
.B(n_12),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_200),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_112),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_115),
.B(n_12),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_157),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_215),
.A2(n_220),
.B1(n_235),
.B2(n_247),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_177),
.A2(n_134),
.B1(n_153),
.B2(n_127),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_153),
.B1(n_134),
.B2(n_127),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_221),
.A2(n_227),
.B1(n_167),
.B2(n_203),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_106),
.B1(n_125),
.B2(n_138),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_231),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_125),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_175),
.C(n_163),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_234),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_163),
.A2(n_106),
.B1(n_148),
.B2(n_149),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_193),
.B(n_190),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_156),
.A2(n_128),
.B1(n_109),
.B2(n_112),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_178),
.B(n_151),
.C(n_109),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_248),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_155),
.B(n_151),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_156),
.A2(n_129),
.B1(n_107),
.B2(n_145),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_264),
.Y(n_306)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_211),
.B(n_205),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_257),
.B(n_268),
.Y(n_295)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_169),
.B(n_185),
.C(n_183),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_259),
.A2(n_263),
.B(n_232),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_201),
.B(n_175),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_269),
.B(n_279),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_258),
.B1(n_215),
.B2(n_220),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_158),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_273),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_214),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_168),
.B(n_199),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_225),
.A2(n_198),
.B1(n_199),
.B2(n_169),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_270),
.A2(n_184),
.B1(n_196),
.B2(n_167),
.Y(n_317)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_210),
.Y(n_272)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_245),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_232),
.B(n_228),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_269),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_230),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_278),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_204),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_174),
.B(n_181),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_173),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_208),
.B(n_224),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_224),
.B(n_208),
.Y(n_290)
);

NOR2x1_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_263),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_231),
.C(n_238),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_293),
.C(n_303),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_298),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_291),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_241),
.C(n_232),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_270),
.A2(n_266),
.B1(n_274),
.B2(n_261),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_300),
.B1(n_305),
.B2(n_308),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_235),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_243),
.C(n_223),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_315),
.C(n_283),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_221),
.B1(n_244),
.B2(n_219),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_244),
.B1(n_243),
.B2(n_236),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_209),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_275),
.A2(n_216),
.B(n_222),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_321),
.B(n_259),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_319),
.B1(n_320),
.B2(n_260),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_278),
.A2(n_268),
.B1(n_252),
.B2(n_267),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_267),
.A2(n_184),
.B1(n_160),
.B2(n_202),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_260),
.A2(n_216),
.B(n_222),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_322),
.A2(n_301),
.B(n_321),
.Y(n_363)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_324),
.Y(n_364)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_276),
.C(n_287),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_313),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_307),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_329),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_347),
.B(n_348),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_315),
.B(n_263),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_333),
.B(n_344),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_263),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_340),
.C(n_341),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_339),
.Y(n_357)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_337),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_257),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_264),
.C(n_272),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_281),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_282),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_309),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_295),
.B(n_189),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_297),
.B(n_265),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_345),
.B(n_351),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_346),
.A2(n_285),
.B1(n_284),
.B2(n_309),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_298),
.A2(n_259),
.B(n_260),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_296),
.A2(n_256),
.B(n_255),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_350),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_296),
.B(n_279),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_342),
.A2(n_299),
.B1(n_288),
.B2(n_320),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_352),
.A2(n_358),
.B1(n_349),
.B2(n_351),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_304),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_355),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_291),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_342),
.A2(n_300),
.B1(n_303),
.B2(n_298),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_301),
.C(n_314),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_369),
.C(n_375),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_363),
.A2(n_331),
.B(n_347),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_346),
.A2(n_305),
.B1(n_308),
.B2(n_310),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_373),
.B1(n_371),
.B2(n_341),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_292),
.C(n_302),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_338),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_335),
.B(n_253),
.Y(n_375)
);

AO22x1_ASAP7_75t_SL g376 ( 
.A1(n_351),
.A2(n_294),
.B1(n_253),
.B2(n_286),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_294),
.C(n_166),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_332),
.C(n_350),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_397),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_327),
.Y(n_383)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_392),
.Y(n_401)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_367),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_387),
.A2(n_388),
.B1(n_391),
.B2(n_394),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_360),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_368),
.C(n_357),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_396),
.B(n_358),
.Y(n_411)
);

FAx1_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_349),
.CI(n_322),
.CON(n_398),
.SN(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g416 ( 
.A1(n_398),
.A2(n_376),
.B(n_280),
.C(n_271),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_377),
.A2(n_348),
.B(n_329),
.Y(n_399)
);

AOI21x1_ASAP7_75t_L g408 ( 
.A1(n_399),
.A2(n_376),
.B(n_365),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_369),
.B(n_339),
.Y(n_400)
);

OAI322xp33_ASAP7_75t_L g406 ( 
.A1(n_400),
.A2(n_355),
.A3(n_344),
.B1(n_368),
.B2(n_357),
.C1(n_356),
.C2(n_375),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_402),
.B(n_400),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_353),
.C(n_378),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_406),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_374),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_416),
.Y(n_424)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_352),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_413),
.C(n_398),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_356),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_420),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_395),
.C(n_388),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_383),
.Y(n_421)
);

OAI21x1_ASAP7_75t_SL g444 ( 
.A1(n_421),
.A2(n_398),
.B(n_380),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_387),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_427),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_415),
.A2(n_392),
.B1(n_397),
.B2(n_381),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_401),
.B1(n_416),
.B2(n_408),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_405),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_407),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_429),
.B(n_430),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_379),
.C(n_385),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_399),
.C(n_380),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_413),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_401),
.Y(n_433)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_436),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_410),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_437),
.A2(n_418),
.B1(n_394),
.B2(n_389),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_440),
.B(n_423),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_417),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_441),
.B(n_414),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_424),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_443),
.A2(n_444),
.B1(n_405),
.B2(n_384),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_445),
.B(n_446),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_431),
.C(n_428),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_425),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_447),
.B(n_448),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_425),
.C(n_382),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_443),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_SL g454 ( 
.A(n_451),
.B(n_453),
.Y(n_454)
);

NAND3xp33_ASAP7_75t_SL g455 ( 
.A(n_450),
.B(n_438),
.C(n_439),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_455),
.A2(n_456),
.B(n_457),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_435),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_458),
.A2(n_451),
.B(n_446),
.Y(n_461)
);

AOI21x1_ASAP7_75t_L g465 ( 
.A1(n_461),
.A2(n_454),
.B(n_218),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_459),
.B(n_449),
.C(n_386),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_462),
.B(n_463),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_454),
.A2(n_187),
.B(n_149),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_465),
.A2(n_464),
.B1(n_460),
.B2(n_206),
.Y(n_466)
);

OA21x2_ASAP7_75t_SL g467 ( 
.A1(n_466),
.A2(n_218),
.B(n_159),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_171),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_164),
.Y(n_469)
);


endmodule