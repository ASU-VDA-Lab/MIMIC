module real_jpeg_32984_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_0),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_0),
.Y(n_400)
);

OAI211xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_19),
.C(n_525),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_18),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_2),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_102),
.B1(n_109),
.B2(n_110),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_3),
.A2(n_109),
.B1(n_141),
.B2(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_3),
.A2(n_109),
.B1(n_323),
.B2(n_325),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_3),
.A2(n_109),
.B1(n_507),
.B2(n_513),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_4),
.Y(n_360)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_5),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_5),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_6),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_8),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_8),
.A2(n_191),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_8),
.A2(n_178),
.B1(n_191),
.B2(n_280),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_8),
.A2(n_191),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

OAI22x1_ASAP7_75t_L g115 ( 
.A1(n_10),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_10),
.Y(n_119)
);

AO22x2_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_119),
.B1(n_152),
.B2(n_155),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_119),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_10),
.A2(n_119),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_11),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_12),
.A2(n_46),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22x1_ASAP7_75t_SL g215 ( 
.A1(n_12),
.A2(n_46),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_12),
.B(n_295),
.Y(n_294)
);

OAI32xp33_ASAP7_75t_L g354 ( 
.A1(n_12),
.A2(n_355),
.A3(n_361),
.B1(n_363),
.B2(n_367),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_12),
.B(n_127),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NAND4xp25_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_20),
.C(n_493),
.D(n_524),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_17),
.B(n_493),
.Y(n_528)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_20),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_250),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_222),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_23),
.B(n_222),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_123),
.C(n_182),
.Y(n_23)
);

INVxp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_25),
.B(n_124),
.Y(n_474)
);

XNOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_80),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_78),
.B2(n_79),
.Y(n_26)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_27),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_SL g283 ( 
.A(n_27),
.B(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_27),
.A2(n_78),
.B1(n_284),
.B2(n_342),
.Y(n_341)
);

AO21x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_37),
.B(n_39),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_SL g441 ( 
.A1(n_28),
.A2(n_272),
.B(n_322),
.Y(n_441)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_29),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_29),
.B(n_40),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_29),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_30),
.B(n_46),
.Y(n_413)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_37),
.Y(n_203)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_40),
.B(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21x1_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_72),
.B(n_76),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_77),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_46),
.B(n_197),
.Y(n_268)
);

AOI32xp33_ASAP7_75t_L g284 ( 
.A1(n_46),
.A2(n_285),
.A3(n_288),
.B1(n_293),
.B2(n_294),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_46),
.B(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_46),
.B(n_405),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_47),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_70),
.B(n_71),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_48),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_48),
.B(n_71),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_48),
.B(n_238),
.Y(n_456)
);

NOR2x1p5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_55),
.B2(n_58),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_51),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_51),
.Y(n_241)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_54),
.Y(n_309)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_54),
.Y(n_318)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_57),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_57),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_57),
.Y(n_313)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_60),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_60),
.B(n_187),
.Y(n_333)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_71),
.B(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_75),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_76),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_78),
.A2(n_81),
.B1(n_224),
.B2(n_469),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_80),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_81),
.Y(n_469)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_101),
.B1(n_114),
.B2(n_115),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_82),
.B(n_115),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_82),
.A2(n_114),
.B(n_176),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_82),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_82),
.B(n_176),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_93),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_91),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_86),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_90),
.Y(n_375)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_92),
.Y(n_296)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_97),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_97),
.Y(n_366)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_101),
.B(n_114),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_114),
.B(n_279),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_114),
.B(n_115),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_114),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_173),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_125),
.B(n_173),
.Y(n_249)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_148),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_139),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_127),
.B(n_151),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_L g235 ( 
.A(n_127),
.B(n_151),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_127),
.B(n_259),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_127),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_127),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AO21x2_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_161),
.B(n_169),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_128)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_129),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_140),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_146),
.A2(n_315),
.B(n_319),
.Y(n_314)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_148),
.B(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g522 ( 
.A(n_149),
.B(n_232),
.C(n_521),
.Y(n_522)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_150),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_159),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_154),
.Y(n_261)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_154),
.Y(n_305)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_159),
.B(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_215),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_161),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_164),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_174),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_174),
.B(n_200),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_175),
.B(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_180),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_181),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_183),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_198),
.C(n_212),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_185),
.B(n_213),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_195),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_186),
.B(n_237),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_197),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_199),
.B(n_467),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_201),
.B(n_449),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_202),
.B(n_388),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_204),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_204),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_209),
.Y(n_324)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2x1p5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_214),
.Y(n_345)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_215),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_215),
.A2(n_234),
.B(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_221),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_223),
.B(n_248),
.C(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_248),
.B2(n_249),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_229),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_236),
.B1(n_246),
.B2(n_247),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_232),
.B(n_330),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_232),
.B(n_330),
.C(n_332),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_232),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_232),
.A2(n_519),
.B(n_522),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_233),
.Y(n_500)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_236),
.A2(n_246),
.B1(n_503),
.B2(n_504),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_245),
.Y(n_236)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_245),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_246),
.B(n_500),
.C(n_501),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_483),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_425),
.B(n_482),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_334),
.B(n_424),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_297),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_254),
.B(n_297),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_277),
.C(n_283),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_255),
.A2(n_256),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_267),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_276),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_258),
.B(n_436),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B(n_276),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_268),
.B(n_269),
.Y(n_300)
);

NOR2x1p5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_270),
.Y(n_409)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g406 ( 
.A(n_272),
.B(n_388),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_273),
.Y(n_321)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_283),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_278),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_328),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_299),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_301),
.B(n_328),
.C(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_320),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_302),
.B(n_320),
.Y(n_431)
);

OAI31xp33_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_306),
.A3(n_310),
.B(n_314),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_333),
.B(n_456),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_349),
.B(n_423),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_336),
.B(n_339),
.Y(n_423)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.C(n_346),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_341),
.B(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_343),
.A2(n_344),
.B1(n_346),
.B2(n_347),
.Y(n_419)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_378),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_417),
.B(n_422),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_395),
.B(n_416),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_379),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_352),
.B(n_379),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_376),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_353),
.A2(n_354),
.B1(n_376),
.B2(n_377),
.Y(n_401)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_378),
.B(n_385),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_386),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_387),
.C(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI21x1_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_402),
.B(n_415),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_401),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_401),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_409),
.Y(n_408)
);

BUFx4f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_407),
.B(n_414),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_406),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_420),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_463),
.C(n_475),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_458),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_427),
.B(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_443),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_428),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_439),
.C(n_440),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_429),
.B(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_438),
.C(n_447),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_434),
.B1(n_435),
.B2(n_438),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_435),
.Y(n_438)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_436),
.Y(n_521)
);

XOR2x1_ASAP7_75t_SL g462 ( 
.A(n_439),
.B(n_440),
.Y(n_462)
);

XOR2x2_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_442),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_450),
.B2(n_451),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_477),
.C(n_479),
.Y(n_476)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_457),
.C(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_456),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_461),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_461),
.Y(n_486)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_463),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_473),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_464),
.B(n_473),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.C(n_470),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_468),
.Y(n_481)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_481),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_475),
.A2(n_485),
.B(n_487),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_480),
.Y(n_491)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_484),
.A2(n_490),
.B(n_492),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_523),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NOR2x1_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_496),
.B(n_498),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_518),
.Y(n_504)
);

OA21x2_ASAP7_75t_SL g505 ( 
.A1(n_506),
.A2(n_516),
.B(n_517),
.Y(n_505)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx3_ASAP7_75t_SL g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx6_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_524),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_527),
.B(n_528),
.Y(n_525)
);


endmodule