module fake_jpeg_31649_n_52 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_52);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_0),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_39),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_R g38 ( 
.A(n_32),
.B(n_31),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_32),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_48),
.C(n_41),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_30),
.C(n_29),
.Y(n_48)
);

OAI221xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_4),
.B2(n_8),
.C(n_9),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_45),
.C(n_7),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_14),
.B(n_15),
.Y(n_52)
);


endmodule