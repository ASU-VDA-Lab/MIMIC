module fake_jpeg_20739_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_58),
.Y(n_107)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_20),
.B1(n_22),
.B2(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_47),
.B1(n_40),
.B2(n_35),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_96),
.B1(n_40),
.B2(n_31),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_69),
.B(n_77),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_75),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_43),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_87),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_76),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_79),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_81),
.Y(n_132)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_22),
.B1(n_20),
.B2(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_88),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_32),
.B(n_30),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_38),
.C(n_41),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_26),
.B1(n_45),
.B2(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_95),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_92),
.B(n_94),
.Y(n_140)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_44),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_57),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_40),
.B1(n_25),
.B2(n_26),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_32),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_21),
.Y(n_142)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_25),
.B1(n_26),
.B2(n_48),
.Y(n_103)
);

OAI22x1_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_21),
.B1(n_39),
.B2(n_40),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_50),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx5_ASAP7_75t_SL g136 ( 
.A(n_109),
.Y(n_136)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_120),
.B1(n_133),
.B2(n_80),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_31),
.B1(n_44),
.B2(n_42),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_72),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_90),
.B(n_21),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_27),
.B1(n_34),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_80),
.B1(n_21),
.B2(n_100),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_38),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_75),
.B1(n_70),
.B2(n_72),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_146),
.B1(n_155),
.B2(n_166),
.Y(n_184)
);

NAND2x1p5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_86),
.Y(n_145)
);

AND2x4_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_136),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_107),
.B1(n_90),
.B2(n_110),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_87),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_147),
.A2(n_153),
.B(n_156),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_71),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_152),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_71),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_41),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_167),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_74),
.B1(n_106),
.B2(n_105),
.Y(n_155)
);

XOR2x2_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_41),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_157),
.A2(n_171),
.B1(n_162),
.B2(n_173),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_41),
.C(n_91),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_143),
.C(n_99),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_34),
.B(n_27),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_161),
.B(n_0),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_165),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_21),
.B(n_39),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_163),
.B1(n_170),
.B2(n_116),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_95),
.B1(n_93),
.B2(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_132),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_83),
.B1(n_44),
.B2(n_42),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_140),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_111),
.A2(n_44),
.B1(n_42),
.B2(n_80),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_80),
.B(n_99),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_143),
.B(n_18),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_24),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_119),
.C(n_139),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_18),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_113),
.B1(n_136),
.B2(n_141),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_178),
.A2(n_196),
.B(n_197),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_168),
.A2(n_113),
.B1(n_129),
.B2(n_141),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_182),
.B1(n_206),
.B2(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_125),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_200),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_164),
.B1(n_145),
.B2(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_192),
.B1(n_194),
.B2(n_201),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_147),
.B1(n_163),
.B2(n_164),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_203),
.B1(n_17),
.B2(n_16),
.Y(n_227)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_42),
.B1(n_115),
.B2(n_39),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_191),
.Y(n_219)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_126),
.B(n_117),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_126),
.B1(n_117),
.B2(n_116),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_122),
.B1(n_129),
.B2(n_115),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_172),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_115),
.B(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_148),
.B1(n_152),
.B2(n_169),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_161),
.B(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_147),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_204),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_158),
.A2(n_18),
.B1(n_17),
.B2(n_24),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_153),
.B1(n_151),
.B2(n_157),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_207),
.A2(n_229),
.B(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_153),
.C(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_200),
.C(n_217),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_218),
.B1(n_220),
.B2(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_233),
.B1(n_227),
.B2(n_225),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_223),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_216),
.B(n_221),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_167),
.B1(n_154),
.B2(n_150),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_153),
.B1(n_167),
.B2(n_11),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_24),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_222),
.B(n_176),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_227),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_226),
.Y(n_251)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_179),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_178),
.B1(n_193),
.B2(n_198),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_178),
.B(n_174),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_16),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_209),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_199),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_248),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_245),
.B(n_254),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_188),
.B(n_189),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_191),
.B1(n_190),
.B2(n_182),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_230),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_191),
.B(n_175),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_197),
.B(n_179),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_210),
.C(n_208),
.Y(n_263)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_176),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_208),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_257),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_235),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_229),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_262),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_266),
.C(n_271),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_220),
.C(n_231),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_207),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_273),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_275),
.B1(n_1),
.B2(n_2),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_224),
.C(n_205),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_256),
.B(n_237),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_230),
.B1(n_183),
.B2(n_211),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_246),
.A2(n_232),
.B1(n_255),
.B2(n_254),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_255),
.B1(n_251),
.B2(n_241),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_233),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_242),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_244),
.C(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.C(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_211),
.C(n_228),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_283),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_238),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_291),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_293),
.B1(n_267),
.B2(n_261),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_250),
.B1(n_243),
.B2(n_241),
.Y(n_288)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_271),
.A2(n_190),
.B1(n_239),
.B2(n_16),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_272),
.B1(n_260),
.B2(n_274),
.Y(n_299)
);

FAx1_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_1),
.CI(n_2),
.CON(n_291),
.SN(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_13),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_277),
.C(n_264),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_268),
.A2(n_11),
.B1(n_9),
.B2(n_3),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_303),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_306),
.B1(n_291),
.B2(n_294),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_263),
.B1(n_269),
.B2(n_3),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_269),
.B(n_2),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_283),
.C(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_310),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_282),
.C(n_287),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_294),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_316),
.C(n_300),
.Y(n_319)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_287),
.C(n_291),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_298),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_321),
.B(n_323),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_320),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_296),
.C(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_305),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_303),
.B(n_314),
.C(n_311),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_326),
.B(n_327),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_1),
.B(n_4),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_317),
.C(n_4),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_329),
.B(n_5),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_1),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_5),
.B(n_6),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_5),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_8),
.Y(n_335)
);


endmodule