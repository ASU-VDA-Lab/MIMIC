module real_aes_2101_n_15 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_15);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_15;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_55;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_53;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_54;
wire n_51;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_0), .Y(n_31) );
AOI322xp5_ASAP7_75t_SL g35 ( .A1(n_1), .A2(n_11), .A3(n_18), .B1(n_36), .B2(n_37), .C1(n_48), .C2(n_54), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_2), .Y(n_25) );
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_3), .B(n_6), .C(n_24), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_4), .Y(n_24) );
NAND3xp33_ASAP7_75t_SL g27 ( .A(n_5), .B(n_28), .C(n_29), .Y(n_27) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_5), .B(n_22), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_7), .Y(n_30) );
NOR2xp33_ASAP7_75t_R g47 ( .A(n_7), .B(n_9), .Y(n_47) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_8), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g45 ( .A(n_8), .B(n_46), .Y(n_45) );
NAND2xp33_ASAP7_75t_SL g17 ( .A(n_9), .B(n_18), .Y(n_17) );
NAND2xp33_ASAP7_75t_SL g32 ( .A(n_9), .B(n_33), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g36 ( .A(n_9), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_10), .Y(n_16) );
INVx3_ASAP7_75t_L g53 ( .A(n_12), .Y(n_53) );
CKINVDCx20_ASAP7_75t_R g26 ( .A(n_13), .Y(n_26) );
NAND2xp33_ASAP7_75t_SL g34 ( .A(n_13), .B(n_21), .Y(n_34) );
NOR2xp33_ASAP7_75t_R g29 ( .A(n_14), .B(n_30), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g43 ( .A(n_14), .Y(n_43) );
OAI221xp5_ASAP7_75t_R g15 ( .A1(n_16), .A2(n_17), .B1(n_31), .B2(n_32), .C(n_35), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
OR2x2_ASAP7_75t_L g19 ( .A(n_20), .B(n_27), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g20 ( .A(n_21), .B(n_26), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
NAND2xp33_ASAP7_75t_SL g22 ( .A(n_23), .B(n_25), .Y(n_22) );
NAND2xp33_ASAP7_75t_SL g40 ( .A(n_26), .B(n_41), .Y(n_40) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_27), .B(n_34), .Y(n_33) );
NAND2xp33_ASAP7_75t_SL g55 ( .A(n_33), .B(n_36), .Y(n_55) );
CKINVDCx20_ASAP7_75t_R g37 ( .A(n_38), .Y(n_37) );
NAND2xp33_ASAP7_75t_SL g38 ( .A(n_39), .B(n_42), .Y(n_38) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_43), .B(n_44), .Y(n_42) );
CKINVDCx20_ASAP7_75t_R g44 ( .A(n_45), .Y(n_44) );
CKINVDCx14_ASAP7_75t_R g46 ( .A(n_47), .Y(n_46) );
CKINVDCx20_ASAP7_75t_R g48 ( .A(n_49), .Y(n_48) );
CKINVDCx20_ASAP7_75t_R g49 ( .A(n_50), .Y(n_49) );
HB1xp67_ASAP7_75t_L g50 ( .A(n_51), .Y(n_50) );
INVx2_ASAP7_75t_L g51 ( .A(n_52), .Y(n_51) );
HB1xp67_ASAP7_75t_L g52 ( .A(n_53), .Y(n_52) );
INVx1_ASAP7_75t_SL g54 ( .A(n_55), .Y(n_54) );
endmodule