module fake_jpeg_31894_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_58),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_42),
.C(n_41),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_3),
.C(n_4),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_72),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_48),
.B(n_18),
.C(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_16),
.B1(n_38),
.B2(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_3),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_47),
.B1(n_51),
.B2(n_45),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_102)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_51),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_1),
.B(n_2),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_83),
.C(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_15),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_6),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_86),
.B(n_5),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_14),
.B1(n_33),
.B2(n_32),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_39),
.B1(n_30),
.B2(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_99),
.C(n_100),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_82),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_7),
.C(n_8),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_7),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_13),
.C(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_110),
.B(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_114),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_95),
.A3(n_90),
.B1(n_99),
.B2(n_102),
.C1(n_9),
.C2(n_11),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_108),
.B(n_107),
.C(n_103),
.D(n_104),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_111),
.B1(n_116),
.B2(n_88),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_105),
.C(n_112),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_112),
.A3(n_93),
.B1(n_17),
.B2(n_21),
.C1(n_25),
.C2(n_12),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_120),
.Y(n_121)
);


endmodule