module fake_netlist_5_2144_n_1995 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1995);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1995;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_3),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_195),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_90),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_60),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_50),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_114),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_24),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_128),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_122),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_93),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_22),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_1),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_45),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_91),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_150),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_98),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_125),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_60),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_16),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_107),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_192),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_23),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_112),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_111),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_95),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_121),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_133),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_30),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_129),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_131),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_87),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_126),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_45),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_141),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_21),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_51),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_80),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_21),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_74),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_25),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_61),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_69),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_6),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_62),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_20),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_75),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_110),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_136),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_17),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_104),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_139),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_196),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_78),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_169),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_77),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_152),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_47),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_163),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_120),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_145),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_113),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_18),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_144),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_85),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_81),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_46),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_119),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_38),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_162),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_44),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_132),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_33),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_146),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_53),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_156),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_148),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_40),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_56),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_89),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_38),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_137),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_168),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_52),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_179),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_47),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_124),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_69),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_184),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_188),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_191),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_82),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_170),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_23),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_11),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_57),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_72),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_43),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_36),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_58),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_8),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_155),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_50),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_55),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_67),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_29),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_2),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_59),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_159),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_2),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_13),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_70),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_8),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_116),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_12),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_65),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_167),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_178),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_142),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_42),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_46),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_35),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_83),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_62),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_3),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_108),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_193),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_84),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_97),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_40),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_127),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_172),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_32),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_79),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_20),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_6),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_33),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_100),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_73),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_31),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_1),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_160),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_103),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_165),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_14),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_27),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_37),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_34),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_41),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_171),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_189),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_88),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_64),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_109),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_28),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_26),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_30),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_96),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_183),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_49),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_22),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_153),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_106),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_4),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_17),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_26),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_44),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_61),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_41),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_94),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_65),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_187),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_7),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_67),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_31),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_28),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_64),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_271),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_203),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_237),
.B(n_0),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_235),
.B(n_0),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_207),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_228),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_199),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_209),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_203),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_210),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_206),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_216),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_260),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_218),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_222),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_231),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_229),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_232),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_271),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_246),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_282),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_323),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_242),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_260),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_247),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_237),
.B(n_206),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_290),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_208),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_355),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_235),
.B(n_5),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_333),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_208),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_213),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_213),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_252),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_219),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_219),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_333),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_298),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_221),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_221),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_226),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_226),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_201),
.B(n_5),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_230),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_321),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_230),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_258),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_239),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_373),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_239),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_243),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_200),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_212),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_259),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_212),
.B(n_7),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_355),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_220),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_275),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_262),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_262),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_243),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_202),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_253),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_204),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_287),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_263),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_289),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_253),
.B(n_10),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_231),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_231),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_211),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_291),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_268),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_268),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_293),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g483 ( 
.A(n_220),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_249),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_272),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_383),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_296),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_214),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_215),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_269),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_263),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_297),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_269),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_304),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_217),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_224),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_273),
.B(n_10),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_462),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_496),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_401),
.B(n_322),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_458),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_472),
.B(n_318),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_428),
.B(n_225),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_486),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_486),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_415),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_486),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_462),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_418),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_418),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_397),
.B(n_227),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_399),
.B(n_205),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_421),
.B(n_201),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_426),
.B(n_257),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_426),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_427),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

NAND2x1_ASAP7_75t_L g529 ( 
.A(n_449),
.B(n_272),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_432),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_417),
.B(n_233),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_318),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_434),
.B(n_234),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_403),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_465),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_466),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_466),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_482),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_482),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_442),
.B(n_405),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_484),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_407),
.B(n_356),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_487),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_487),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_424),
.B(n_223),
.Y(n_551)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_461),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_431),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_402),
.B(n_349),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_409),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_435),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

AND2x2_ASAP7_75t_SL g559 ( 
.A(n_474),
.B(n_257),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_440),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_441),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_444),
.B(n_266),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_445),
.B(n_356),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_446),
.B(n_266),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_447),
.B(n_450),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_452),
.B(n_236),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_412),
.B(n_231),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_454),
.B(n_238),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_456),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_430),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_457),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_467),
.B(n_240),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_480),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_492),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_495),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_461),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_553),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_516),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_521),
.B(n_408),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_553),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_403),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_509),
.B(n_468),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_SL g586 ( 
.A(n_578),
.B(n_438),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_559),
.A2(n_499),
.B1(n_433),
.B2(n_400),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_525),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_555),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_516),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_553),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_552),
.B(n_578),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_516),
.Y(n_593)
);

BUFx8_ASAP7_75t_SL g594 ( 
.A(n_504),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_538),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_507),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_517),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_507),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_509),
.B(n_404),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_507),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_551),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_517),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_507),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_517),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_517),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_538),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_578),
.B(n_476),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_551),
.B(n_475),
.Y(n_609)
);

INVxp33_ASAP7_75t_SL g610 ( 
.A(n_503),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_519),
.B(n_470),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_518),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_552),
.A2(n_276),
.B1(n_283),
.B2(n_273),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_518),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_538),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_557),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_529),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_518),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_500),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_503),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_503),
.B(n_554),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_500),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_530),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_500),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_578),
.B(n_277),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_519),
.B(n_477),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_518),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_552),
.B(n_506),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_536),
.B(n_404),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_558),
.Y(n_632)
);

INVx8_ASAP7_75t_L g633 ( 
.A(n_525),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_558),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_559),
.A2(n_249),
.B1(n_254),
.B2(n_250),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_520),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_530),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_559),
.A2(n_567),
.B1(n_390),
.B2(n_392),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_552),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_554),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_516),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_532),
.B(n_490),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_560),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_520),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_516),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_532),
.B(n_406),
.Y(n_647)
);

INVxp33_ASAP7_75t_L g648 ( 
.A(n_554),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_560),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_530),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_567),
.B(n_491),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_543),
.B(n_483),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_552),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_529),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_529),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_561),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_557),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_559),
.A2(n_250),
.B1(n_261),
.B2(n_254),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_552),
.A2(n_543),
.B1(n_533),
.B2(n_506),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_574),
.Y(n_662)
);

CKINVDCx6p67_ASAP7_75t_R g663 ( 
.A(n_536),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_520),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_511),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_535),
.B(n_497),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_516),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_498),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_566),
.B(n_406),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_506),
.A2(n_261),
.B1(n_278),
.B2(n_267),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_570),
.B(n_410),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_500),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_500),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_557),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_533),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_557),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_574),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_502),
.A2(n_570),
.B1(n_579),
.B2(n_411),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_504),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_566),
.B(n_568),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_533),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_568),
.B(n_410),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_562),
.A2(n_352),
.B1(n_344),
.B2(n_339),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_575),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_530),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_575),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_562),
.B(n_564),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_516),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_562),
.A2(n_352),
.B1(n_344),
.B2(n_339),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_502),
.B(n_411),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_577),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_562),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_577),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_530),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_546),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_530),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_572),
.B(n_413),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_523),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_530),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_501),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_501),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_579),
.B(n_416),
.C(n_413),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_523),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_508),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_579),
.A2(n_494),
.B1(n_489),
.B2(n_416),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_557),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_530),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_523),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_579),
.B(n_422),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_523),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_524),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_524),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_524),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_562),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_524),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_527),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_572),
.B(n_422),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_511),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_508),
.B(n_425),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_557),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_512),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_511),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_512),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_557),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_527),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_546),
.B(n_463),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_562),
.A2(n_368),
.B1(n_331),
.B2(n_326),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_513),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_546),
.B(n_419),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_557),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_527),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_601),
.B(n_425),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_640),
.B(n_241),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_584),
.B(n_439),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_680),
.B(n_569),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_651),
.B(n_420),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_632),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_675),
.B(n_569),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_619),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_640),
.B(n_244),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_675),
.B(n_569),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_681),
.B(n_569),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_635),
.A2(n_278),
.B1(n_281),
.B2(n_267),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_681),
.B(n_439),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_R g745 ( 
.A(n_679),
.B(n_429),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_661),
.B(n_569),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_659),
.B(n_569),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_599),
.B(n_647),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_653),
.B(n_453),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_653),
.B(n_453),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_592),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_726),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_659),
.B(n_569),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_608),
.B(n_460),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_626),
.B(n_245),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_671),
.B(n_460),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_659),
.B(n_569),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_669),
.B(n_464),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_632),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_654),
.B(n_272),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_660),
.A2(n_281),
.B1(n_317),
.B2(n_285),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_634),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_626),
.B(n_251),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_639),
.A2(n_354),
.B1(n_364),
.B2(n_327),
.Y(n_764)
);

AND2x6_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_276),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_697),
.B(n_464),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_L g767 ( 
.A(n_626),
.B(n_587),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_616),
.Y(n_768)
);

OAI221xp5_ASAP7_75t_L g769 ( 
.A1(n_670),
.A2(n_565),
.B1(n_485),
.B2(n_256),
.C(n_285),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_582),
.B(n_473),
.C(n_471),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_585),
.B(n_471),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_611),
.B(n_473),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_L g773 ( 
.A(n_663),
.B(n_478),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_634),
.Y(n_774)
);

NOR2x2_ASAP7_75t_L g775 ( 
.A(n_639),
.B(n_277),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_607),
.B(n_571),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_627),
.B(n_478),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_607),
.B(n_571),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_626),
.A2(n_368),
.B1(n_375),
.B2(n_379),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_616),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_654),
.B(n_272),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_644),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_626),
.A2(n_375),
.B1(n_379),
.B2(n_396),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_615),
.B(n_571),
.Y(n_784)
);

OAI221xp5_ASAP7_75t_L g785 ( 
.A1(n_683),
.A2(n_565),
.B1(n_396),
.B2(n_317),
.C(n_331),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_643),
.B(n_481),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_608),
.B(n_481),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_622),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_695),
.A2(n_564),
.B(n_337),
.C(n_522),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_644),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_592),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_615),
.B(n_571),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_626),
.B(n_264),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_695),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_580),
.B(n_571),
.Y(n_795)
);

O2A1O1Ixp5_ASAP7_75t_L g796 ( 
.A1(n_622),
.A2(n_672),
.B(n_673),
.C(n_625),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_625),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_580),
.B(n_571),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_583),
.B(n_571),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_583),
.B(n_571),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_591),
.B(n_649),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_654),
.B(n_272),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_591),
.B(n_556),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_726),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_654),
.B(n_564),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_649),
.Y(n_806)
);

NOR3xp33_ASAP7_75t_L g807 ( 
.A(n_609),
.B(n_494),
.C(n_489),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_666),
.B(n_361),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_613),
.A2(n_564),
.B(n_563),
.C(n_576),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_652),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_652),
.B(n_556),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_657),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_657),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_626),
.B(n_265),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_668),
.B(n_563),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_662),
.B(n_556),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_665),
.A2(n_510),
.B(n_505),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_617),
.B(n_564),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_702),
.B(n_563),
.C(n_307),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_662),
.B(n_556),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_677),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_594),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_677),
.B(n_573),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_684),
.B(n_573),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_673),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_630),
.A2(n_443),
.B1(n_451),
.B2(n_455),
.Y(n_826)
);

INVx8_ASAP7_75t_L g827 ( 
.A(n_592),
.Y(n_827)
);

OAI22xp33_ASAP7_75t_L g828 ( 
.A1(n_592),
.A2(n_326),
.B1(n_386),
.B2(n_300),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_684),
.B(n_686),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_686),
.B(n_573),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_589),
.B(n_534),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_690),
.B(n_270),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_592),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_691),
.B(n_573),
.Y(n_834)
);

BUFx5_ASAP7_75t_L g835 ( 
.A(n_617),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_691),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_693),
.B(n_576),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_630),
.A2(n_358),
.B1(n_338),
.B2(n_283),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_678),
.B(n_705),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_693),
.B(n_576),
.Y(n_840)
);

AOI22x1_ASAP7_75t_L g841 ( 
.A1(n_596),
.A2(n_337),
.B1(n_301),
.B2(n_288),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_700),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_589),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_671),
.B(n_534),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_SL g845 ( 
.A(n_655),
.B(n_288),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_629),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_719),
.B(n_537),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_700),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_630),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_701),
.B(n_576),
.Y(n_850)
);

AOI221x1_ASAP7_75t_L g851 ( 
.A1(n_596),
.A2(n_255),
.B1(n_363),
.B2(n_300),
.C(n_301),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_630),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_655),
.B(n_564),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_701),
.B(n_522),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_704),
.B(n_522),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_704),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_630),
.A2(n_248),
.B1(n_342),
.B2(n_357),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_721),
.B(n_522),
.Y(n_858)
);

O2A1O1Ixp5_ASAP7_75t_L g859 ( 
.A1(n_598),
.A2(n_522),
.B(n_526),
.C(n_531),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_721),
.B(n_522),
.Y(n_860)
);

AO221x1_ASAP7_75t_L g861 ( 
.A1(n_629),
.A2(n_338),
.B1(n_305),
.B2(n_346),
.C(n_363),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_723),
.B(n_513),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_663),
.B(n_537),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_709),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_655),
.Y(n_865)
);

BUFx5_ASAP7_75t_L g866 ( 
.A(n_656),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_656),
.B(n_305),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_597),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_723),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_631),
.B(n_313),
.C(n_306),
.Y(n_870)
);

NOR2xp67_ASAP7_75t_L g871 ( 
.A(n_598),
.B(n_539),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_682),
.A2(n_310),
.B1(n_274),
.B2(n_280),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_728),
.B(n_544),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_620),
.B(n_315),
.C(n_314),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_717),
.B(n_319),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_729),
.B(n_279),
.Y(n_876)
);

O2A1O1Ixp5_ASAP7_75t_L g877 ( 
.A1(n_600),
.A2(n_526),
.B(n_531),
.C(n_308),
.Y(n_877)
);

OAI22x1_ASAP7_75t_L g878 ( 
.A1(n_621),
.A2(n_380),
.B1(n_359),
.B2(n_360),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_687),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_687),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_586),
.B(n_320),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_595),
.B(n_544),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_687),
.B(n_308),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_595),
.B(n_544),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_656),
.B(n_284),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_595),
.B(n_544),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_687),
.Y(n_887)
);

INVx8_ASAP7_75t_L g888 ( 
.A(n_633),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_692),
.B(n_286),
.Y(n_889)
);

O2A1O1Ixp5_ASAP7_75t_L g890 ( 
.A1(n_600),
.A2(n_526),
.B(n_531),
.C(n_358),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_604),
.B(n_539),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_603),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_604),
.A2(n_303),
.B1(n_292),
.B2(n_295),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_604),
.B(n_324),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_603),
.B(n_325),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_722),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_602),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_843),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_805),
.A2(n_720),
.B(n_637),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_839),
.A2(n_689),
.B(n_727),
.C(n_378),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_805),
.A2(n_720),
.B(n_637),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_735),
.A2(n_720),
.B(n_637),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_748),
.B(n_718),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_835),
.B(n_692),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_748),
.B(n_718),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_756),
.B(n_641),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_818),
.A2(n_720),
.B(n_637),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_808),
.A2(n_346),
.B(n_348),
.C(n_378),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_853),
.A2(n_650),
.B(n_624),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_883),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_853),
.A2(n_650),
.B(n_624),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_835),
.B(n_692),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_888),
.A2(n_650),
.B(n_624),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_808),
.B(n_718),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_815),
.B(n_718),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_888),
.A2(n_650),
.B(n_624),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_732),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_815),
.A2(n_692),
.B1(n_714),
.B2(n_722),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_771),
.B(n_722),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_739),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_831),
.B(n_648),
.Y(n_921)
);

OAI321xp33_ASAP7_75t_L g922 ( 
.A1(n_839),
.A2(n_348),
.A3(n_547),
.B1(n_549),
.B2(n_541),
.C(n_540),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_788),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_734),
.B(n_865),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_772),
.A2(n_786),
.B(n_777),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_771),
.B(n_610),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_888),
.A2(n_694),
.B(n_685),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_734),
.B(n_714),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_865),
.B(n_714),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_772),
.B(n_714),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_SL g931 ( 
.A1(n_789),
.A2(n_581),
.B(n_590),
.C(n_593),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_777),
.A2(n_707),
.B1(n_581),
.B2(n_590),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_822),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_752),
.A2(n_698),
.B(n_708),
.C(n_710),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_859),
.A2(n_731),
.B(n_605),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_768),
.A2(n_694),
.B(n_685),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_804),
.A2(n_794),
.B(n_767),
.C(n_838),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_780),
.A2(n_694),
.B(n_685),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_796),
.A2(n_731),
.B(n_605),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_797),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_786),
.B(n_581),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_746),
.A2(n_694),
.B(n_685),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_791),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_758),
.B(n_329),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_794),
.B(n_581),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_745),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_758),
.B(n_766),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_747),
.A2(n_699),
.B(n_696),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_753),
.A2(n_731),
.B(n_605),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_SL g950 ( 
.A1(n_883),
.A2(n_540),
.B(n_541),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_766),
.B(n_330),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_791),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_737),
.B(n_590),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_759),
.B(n_590),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_762),
.B(n_593),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_757),
.A2(n_699),
.B(n_696),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_825),
.Y(n_957)
);

AO21x1_ASAP7_75t_L g958 ( 
.A1(n_838),
.A2(n_699),
.B(n_696),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_828),
.A2(n_710),
.B(n_711),
.C(n_712),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_760),
.A2(n_699),
.B(n_696),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_791),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_760),
.A2(n_633),
.B(n_616),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_774),
.B(n_593),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_782),
.B(n_593),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_863),
.B(n_299),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_754),
.B(n_299),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_892),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_846),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_790),
.B(n_623),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_806),
.B(n_623),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_781),
.A2(n_633),
.B(n_616),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_810),
.B(n_623),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_877),
.A2(n_606),
.B(n_602),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_781),
.A2(n_633),
.B(n_616),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_749),
.B(n_332),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_745),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_750),
.B(n_335),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_787),
.B(n_340),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_736),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_751),
.A2(n_623),
.B1(n_642),
.B2(n_688),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_802),
.A2(n_633),
.B(n_616),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_764),
.B(n_341),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_812),
.B(n_642),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_764),
.B(n_343),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_828),
.B(n_365),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_835),
.B(n_658),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_802),
.A2(n_674),
.B(n_658),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_882),
.A2(n_674),
.B(n_658),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_875),
.B(n_367),
.C(n_366),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_813),
.B(n_642),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_890),
.A2(n_741),
.B(n_738),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_884),
.A2(n_674),
.B(n_658),
.Y(n_992)
);

CKINVDCx10_ASAP7_75t_R g993 ( 
.A(n_878),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_886),
.A2(n_674),
.B(n_658),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_829),
.A2(n_711),
.B(n_712),
.C(n_716),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_844),
.B(n_299),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_821),
.B(n_836),
.Y(n_997)
);

AO21x2_ASAP7_75t_L g998 ( 
.A1(n_889),
.A2(n_606),
.B(n_602),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_742),
.A2(n_674),
.B(n_658),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_873),
.A2(n_612),
.B(n_606),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_879),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_854),
.A2(n_676),
.B(n_674),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_842),
.B(n_642),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_848),
.B(n_646),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_855),
.A2(n_860),
.B(n_858),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_791),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_875),
.A2(n_646),
.B(n_667),
.C(n_688),
.Y(n_1007)
);

AO21x1_ASAP7_75t_L g1008 ( 
.A1(n_889),
.A2(n_614),
.B(n_612),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_801),
.A2(n_706),
.B(n_676),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_751),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_743),
.A2(n_761),
.B1(n_785),
.B2(n_783),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_856),
.B(n_646),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_880),
.B(n_547),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_776),
.A2(n_706),
.B(n_676),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_887),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_881),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_881),
.A2(n_646),
.B(n_667),
.C(n_688),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_869),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_778),
.A2(n_614),
.B(n_612),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_784),
.A2(n_706),
.B(n_676),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_792),
.A2(n_896),
.B(n_740),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_809),
.A2(n_618),
.B(n_614),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_835),
.B(n_676),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_744),
.B(n_372),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_896),
.A2(n_676),
.B(n_706),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_826),
.B(n_621),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_833),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_847),
.B(n_667),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_864),
.B(n_770),
.Y(n_1029)
);

NOR2xp67_ASAP7_75t_L g1030 ( 
.A(n_819),
.B(n_549),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_835),
.B(n_706),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_835),
.B(n_667),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_876),
.A2(n_393),
.B(n_376),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_891),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_733),
.A2(n_724),
.B(n_706),
.Y(n_1035)
);

AND2x2_ASAP7_75t_SL g1036 ( 
.A(n_743),
.B(n_724),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_833),
.A2(n_730),
.B(n_724),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_866),
.B(n_688),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_827),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_866),
.B(n_707),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_891),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_832),
.B(n_384),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_866),
.B(n_707),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_827),
.B(n_540),
.Y(n_1044)
);

NOR2xp67_ASAP7_75t_L g1045 ( 
.A(n_894),
.B(n_309),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_866),
.B(n_707),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_849),
.B(n_588),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_811),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_866),
.B(n_618),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_885),
.A2(n_628),
.B(n_725),
.C(n_716),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_773),
.B(n_526),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_866),
.B(n_895),
.Y(n_1052)
);

AOI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_894),
.A2(n_395),
.B(n_394),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_849),
.A2(n_724),
.B(n_730),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_895),
.B(n_618),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_795),
.A2(n_628),
.B(n_725),
.C(n_636),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_816),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_769),
.A2(n_636),
.B(n_716),
.C(n_715),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_775),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_798),
.A2(n_628),
.B(n_725),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_827),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_852),
.A2(n_544),
.B(n_548),
.C(n_715),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_852),
.A2(n_730),
.B(n_724),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_862),
.B(n_387),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_872),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_761),
.B(n_871),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_857),
.A2(n_548),
.B(n_636),
.C(n_715),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_765),
.B(n_638),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_820),
.B(n_724),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_807),
.B(n_388),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_765),
.A2(n_389),
.B1(n_311),
.B2(n_312),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_765),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_823),
.A2(n_730),
.B(n_588),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_765),
.B(n_638),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_799),
.A2(n_638),
.B(n_713),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_765),
.B(n_645),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_867),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_800),
.A2(n_645),
.B(n_713),
.Y(n_1078)
);

BUFx2_ASAP7_75t_SL g1079 ( 
.A(n_867),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_874),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_824),
.B(n_316),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_L g1082 ( 
.A(n_830),
.B(n_526),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_929),
.A2(n_814),
.B(n_755),
.Y(n_1083)
);

OR2x6_ASAP7_75t_L g1084 ( 
.A(n_1039),
.B(n_834),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_921),
.B(n_870),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1052),
.A2(n_1005),
.B(n_912),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_925),
.A2(n_837),
.B(n_840),
.C(n_850),
.Y(n_1087)
);

BUFx8_ASAP7_75t_SL g1088 ( 
.A(n_933),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_968),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_947),
.B(n_867),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_930),
.B(n_867),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_965),
.B(n_861),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_968),
.Y(n_1093)
);

INVx3_ASAP7_75t_SL g1094 ( 
.A(n_906),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_904),
.A2(n_763),
.B(n_793),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1061),
.B(n_867),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_930),
.B(n_919),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_R g1098 ( 
.A(n_1065),
.B(n_803),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_898),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_904),
.A2(n_817),
.B(n_730),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1018),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1059),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_944),
.A2(n_845),
.B(n_893),
.C(n_868),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_910),
.A2(n_779),
.B1(n_783),
.B2(n_897),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_919),
.B(n_779),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_910),
.A2(n_362),
.B1(n_369),
.B2(n_370),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_946),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_944),
.A2(n_951),
.B(n_937),
.C(n_1042),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1039),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_951),
.B(n_851),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_SL g1111 ( 
.A(n_1077),
.B(n_279),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_926),
.B(n_299),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1016),
.B(n_328),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_926),
.B(n_966),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_917),
.B(n_336),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1053),
.A2(n_548),
.B(n_713),
.C(n_703),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_R g1117 ( 
.A(n_943),
.B(n_345),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1042),
.A2(n_548),
.B(n_377),
.C(n_350),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1064),
.B(n_645),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_1008),
.A2(n_703),
.A3(n_664),
.B(n_528),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1064),
.B(n_664),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_900),
.A2(n_381),
.B(n_351),
.C(n_353),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1039),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_913),
.A2(n_927),
.B(n_916),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_908),
.A2(n_984),
.B(n_982),
.C(n_985),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1036),
.A2(n_371),
.B1(n_347),
.B2(n_382),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_L g1127 ( 
.A(n_982),
.B(n_550),
.C(n_542),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_920),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_914),
.B(n_664),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_986),
.A2(n_1031),
.B(n_1023),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_914),
.B(n_703),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_985),
.A2(n_550),
.B(n_542),
.C(n_531),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_986),
.A2(n_588),
.B(n_511),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1006),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_940),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_924),
.B(n_841),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_984),
.A2(n_550),
.B(n_542),
.C(n_531),
.Y(n_1137)
);

BUFx8_ASAP7_75t_L g1138 ( 
.A(n_1029),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_1039),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1048),
.B(n_542),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1024),
.A2(n_550),
.B(n_527),
.C(n_528),
.Y(n_1141)
);

AOI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_1024),
.A2(n_302),
.B1(n_385),
.B2(n_545),
.C(n_528),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1023),
.A2(n_588),
.B(n_511),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1044),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1044),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1044),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_928),
.A2(n_1011),
.B1(n_905),
.B2(n_903),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1011),
.A2(n_588),
.B1(n_528),
.B2(n_545),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_967),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_978),
.B(n_302),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_979),
.B(n_279),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1077),
.B(n_545),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1006),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_978),
.B(n_302),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_943),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_1077),
.B(n_545),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1057),
.B(n_545),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1080),
.A2(n_515),
.B(n_514),
.C(n_510),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1032),
.A2(n_1038),
.B(n_1021),
.Y(n_1159)
);

AOI211xp5_ASAP7_75t_L g1160 ( 
.A1(n_975),
.A2(n_385),
.B(n_302),
.C(n_391),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1079),
.B(n_545),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_996),
.B(n_279),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1036),
.A2(n_545),
.B1(n_515),
.B2(n_514),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_975),
.A2(n_977),
.B(n_1070),
.C(n_997),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1026),
.B(n_545),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_915),
.B(n_505),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1081),
.B(n_505),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_976),
.B(n_11),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1077),
.B(n_505),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_952),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_936),
.A2(n_510),
.B(n_515),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_977),
.A2(n_514),
.B(n_510),
.C(n_391),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1066),
.A2(n_525),
.B1(n_391),
.B2(n_294),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_989),
.A2(n_391),
.B1(n_294),
.B2(n_385),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1033),
.B(n_385),
.Y(n_1175)
);

INVx8_ASAP7_75t_L g1176 ( 
.A(n_952),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1034),
.B(n_1041),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1001),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1081),
.B(n_1015),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_941),
.A2(n_294),
.B1(n_198),
.B2(n_190),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_961),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_918),
.A2(n_294),
.B1(n_186),
.B2(n_176),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_950),
.A2(n_525),
.B1(n_175),
.B2(n_174),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_945),
.B(n_525),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1010),
.B(n_525),
.Y(n_1185)
);

O2A1O1Ixp5_ASAP7_75t_L g1186 ( 
.A1(n_958),
.A2(n_130),
.B(n_166),
.C(n_157),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1010),
.B(n_1027),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1027),
.B(n_525),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_961),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1013),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_938),
.A2(n_105),
.B(n_154),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1072),
.A2(n_151),
.B1(n_147),
.B2(n_143),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_923),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_899),
.A2(n_101),
.B(n_140),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_957),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_1013),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1030),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1062),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_901),
.A2(n_99),
.B(n_138),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1040),
.A2(n_118),
.B(n_102),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1043),
.A2(n_92),
.B(n_86),
.Y(n_1201)
);

AOI221xp5_ASAP7_75t_L g1202 ( 
.A1(n_922),
.A2(n_15),
.B1(n_19),
.B2(n_25),
.C(n_27),
.Y(n_1202)
);

NAND2xp33_ASAP7_75t_SL g1203 ( 
.A(n_1055),
.B(n_19),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1045),
.B(n_953),
.Y(n_1204)
);

AOI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1069),
.A2(n_525),
.B(n_76),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_954),
.A2(n_525),
.B1(n_71),
.B2(n_34),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_955),
.B(n_29),
.Y(n_1207)
);

NAND2x1_ASAP7_75t_L g1208 ( 
.A(n_1054),
.B(n_525),
.Y(n_1208)
);

NOR3xp33_ASAP7_75t_SL g1209 ( 
.A(n_993),
.B(n_32),
.C(n_35),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1051),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1071),
.B(n_36),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1028),
.B(n_37),
.Y(n_1212)
);

O2A1O1Ixp5_ASAP7_75t_SL g1213 ( 
.A1(n_1069),
.A2(n_39),
.B(n_42),
.C(n_43),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_963),
.B(n_39),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_964),
.A2(n_525),
.B1(n_49),
.B2(n_51),
.Y(n_1215)
);

BUFx8_ASAP7_75t_SL g1216 ( 
.A(n_1068),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_969),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1046),
.A2(n_70),
.B(n_52),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_970),
.B(n_48),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1074),
.B(n_48),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1049),
.A2(n_53),
.B(n_54),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_972),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_902),
.A2(n_68),
.B(n_55),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_983),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_959),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_907),
.A2(n_58),
.B(n_59),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1050),
.A2(n_63),
.B(n_66),
.C(n_942),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_SL g1228 ( 
.A(n_1076),
.B(n_63),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_R g1229 ( 
.A(n_990),
.B(n_66),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1022),
.B(n_932),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1003),
.B(n_1012),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1007),
.A2(n_1067),
.B(n_1017),
.C(n_934),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_909),
.A2(n_911),
.B(n_1058),
.C(n_991),
.Y(n_1233)
);

BUFx4f_ASAP7_75t_L g1234 ( 
.A(n_1047),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_995),
.A2(n_1009),
.B(n_1004),
.C(n_1002),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_998),
.Y(n_1236)
);

OAI22x1_ASAP7_75t_L g1237 ( 
.A1(n_1047),
.A2(n_1082),
.B1(n_931),
.B2(n_998),
.Y(n_1237)
);

OAI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1154),
.A2(n_1108),
.B(n_1112),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1101),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1124),
.A2(n_939),
.B(n_994),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1114),
.B(n_1063),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1233),
.A2(n_1147),
.A3(n_1237),
.B(n_1235),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1086),
.A2(n_949),
.B(n_935),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1234),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1088),
.Y(n_1245)
);

AOI221x1_ASAP7_75t_L g1246 ( 
.A1(n_1225),
.A2(n_980),
.B1(n_992),
.B2(n_988),
.C(n_1035),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1099),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1125),
.A2(n_1037),
.B(n_981),
.C(n_974),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1100),
.A2(n_999),
.B(n_1020),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1093),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1164),
.A2(n_962),
.B(n_971),
.C(n_948),
.Y(n_1251)
);

NAND2xp33_ASAP7_75t_L g1252 ( 
.A(n_1097),
.B(n_973),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1236),
.A2(n_1014),
.A3(n_956),
.B(n_987),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1232),
.A2(n_1000),
.B(n_1078),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_L g1255 ( 
.A(n_1179),
.B(n_1073),
.Y(n_1255)
);

AND2x6_ASAP7_75t_L g1256 ( 
.A(n_1109),
.B(n_1056),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1083),
.A2(n_960),
.B(n_1025),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1159),
.A2(n_1019),
.B(n_1060),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1110),
.A2(n_1230),
.B(n_1087),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1211),
.A2(n_1175),
.B1(n_1150),
.B2(n_1174),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1105),
.B(n_1075),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1130),
.A2(n_1171),
.B(n_1095),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1089),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1094),
.B(n_1102),
.Y(n_1264)
);

NAND3x1_ASAP7_75t_L g1265 ( 
.A(n_1085),
.B(n_1106),
.C(n_1202),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1139),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1122),
.A2(n_1090),
.B(n_1103),
.C(n_1091),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1205),
.A2(n_1163),
.B(n_1133),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1149),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1119),
.A2(n_1121),
.B(n_1167),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1176),
.B(n_1144),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1153),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1160),
.A2(n_1162),
.B(n_1151),
.C(n_1197),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1132),
.A2(n_1227),
.B(n_1116),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1160),
.A2(n_1092),
.B(n_1204),
.C(n_1126),
.Y(n_1275)
);

AOI221xp5_ASAP7_75t_L g1276 ( 
.A1(n_1203),
.A2(n_1115),
.B1(n_1142),
.B2(n_1180),
.C(n_1198),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1217),
.B(n_1222),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1129),
.A2(n_1131),
.B(n_1136),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1163),
.A2(n_1143),
.B(n_1208),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1178),
.Y(n_1280)
);

NAND2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1098),
.B(n_1144),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1118),
.A2(n_1212),
.B(n_1172),
.C(n_1219),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1168),
.A2(n_1113),
.B(n_1226),
.C(n_1223),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1234),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1176),
.B(n_1144),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1107),
.B(n_1196),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1224),
.B(n_1187),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1123),
.B(n_1109),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1231),
.A2(n_1161),
.B(n_1166),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1220),
.A2(n_1214),
.B1(n_1207),
.B2(n_1126),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1194),
.A2(n_1199),
.B(n_1157),
.Y(n_1291)
);

INVx3_ASAP7_75t_SL g1292 ( 
.A(n_1109),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1155),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1134),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1161),
.A2(n_1140),
.B(n_1111),
.Y(n_1295)
);

INVx5_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1141),
.A2(n_1182),
.A3(n_1148),
.B(n_1104),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1111),
.A2(n_1191),
.B(n_1184),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1193),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1137),
.A2(n_1186),
.B(n_1213),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1221),
.A2(n_1218),
.A3(n_1200),
.B(n_1201),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1165),
.B(n_1190),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1192),
.A2(n_1120),
.A3(n_1185),
.B(n_1188),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1190),
.B(n_1177),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1195),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1152),
.A2(n_1156),
.B(n_1169),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1138),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1152),
.A2(n_1156),
.B(n_1169),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1190),
.B(n_1220),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1210),
.B(n_1216),
.Y(n_1310)
);

CKINVDCx6p67_ASAP7_75t_R g1311 ( 
.A(n_1145),
.Y(n_1311)
);

AO32x2_ASAP7_75t_L g1312 ( 
.A1(n_1120),
.A2(n_1228),
.A3(n_1173),
.B1(n_1215),
.B2(n_1127),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1145),
.B(n_1146),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1128),
.B(n_1135),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1181),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1170),
.Y(n_1316)
);

BUFx12f_ASAP7_75t_L g1317 ( 
.A(n_1138),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1084),
.A2(n_1183),
.B(n_1176),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1170),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1106),
.B(n_1096),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1096),
.B(n_1173),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1084),
.A2(n_1145),
.B1(n_1146),
.B2(n_1183),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1206),
.A2(n_1158),
.B(n_1215),
.C(n_1209),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1206),
.A2(n_1084),
.A3(n_1229),
.B(n_1117),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1146),
.B(n_1155),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1155),
.A2(n_1124),
.B(n_1086),
.Y(n_1326)
);

CKINVDCx16_ASAP7_75t_R g1327 ( 
.A(n_1189),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1189),
.A2(n_1124),
.B(n_1086),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1189),
.A2(n_925),
.B(n_1125),
.C(n_947),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_L g1330 ( 
.A(n_1179),
.B(n_1016),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1124),
.A2(n_1100),
.B(n_1159),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1108),
.A2(n_1097),
.B(n_1147),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1114),
.B(n_947),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1125),
.A2(n_925),
.B(n_947),
.C(n_1108),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1097),
.A2(n_947),
.B1(n_1011),
.B2(n_910),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1114),
.B(n_947),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1124),
.A2(n_1100),
.B(n_1159),
.Y(n_1338)
);

AOI221x1_ASAP7_75t_L g1339 ( 
.A1(n_1108),
.A2(n_925),
.B1(n_947),
.B2(n_951),
.C(n_944),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1101),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1108),
.B(n_947),
.C(n_925),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1093),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1114),
.B(n_947),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1097),
.A2(n_947),
.B1(n_925),
.B2(n_1108),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1123),
.B(n_1039),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1101),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1114),
.B(n_947),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1114),
.B(n_947),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1101),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1124),
.A2(n_1100),
.B(n_1159),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1114),
.B(n_947),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1144),
.B(n_1061),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1108),
.A2(n_1097),
.B(n_1147),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1233),
.A2(n_1108),
.A3(n_1147),
.B(n_1237),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_SL g1358 ( 
.A1(n_1108),
.A2(n_947),
.B(n_1125),
.C(n_1225),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1101),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1114),
.B(n_947),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1125),
.A2(n_925),
.B(n_947),
.C(n_1108),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1362)
);

A2O1A1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1125),
.A2(n_925),
.B(n_947),
.C(n_1108),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1088),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1108),
.A2(n_1097),
.B(n_1147),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1114),
.B(n_947),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1124),
.A2(n_1100),
.B(n_1159),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1102),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1088),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1102),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1108),
.A2(n_1097),
.B(n_1147),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1101),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1099),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1097),
.A2(n_947),
.B1(n_925),
.B2(n_1108),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_SL g1378 ( 
.A1(n_1108),
.A2(n_947),
.B(n_1125),
.C(n_1225),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1108),
.A2(n_947),
.B(n_925),
.C(n_808),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1088),
.Y(n_1380)
);

AND2x6_ASAP7_75t_L g1381 ( 
.A(n_1109),
.B(n_791),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1114),
.B(n_947),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1102),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1124),
.A2(n_1100),
.B(n_1159),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1114),
.B(n_947),
.Y(n_1386)
);

NAND2x1_ASAP7_75t_L g1387 ( 
.A(n_1170),
.B(n_849),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1233),
.A2(n_1086),
.B(n_1159),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1125),
.A2(n_925),
.B(n_947),
.C(n_1108),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1101),
.Y(n_1391)
);

AOI221xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1125),
.A2(n_1202),
.B1(n_925),
.B2(n_839),
.C(n_1108),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1114),
.B(n_947),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1124),
.A2(n_1086),
.B(n_1052),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1124),
.A2(n_1100),
.B(n_1159),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1125),
.A2(n_925),
.B(n_947),
.C(n_1108),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1124),
.A2(n_1100),
.B(n_1159),
.Y(n_1398)
);

INVx8_ASAP7_75t_L g1399 ( 
.A(n_1139),
.Y(n_1399)
);

BUFx10_ASAP7_75t_L g1400 ( 
.A(n_1115),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1088),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1238),
.A2(n_1260),
.B1(n_1276),
.B2(n_1290),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1238),
.A2(n_1290),
.B1(n_1342),
.B2(n_1377),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1317),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1292),
.Y(n_1405)
);

BUFx12f_ASAP7_75t_L g1406 ( 
.A(n_1371),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1272),
.Y(n_1407)
);

BUFx8_ASAP7_75t_L g1408 ( 
.A(n_1369),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1269),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1280),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1265),
.A2(n_1333),
.B1(n_1386),
.B2(n_1281),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1342),
.A2(n_1345),
.B1(n_1330),
.B2(n_1241),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1379),
.A2(n_1392),
.B(n_1283),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1272),
.Y(n_1414)
);

BUFx8_ASAP7_75t_SL g1415 ( 
.A(n_1380),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1330),
.A2(n_1367),
.B1(n_1360),
.B2(n_1337),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1296),
.B(n_1244),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1245),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1344),
.B(n_1350),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1364),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1374),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1351),
.A2(n_1394),
.B1(n_1382),
.B2(n_1354),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1339),
.A2(n_1264),
.B1(n_1336),
.B2(n_1287),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1244),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1341),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1250),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1305),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1314),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1348),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1336),
.A2(n_1320),
.B1(n_1321),
.B2(n_1307),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1372),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1332),
.A2(n_1373),
.B1(n_1366),
.B2(n_1356),
.Y(n_1432)
);

INVx8_ASAP7_75t_L g1433 ( 
.A(n_1381),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1273),
.A2(n_1275),
.B(n_1363),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1392),
.A2(n_1309),
.B1(n_1310),
.B2(n_1322),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1401),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1332),
.A2(n_1356),
.B1(n_1373),
.B2(n_1366),
.Y(n_1437)
);

BUFx10_ASAP7_75t_L g1438 ( 
.A(n_1286),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1334),
.A2(n_1389),
.B1(n_1361),
.B2(n_1397),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1335),
.A2(n_1390),
.B(n_1384),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1352),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_1355),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1400),
.A2(n_1302),
.B1(n_1383),
.B2(n_1259),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1400),
.A2(n_1259),
.B1(n_1255),
.B2(n_1263),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1399),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1255),
.A2(n_1343),
.B1(n_1252),
.B2(n_1261),
.Y(n_1446)
);

BUFx12f_ASAP7_75t_L g1447 ( 
.A(n_1266),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1296),
.A2(n_1323),
.B1(n_1329),
.B2(n_1277),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1359),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1294),
.A2(n_1304),
.B1(n_1315),
.B2(n_1274),
.Y(n_1450)
);

INVx8_ASAP7_75t_L g1451 ( 
.A(n_1381),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1296),
.A2(n_1391),
.B1(n_1299),
.B2(n_1254),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1274),
.A2(n_1318),
.B1(n_1254),
.B2(n_1300),
.Y(n_1453)
);

BUFx4f_ASAP7_75t_SL g1454 ( 
.A(n_1311),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1284),
.A2(n_1285),
.B1(n_1271),
.B2(n_1289),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1284),
.A2(n_1285),
.B1(n_1271),
.B2(n_1278),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1327),
.B(n_1278),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1399),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1399),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1381),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1300),
.A2(n_1313),
.B1(n_1266),
.B2(n_1316),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1295),
.A2(n_1248),
.B(n_1247),
.Y(n_1462)
);

BUFx5_ASAP7_75t_L g1463 ( 
.A(n_1256),
.Y(n_1463)
);

BUFx2_ASAP7_75t_SL g1464 ( 
.A(n_1376),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1355),
.Y(n_1465)
);

CKINVDCx16_ASAP7_75t_R g1466 ( 
.A(n_1313),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1358),
.B(n_1378),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1319),
.A2(n_1388),
.B1(n_1256),
.B2(n_1381),
.Y(n_1468)
);

INVx6_ASAP7_75t_L g1469 ( 
.A(n_1271),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1285),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1256),
.A2(n_1388),
.B1(n_1324),
.B2(n_1325),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1293),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1270),
.A2(n_1347),
.B1(n_1288),
.B2(n_1251),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1324),
.B(n_1293),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1326),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1243),
.A2(n_1328),
.B1(n_1387),
.B2(n_1349),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1256),
.A2(n_1298),
.B1(n_1243),
.B2(n_1395),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1324),
.B(n_1357),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1306),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1340),
.A2(n_1365),
.B1(n_1393),
.B2(n_1375),
.Y(n_1480)
);

INVx4_ASAP7_75t_R g1481 ( 
.A(n_1267),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1346),
.A2(n_1370),
.B1(n_1362),
.B2(n_1279),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1242),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1308),
.Y(n_1484)
);

BUFx10_ASAP7_75t_L g1485 ( 
.A(n_1282),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1303),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1297),
.A2(n_1312),
.B1(n_1257),
.B2(n_1246),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1253),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1297),
.A2(n_1312),
.B1(n_1301),
.B2(n_1258),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1301),
.Y(n_1490)
);

CKINVDCx11_ASAP7_75t_R g1491 ( 
.A(n_1312),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1268),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1297),
.A2(n_1291),
.B1(n_1262),
.B2(n_1240),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1331),
.A2(n_1368),
.B1(n_1398),
.B2(n_1338),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1253),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1249),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1353),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1385),
.Y(n_1498)
);

BUFx8_ASAP7_75t_L g1499 ( 
.A(n_1396),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1260),
.A2(n_947),
.B1(n_1011),
.B2(n_910),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1333),
.B(n_1386),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1239),
.Y(n_1502)
);

BUFx12f_ASAP7_75t_L g1503 ( 
.A(n_1371),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1317),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1239),
.Y(n_1505)
);

BUFx12f_ASAP7_75t_L g1506 ( 
.A(n_1371),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_L g1507 ( 
.A(n_1371),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1239),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1260),
.A2(n_947),
.B1(n_1011),
.B2(n_910),
.Y(n_1509)
);

NAND2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1296),
.B(n_1244),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1250),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1238),
.A2(n_925),
.B1(n_808),
.B2(n_947),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1239),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1369),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1399),
.Y(n_1515)
);

INVx6_ASAP7_75t_L g1516 ( 
.A(n_1399),
.Y(n_1516)
);

BUFx10_ASAP7_75t_L g1517 ( 
.A(n_1286),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1371),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1239),
.Y(n_1519)
);

OAI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1290),
.A2(n_947),
.B1(n_651),
.B2(n_876),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1238),
.A2(n_925),
.B1(n_808),
.B2(n_947),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1272),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1400),
.A2(n_651),
.B1(n_736),
.B2(n_926),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1292),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1260),
.A2(n_947),
.B1(n_1011),
.B2(n_910),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1239),
.Y(n_1526)
);

BUFx8_ASAP7_75t_L g1527 ( 
.A(n_1317),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1333),
.B(n_1386),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1290),
.A2(n_947),
.B1(n_651),
.B2(n_876),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1272),
.Y(n_1530)
);

CKINVDCx11_ASAP7_75t_R g1531 ( 
.A(n_1317),
.Y(n_1531)
);

BUFx2_ASAP7_75t_R g1532 ( 
.A(n_1371),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1400),
.A2(n_651),
.B1(n_736),
.B2(n_926),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1239),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1239),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1239),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1239),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1272),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1400),
.A2(n_651),
.B1(n_736),
.B2(n_926),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1260),
.A2(n_947),
.B1(n_1011),
.B2(n_910),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1239),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_SL g1542 ( 
.A(n_1245),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1369),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1260),
.A2(n_926),
.B1(n_808),
.B2(n_925),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1333),
.B(n_1386),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1544),
.A2(n_1521),
.B(n_1512),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1440),
.A2(n_1476),
.B(n_1494),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1407),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1478),
.B(n_1432),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1475),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1488),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1407),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1476),
.A2(n_1482),
.B(n_1480),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1437),
.B(n_1491),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1501),
.B(n_1528),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1474),
.B(n_1484),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1452),
.B(n_1462),
.Y(n_1557)
);

CKINVDCx6p67_ASAP7_75t_R g1558 ( 
.A(n_1445),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1520),
.A2(n_1529),
.B(n_1434),
.Y(n_1559)
);

AOI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1452),
.A2(n_1498),
.B(n_1496),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1414),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1414),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1483),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1477),
.A2(n_1479),
.B(n_1473),
.Y(n_1564)
);

AO31x2_ASAP7_75t_L g1565 ( 
.A1(n_1487),
.A2(n_1489),
.A3(n_1495),
.B(n_1439),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1489),
.B(n_1487),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1469),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1479),
.A2(n_1473),
.B(n_1439),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1469),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1497),
.B(n_1490),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1402),
.A2(n_1539),
.B1(n_1533),
.B2(n_1523),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1434),
.A2(n_1403),
.B(n_1411),
.Y(n_1572)
);

AO21x2_ASAP7_75t_L g1573 ( 
.A1(n_1493),
.A2(n_1413),
.B(n_1462),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1459),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1459),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1425),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1429),
.Y(n_1577)
);

NAND2x1p5_ASAP7_75t_L g1578 ( 
.A(n_1460),
.B(n_1467),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1522),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1499),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1463),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1468),
.A2(n_1453),
.B(n_1455),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1441),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1412),
.A2(n_1435),
.B1(n_1444),
.B2(n_1416),
.C(n_1430),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1449),
.Y(n_1585)
);

AOI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1455),
.A2(n_1448),
.B(n_1456),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1499),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1492),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1463),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1486),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1471),
.B(n_1457),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1423),
.A2(n_1448),
.B(n_1509),
.Y(n_1592)
);

CKINVDCx11_ASAP7_75t_R g1593 ( 
.A(n_1404),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1485),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1485),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1426),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1522),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1409),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1410),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1500),
.A2(n_1540),
.B(n_1509),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1421),
.Y(n_1601)
);

BUFx12f_ASAP7_75t_L g1602 ( 
.A(n_1504),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_SL g1603 ( 
.A(n_1527),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1456),
.A2(n_1460),
.B(n_1461),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1502),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1505),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1508),
.B(n_1513),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1519),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1526),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1433),
.Y(n_1610)
);

AO21x2_ASAP7_75t_L g1611 ( 
.A1(n_1500),
.A2(n_1525),
.B(n_1540),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1534),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1535),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1545),
.B(n_1419),
.Y(n_1614)
);

NOR2x1_ASAP7_75t_R g1615 ( 
.A(n_1531),
.B(n_1436),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1536),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1525),
.A2(n_1422),
.B(n_1472),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1427),
.B(n_1541),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_SL g1619 ( 
.A1(n_1446),
.A2(n_1450),
.B(n_1443),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1417),
.A2(n_1510),
.B(n_1537),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1428),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1433),
.B(n_1451),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1530),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1530),
.B(n_1538),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1417),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1510),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1515),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1431),
.Y(n_1628)
);

CKINVDCx11_ASAP7_75t_R g1629 ( 
.A(n_1518),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1481),
.A2(n_1511),
.B(n_1538),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1408),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1515),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1424),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1466),
.B(n_1514),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1543),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1470),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1408),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_SL g1638 ( 
.A1(n_1405),
.A2(n_1524),
.B(n_1527),
.Y(n_1638)
);

INVx4_ASAP7_75t_L g1639 ( 
.A(n_1516),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1442),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1442),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1464),
.A2(n_1454),
.B(n_1447),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1438),
.B(n_1517),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1524),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1465),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1438),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1517),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1542),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1458),
.B(n_1418),
.Y(n_1649)
);

AO31x2_ASAP7_75t_L g1650 ( 
.A1(n_1542),
.A2(n_1532),
.A3(n_1420),
.B(n_1406),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1503),
.Y(n_1651)
);

INVxp33_ASAP7_75t_L g1652 ( 
.A(n_1415),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1506),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1507),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_SL g1655 ( 
.A(n_1557),
.B(n_1622),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1621),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1546),
.A2(n_1559),
.B(n_1571),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1621),
.B(n_1548),
.Y(n_1658)
);

OAI211xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1572),
.A2(n_1628),
.B(n_1555),
.C(n_1600),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1584),
.A2(n_1550),
.B(n_1582),
.C(n_1554),
.Y(n_1660)
);

AND2x6_ASAP7_75t_L g1661 ( 
.A(n_1587),
.B(n_1581),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1550),
.A2(n_1557),
.B1(n_1554),
.B2(n_1590),
.Y(n_1662)
);

A2O1A1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1550),
.A2(n_1582),
.B(n_1570),
.C(n_1604),
.Y(n_1663)
);

BUFx8_ASAP7_75t_SL g1664 ( 
.A(n_1602),
.Y(n_1664)
);

NOR3xp33_ASAP7_75t_SL g1665 ( 
.A(n_1638),
.B(n_1648),
.C(n_1647),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1630),
.Y(n_1666)
);

O2A1O1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1619),
.A2(n_1592),
.B(n_1557),
.C(n_1561),
.Y(n_1667)
);

A2O1A1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1570),
.A2(n_1553),
.B(n_1604),
.C(n_1568),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1621),
.B(n_1552),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1591),
.B(n_1634),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1623),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1596),
.B(n_1562),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1557),
.A2(n_1590),
.B1(n_1646),
.B2(n_1647),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1557),
.A2(n_1646),
.B1(n_1595),
.B2(n_1567),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1579),
.B(n_1597),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1568),
.A2(n_1564),
.B(n_1547),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1553),
.A2(n_1587),
.B(n_1642),
.C(n_1564),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1595),
.B(n_1549),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1566),
.A2(n_1587),
.B(n_1592),
.C(n_1595),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1586),
.A2(n_1617),
.B(n_1620),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1556),
.B(n_1581),
.Y(n_1681)
);

BUFx2_ASAP7_75t_SL g1682 ( 
.A(n_1631),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1576),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_SL g1684 ( 
.A(n_1622),
.B(n_1592),
.Y(n_1684)
);

NAND4xp25_ASAP7_75t_L g1685 ( 
.A(n_1624),
.B(n_1648),
.C(n_1607),
.D(n_1608),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1611),
.A2(n_1580),
.B1(n_1643),
.B2(n_1645),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1586),
.A2(n_1617),
.B(n_1620),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1630),
.B(n_1607),
.Y(n_1688)
);

AO32x2_ASAP7_75t_L g1689 ( 
.A1(n_1567),
.A2(n_1569),
.A3(n_1565),
.B1(n_1630),
.B2(n_1566),
.Y(n_1689)
);

OAI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1593),
.A2(n_1587),
.B(n_1580),
.C(n_1635),
.Y(n_1690)
);

AO21x1_ASAP7_75t_L g1691 ( 
.A1(n_1578),
.A2(n_1633),
.B(n_1612),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1594),
.B(n_1580),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1629),
.Y(n_1693)
);

OAI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1643),
.A2(n_1636),
.B(n_1606),
.C(n_1599),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1563),
.Y(n_1695)
);

AO21x2_ASAP7_75t_L g1696 ( 
.A1(n_1560),
.A2(n_1547),
.B(n_1573),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_R g1697 ( 
.A(n_1622),
.B(n_1594),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_SL g1698 ( 
.A(n_1622),
.B(n_1573),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1577),
.B(n_1583),
.Y(n_1699)
);

INVx5_ASAP7_75t_SL g1700 ( 
.A(n_1558),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1558),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1631),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_SL g1703 ( 
.A1(n_1574),
.A2(n_1575),
.B(n_1627),
.C(n_1632),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1611),
.A2(n_1619),
.B1(n_1573),
.B2(n_1602),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1642),
.A2(n_1625),
.B(n_1626),
.Y(n_1705)
);

AO32x2_ASAP7_75t_L g1706 ( 
.A1(n_1569),
.A2(n_1565),
.A3(n_1639),
.B1(n_1575),
.B2(n_1574),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1625),
.A2(n_1626),
.B(n_1640),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1625),
.A2(n_1626),
.B(n_1641),
.Y(n_1708)
);

NOR2xp67_ASAP7_75t_SL g1709 ( 
.A(n_1631),
.B(n_1645),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1710)
);

NAND2xp33_ASAP7_75t_L g1711 ( 
.A(n_1610),
.B(n_1627),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1609),
.B(n_1613),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1641),
.A2(n_1644),
.B(n_1578),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1598),
.A2(n_1612),
.B1(n_1616),
.B2(n_1608),
.C(n_1605),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1661),
.Y(n_1715)
);

NAND2x1_ASAP7_75t_L g1716 ( 
.A(n_1661),
.B(n_1589),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1688),
.B(n_1706),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1657),
.B(n_1641),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1666),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1666),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1565),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1710),
.B(n_1565),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1658),
.B(n_1669),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1679),
.B(n_1565),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1678),
.B(n_1565),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1695),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1659),
.A2(n_1653),
.B1(n_1651),
.B2(n_1645),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1660),
.A2(n_1603),
.B1(n_1622),
.B2(n_1578),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1678),
.B(n_1585),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1706),
.B(n_1551),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1706),
.B(n_1551),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1683),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1679),
.B(n_1675),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1705),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1689),
.B(n_1551),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1659),
.A2(n_1653),
.B1(n_1651),
.B2(n_1645),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1691),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1661),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1712),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1699),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1714),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1733),
.B(n_1694),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1715),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1730),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1725),
.B(n_1686),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1716),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1726),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1722),
.B(n_1668),
.Y(n_1748)
);

OAI33xp33_ASAP7_75t_L g1749 ( 
.A1(n_1741),
.A2(n_1673),
.A3(n_1662),
.B1(n_1667),
.B2(n_1656),
.B3(n_1674),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1717),
.B(n_1670),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1726),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1730),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1727),
.A2(n_1704),
.B1(n_1663),
.B2(n_1667),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1727),
.A2(n_1704),
.B(n_1694),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1715),
.B(n_1684),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1719),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1732),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1717),
.B(n_1698),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1717),
.B(n_1681),
.Y(n_1759)
);

AOI33xp33_ASAP7_75t_L g1760 ( 
.A1(n_1741),
.A2(n_1671),
.A3(n_1616),
.B1(n_1703),
.B2(n_1632),
.B3(n_1588),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1715),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1728),
.A2(n_1655),
.B1(n_1690),
.B2(n_1700),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1725),
.B(n_1707),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1723),
.B(n_1690),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1732),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1736),
.A2(n_1664),
.B1(n_1685),
.B2(n_1682),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1715),
.B(n_1677),
.Y(n_1767)
);

OAI21xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1724),
.A2(n_1713),
.B(n_1692),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1730),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1721),
.B(n_1733),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1724),
.A2(n_1696),
.B(n_1711),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1729),
.B(n_1708),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1736),
.B(n_1665),
.C(n_1709),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1731),
.Y(n_1774)
);

NOR3xp33_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1615),
.C(n_1680),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1687),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1721),
.B(n_1676),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1747),
.Y(n_1778)
);

INVxp67_ASAP7_75t_SL g1779 ( 
.A(n_1742),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1747),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1744),
.B(n_1752),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1742),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1751),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1763),
.B(n_1719),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1751),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1743),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1763),
.B(n_1745),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1757),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1745),
.B(n_1720),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1746),
.B(n_1738),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1770),
.B(n_1733),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1746),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1770),
.B(n_1734),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1757),
.Y(n_1794)
);

NOR3xp33_ASAP7_75t_SL g1795 ( 
.A(n_1749),
.B(n_1693),
.C(n_1718),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1758),
.B(n_1734),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1743),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1748),
.B(n_1734),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1769),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1765),
.Y(n_1800)
);

AND2x4_ASAP7_75t_SL g1801 ( 
.A(n_1743),
.B(n_1665),
.Y(n_1801)
);

OAI211xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1754),
.A2(n_1718),
.B(n_1724),
.C(n_1637),
.Y(n_1802)
);

INVx4_ASAP7_75t_L g1803 ( 
.A(n_1743),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1774),
.B(n_1731),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1774),
.B(n_1731),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1772),
.B(n_1720),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1772),
.B(n_1740),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1758),
.B(n_1735),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1778),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1779),
.B(n_1808),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1779),
.B(n_1746),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1781),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1778),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1808),
.B(n_1746),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1808),
.B(n_1804),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1781),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1780),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1756),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1804),
.B(n_1750),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1795),
.B(n_1754),
.C(n_1775),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1780),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1781),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1783),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1799),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1782),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1783),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1791),
.B(n_1748),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1791),
.B(n_1777),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1790),
.B(n_1755),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1785),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1785),
.Y(n_1831)
);

OR2x6_ASAP7_75t_L g1832 ( 
.A(n_1803),
.B(n_1753),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1787),
.B(n_1756),
.Y(n_1833)
);

INVxp67_ASAP7_75t_SL g1834 ( 
.A(n_1798),
.Y(n_1834)
);

NOR4xp25_ASAP7_75t_L g1835 ( 
.A(n_1782),
.B(n_1773),
.C(n_1753),
.D(n_1760),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1789),
.B(n_1776),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1786),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1788),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1789),
.B(n_1776),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1786),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1805),
.B(n_1759),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1799),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1788),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1794),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1790),
.B(n_1755),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1805),
.B(n_1759),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1794),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1797),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1784),
.B(n_1777),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1800),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1799),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1809),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1810),
.B(n_1829),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1809),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1848),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1813),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1810),
.B(n_1790),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1810),
.B(n_1790),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1815),
.B(n_1803),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1824),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1835),
.B(n_1764),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1825),
.B(n_1784),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1825),
.B(n_1806),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1829),
.B(n_1790),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1845),
.B(n_1796),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1813),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1845),
.B(n_1796),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1827),
.B(n_1834),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1817),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1835),
.B(n_1834),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1815),
.B(n_1797),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1827),
.B(n_1798),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1815),
.B(n_1803),
.Y(n_1873)
);

OAI21xp33_ASAP7_75t_L g1874 ( 
.A1(n_1820),
.A2(n_1802),
.B(n_1766),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1811),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1818),
.B(n_1806),
.Y(n_1876)
);

INVx4_ASAP7_75t_L g1877 ( 
.A(n_1832),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1841),
.B(n_1803),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1841),
.B(n_1801),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1820),
.B(n_1807),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1817),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1818),
.B(n_1807),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1821),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1841),
.B(n_1801),
.Y(n_1884)
);

NAND2xp33_ASAP7_75t_L g1885 ( 
.A(n_1837),
.B(n_1775),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1833),
.B(n_1793),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1846),
.B(n_1801),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1821),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1833),
.B(n_1837),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1861),
.A2(n_1832),
.B(n_1802),
.Y(n_1890)
);

O2A1O1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1870),
.A2(n_1832),
.B(n_1840),
.C(n_1749),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1872),
.B(n_1836),
.Y(n_1892)
);

NAND2x1_ASAP7_75t_L g1893 ( 
.A(n_1877),
.B(n_1879),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1853),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1874),
.A2(n_1832),
.B1(n_1762),
.B2(n_1773),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1852),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_SL g1897 ( 
.A1(n_1880),
.A2(n_1832),
.B1(n_1768),
.B2(n_1737),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1855),
.B(n_1840),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1899)
);

NAND4xp25_ASAP7_75t_L g1900 ( 
.A(n_1874),
.B(n_1766),
.C(n_1762),
.D(n_1771),
.Y(n_1900)
);

NAND2x1p5_ASAP7_75t_L g1901 ( 
.A(n_1877),
.B(n_1879),
.Y(n_1901)
);

XNOR2x1_ASAP7_75t_L g1902 ( 
.A(n_1884),
.B(n_1649),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1868),
.Y(n_1903)
);

OAI322xp33_ASAP7_75t_L g1904 ( 
.A1(n_1862),
.A2(n_1849),
.A3(n_1831),
.B1(n_1830),
.B2(n_1826),
.C1(n_1823),
.C2(n_1793),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1877),
.A2(n_1737),
.B1(n_1767),
.B2(n_1771),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1884),
.B(n_1846),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1852),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1885),
.A2(n_1768),
.B1(n_1836),
.B2(n_1839),
.C(n_1849),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1877),
.B(n_1839),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1862),
.A2(n_1767),
.B1(n_1701),
.B2(n_1700),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1854),
.Y(n_1911)
);

OAI32xp33_ASAP7_75t_L g1912 ( 
.A1(n_1863),
.A2(n_1828),
.A3(n_1814),
.B1(n_1816),
.B2(n_1822),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1887),
.A2(n_1767),
.B1(n_1761),
.B2(n_1811),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1868),
.A2(n_1767),
.B1(n_1761),
.B2(n_1755),
.Y(n_1914)
);

AND2x4_ASAP7_75t_SL g1915 ( 
.A(n_1887),
.B(n_1654),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1871),
.B(n_1846),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1906),
.B(n_1864),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1893),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1895),
.A2(n_1878),
.B1(n_1859),
.B2(n_1873),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1894),
.B(n_1872),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1896),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_SL g1922 ( 
.A1(n_1890),
.A2(n_1901),
.B1(n_1915),
.B2(n_1899),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1907),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1903),
.B(n_1889),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1911),
.Y(n_1925)
);

OAI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1900),
.A2(n_1863),
.B1(n_1889),
.B2(n_1875),
.C(n_1876),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1900),
.A2(n_1878),
.B(n_1873),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1898),
.Y(n_1928)
);

OAI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1891),
.A2(n_1875),
.B1(n_1876),
.B2(n_1882),
.C(n_1886),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1902),
.B(n_1864),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_1909),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1916),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1892),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1904),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1904),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1897),
.A2(n_1908),
.B(n_1905),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1910),
.B(n_1871),
.Y(n_1937)
);

OAI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1929),
.A2(n_1910),
.B1(n_1914),
.B2(n_1886),
.Y(n_1938)
);

XOR2x2_ASAP7_75t_L g1939 ( 
.A(n_1929),
.B(n_1615),
.Y(n_1939)
);

AOI21xp33_ASAP7_75t_SL g1940 ( 
.A1(n_1934),
.A2(n_1652),
.B(n_1913),
.Y(n_1940)
);

OA22x2_ASAP7_75t_SL g1941 ( 
.A1(n_1935),
.A2(n_1866),
.B1(n_1888),
.B2(n_1883),
.Y(n_1941)
);

AND2x2_ASAP7_75t_SL g1942 ( 
.A(n_1924),
.B(n_1859),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1917),
.B(n_1857),
.Y(n_1943)
);

AOI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1936),
.A2(n_1912),
.B1(n_1859),
.B2(n_1882),
.C(n_1883),
.Y(n_1944)
);

OAI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1919),
.A2(n_1857),
.B1(n_1858),
.B2(n_1859),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1922),
.A2(n_1653),
.B(n_1649),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1930),
.B(n_1858),
.Y(n_1947)
);

AOI211xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1918),
.A2(n_1888),
.B(n_1881),
.C(n_1869),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1931),
.B(n_1928),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1946),
.B(n_1933),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1947),
.B(n_1932),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1942),
.Y(n_1952)
);

NAND3xp33_ASAP7_75t_L g1953 ( 
.A(n_1948),
.B(n_1926),
.C(n_1937),
.Y(n_1953)
);

OAI211xp5_ASAP7_75t_SL g1954 ( 
.A1(n_1946),
.A2(n_1926),
.B(n_1937),
.C(n_1927),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1939),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1938),
.B(n_1920),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1949),
.Y(n_1957)
);

AOI21xp33_ASAP7_75t_L g1958 ( 
.A1(n_1945),
.A2(n_1923),
.B(n_1921),
.Y(n_1958)
);

AOI211xp5_ASAP7_75t_L g1959 ( 
.A1(n_1940),
.A2(n_1925),
.B(n_1881),
.C(n_1869),
.Y(n_1959)
);

A2O1A1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1953),
.A2(n_1944),
.B(n_1941),
.C(n_1943),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_R g1961 ( 
.A(n_1957),
.B(n_1702),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_1955),
.Y(n_1962)
);

OAI31xp33_ASAP7_75t_L g1963 ( 
.A1(n_1954),
.A2(n_1811),
.A3(n_1856),
.B(n_1866),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1956),
.A2(n_1856),
.B(n_1854),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1952),
.Y(n_1965)
);

AOI221xp5_ASAP7_75t_L g1966 ( 
.A1(n_1960),
.A2(n_1958),
.B1(n_1950),
.B2(n_1959),
.C(n_1951),
.Y(n_1966)
);

OAI211xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1963),
.A2(n_1860),
.B(n_1828),
.C(n_1700),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1962),
.A2(n_1811),
.B1(n_1831),
.B2(n_1823),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_SL g1969 ( 
.A1(n_1965),
.A2(n_1865),
.B(n_1867),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1964),
.A2(n_1860),
.B1(n_1865),
.B2(n_1867),
.C(n_1826),
.Y(n_1970)
);

OAI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1961),
.A2(n_1860),
.B(n_1639),
.C(n_1830),
.Y(n_1971)
);

AOI211xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1962),
.A2(n_1703),
.B(n_1814),
.C(n_1844),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1969),
.B(n_1814),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1968),
.B(n_1812),
.Y(n_1974)
);

AOI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1966),
.A2(n_1816),
.B1(n_1822),
.B2(n_1812),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1972),
.B(n_1819),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1971),
.Y(n_1977)
);

NOR2x1_ASAP7_75t_L g1978 ( 
.A(n_1967),
.B(n_1838),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1973),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1976),
.A2(n_1970),
.B1(n_1812),
.B2(n_1816),
.Y(n_1980)
);

XNOR2x1_ASAP7_75t_SL g1981 ( 
.A(n_1977),
.B(n_1792),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1978),
.B(n_1838),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1980),
.B(n_1975),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1983),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1984),
.B(n_1979),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1984),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1986),
.A2(n_1982),
.B(n_1974),
.Y(n_1987)
);

OAI22x1_ASAP7_75t_L g1988 ( 
.A1(n_1985),
.A2(n_1981),
.B1(n_1792),
.B2(n_1822),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1987),
.A2(n_1842),
.B(n_1824),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1988),
.A2(n_1851),
.B1(n_1824),
.B2(n_1842),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1989),
.A2(n_1851),
.B(n_1842),
.Y(n_1991)
);

OAI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1991),
.A2(n_1990),
.B(n_1851),
.Y(n_1992)
);

OAI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1992),
.A2(n_1792),
.B1(n_1850),
.B2(n_1847),
.Y(n_1993)
);

OAI221xp5_ASAP7_75t_R g1994 ( 
.A1(n_1993),
.A2(n_1650),
.B1(n_1697),
.B2(n_1850),
.C(n_1847),
.Y(n_1994)
);

AOI211xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1844),
.B(n_1843),
.C(n_1650),
.Y(n_1995)
);


endmodule