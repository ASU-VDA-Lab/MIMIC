module fake_jpeg_26127_n_168 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_43),
.B(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_27),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_17),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_36),
.B1(n_20),
.B2(n_19),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_70),
.B1(n_85),
.B2(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_21),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_42),
.B1(n_20),
.B2(n_19),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_26),
.B(n_15),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_82),
.B(n_1),
.C(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_30),
.B1(n_22),
.B2(n_26),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_18),
.B1(n_53),
.B2(n_3),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_83),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_28),
.B(n_9),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_55),
.B1(n_25),
.B2(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_68),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_106),
.B1(n_87),
.B2(n_72),
.Y(n_110)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_49),
.B1(n_16),
.B2(n_24),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_99),
.B1(n_101),
.B2(n_2),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_70),
.B1(n_75),
.B2(n_63),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_105),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_102),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_25),
.B1(n_16),
.B2(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_16),
.B1(n_39),
.B2(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_9),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_28),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_116),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_114),
.B(n_121),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_63),
.B1(n_64),
.B2(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_119),
.B1(n_121),
.B2(n_93),
.Y(n_123)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_118),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_64),
.B(n_53),
.C(n_79),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_64),
.B1(n_69),
.B2(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_6),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_126),
.B1(n_118),
.B2(n_111),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_105),
.B1(n_97),
.B2(n_101),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_130),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_90),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_97),
.C(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_117),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_113),
.B(n_120),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_135),
.A2(n_127),
.B(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_139),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_142),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_134),
.C(n_113),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_151),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_142),
.B(n_144),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_135),
.B(n_136),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_113),
.C(n_130),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_156),
.B(n_152),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_140),
.B(n_141),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_147),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_158),
.B(n_160),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_147),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_158),
.B(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_109),
.C(n_94),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_88),
.B(n_113),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_91),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_162),
.C(n_165),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_167),
.Y(n_168)
);


endmodule